
/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 19:04:52 2023
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module kanwa ( p_reset , m_clock , data_in33 , data_in34 , data_in35 , data_in36 , data_in37 , data_in38 , data_in39 , data_in40 , data_in41 , data_in42 , data_in43 , data_in44 , data_in45 , data_in46 , data_in47 , data_in48 , data_in49 , data_in50 , data_in51 , data_in52 , data_in53 , data_in54 , data_in55 , data_in56 , data_in57 , data_in58 , data_in59 , data_in60 , data_in61 , data_in62 , data_in65 , data_in66 , data_in67 , data_in68 , data_in69 , data_in70 , data_in71 , data_in72 , data_in73 , data_in74 , data_in75 , data_in76 , data_in77 , data_in78 , data_in79 , data_in80 , data_in81 , data_in82 , data_in83 , data_in84 , data_in85 , data_in86 , data_in87 , data_in88 , data_in89 , data_in90 , data_in91 , data_in92 , data_in93 , data_in94 , data_in97 , data_in98 , data_in99 , data_in100 , data_in101 , data_in102 , data_in103 , data_in104 , data_in105 , data_in106 , data_in107 , data_in108 , data_in109 , data_in110 , data_in111 , data_in112 , data_in113 , data_in114 , data_in115 , data_in116 , data_in117 , data_in118 , data_in119 , data_in120 , data_in121 , data_in122 , data_in123 , data_in124 , data_in125 , data_in126 , data_in129 , data_in130 , data_in131 , data_in132 , data_in133 , data_in134 , data_in135 , data_in136 , data_in137 , data_in138 , data_in139 , data_in140 , data_in141 , data_in142 , data_in143 , data_in144 , data_in145 , data_in146 , data_in147 , data_in148 , data_in149 , data_in150 , data_in151 , data_in152 , data_in153 , data_in154 , data_in155 , data_in156 , data_in157 , data_in158 , data_in161 , data_in162 , data_in163 , data_in164 , data_in165 , data_in166 , data_in167 , data_in168 , data_in169 , data_in170 , data_in171 , data_in172 , data_in173 , data_in174 , data_in175 , data_in176 , data_in177 , data_in178 , data_in179 , data_in180 , data_in181 , data_in182 , data_in183 , data_in184 , data_in185 , data_in186 , data_in187 , data_in188 , data_in189 , data_in190 , data_in193 , data_in194 , data_in195 , data_in196 , data_in197 , data_in198 , data_in199 , data_in200 , data_in201 , data_in202 , data_in203 , data_in204 , data_in205 , data_in206 , data_in207 , data_in208 , data_in209 , data_in210 , data_in211 , data_in212 , data_in213 , data_in214 , data_in215 , data_in216 , data_in217 , data_in218 , data_in219 , data_in220 , data_in221 , data_in222 , data_in225 , data_in226 , data_in227 , data_in228 , data_in229 , data_in230 , data_in231 , data_in232 , data_in233 , data_in234 , data_in235 , data_in236 , data_in237 , data_in238 , data_in239 , data_in240 , data_in241 , data_in242 , data_in243 , data_in244 , data_in245 , data_in246 , data_in247 , data_in248 , data_in249 , data_in250 , data_in251 , data_in252 , data_in253 , data_in254 , data_in257 , data_in258 , data_in259 , data_in260 , data_in261 , data_in262 , data_in263 , data_in264 , data_in265 , data_in266 , data_in267 , data_in268 , data_in269 , data_in270 , data_in271 , data_in272 , data_in273 , data_in274 , data_in275 , data_in276 , data_in277 , data_in278 , data_in279 , data_in280 , data_in281 , data_in282 , data_in283 , data_in284 , data_in285 , data_in286 , data_in289 , data_in290 , data_in291 , data_in292 , data_in293 , data_in294 , data_in295 , data_in296 , data_in297 , data_in298 , data_in299 , data_in300 , data_in301 , data_in302 , data_in303 , data_in304 , data_in305 , data_in306 , data_in307 , data_in308 , data_in309 , data_in310 , data_in311 , data_in312 , data_in313 , data_in314 , data_in315 , data_in316 , data_in317 , data_in318 , data_in321 , data_in322 , data_in323 , data_in324 , data_in325 , data_in326 , data_in327 , data_in328 , data_in329 , data_in330 , data_in331 , data_in332 , data_in333 , data_in334 , data_in335 , data_in336 , data_in337 , data_in338 , data_in339 , data_in340 , data_in341 , data_in342 , data_in343 , data_in344 , data_in345 , data_in346 , data_in347 , data_in348 , data_in349 , data_in350 , data_in353 , data_in354 , data_in355 , data_in356 , data_in357 , data_in358 , data_in359 , data_in360 , data_in361 , data_in362 , data_in363 , data_in364 , data_in365 , data_in366 , data_in367 , data_in368 , data_in369 , data_in370 , data_in371 , data_in372 , data_in373 , data_in374 , data_in375 , data_in376 , data_in377 , data_in378 , data_in379 , data_in380 , data_in381 , data_in382 , data_in385 , data_in386 , data_in387 , data_in388 , data_in389 , data_in390 , data_in391 , data_in392 , data_in393 , data_in394 , data_in395 , data_in396 , data_in397 , data_in398 , data_in399 , data_in400 , data_in401 , data_in402 , data_in403 , data_in404 , data_in405 , data_in406 , data_in407 , data_in408 , data_in409 , data_in410 , data_in411 , data_in412 , data_in413 , data_in414 , data_in417 , data_in418 , data_in419 , data_in420 , data_in421 , data_in422 , data_in423 , data_in424 , data_in425 , data_in426 , data_in427 , data_in428 , data_in429 , data_in430 , data_in431 , data_in432 , data_in433 , data_in434 , data_in435 , data_in436 , data_in437 , data_in438 , data_in439 , data_in440 , data_in441 , data_in442 , data_in443 , data_in444 , data_in445 , data_in446 , data_in449 , data_in450 , data_in451 , data_in452 , data_in453 , data_in454 , data_in455 , data_in456 , data_in457 , data_in458 , data_in459 , data_in460 , data_in461 , data_in462 , data_in463 , data_in464 , data_in465 , data_in466 , data_in467 , data_in468 , data_in469 , data_in470 , data_in471 , data_in472 , data_in473 , data_in474 , data_in475 , data_in476 , data_in477 , data_in478 , start , goal , data_out33 , data_out34 , data_out35 , data_out36 , data_out37 , data_out38 , data_out39 , data_out40 , data_out41 , data_out42 , data_out43 , data_out44 , data_out45 , data_out46 , data_out47 , data_out48 , data_out49 , data_out50 , data_out51 , data_out52 , data_out53 , data_out54 , data_out55 , data_out56 , data_out57 , data_out58 , data_out59 , data_out60 , data_out61 , data_out62 , data_out65 , data_out66 , data_out67 , data_out68 , data_out69 , data_out70 , data_out71 , data_out72 , data_out73 , data_out74 , data_out75 , data_out76 , data_out77 , data_out78 , data_out79 , data_out80 , data_out81 , data_out82 , data_out83 , data_out84 , data_out85 , data_out86 , data_out87 , data_out88 , data_out89 , data_out90 , data_out91 , data_out92 , data_out93 , data_out94 , data_out97 , data_out98 , data_out99 , data_out100 , data_out101 , data_out102 , data_out103 , data_out104 , data_out105 , data_out106 , data_out107 , data_out108 , data_out109 , data_out110 , data_out111 , data_out112 , data_out113 , data_out114 , data_out115 , data_out116 , data_out117 , data_out118 , data_out119 , data_out120 , data_out121 , data_out122 , data_out123 , data_out124 , data_out125 , data_out126 , data_out129 , data_out130 , data_out131 , data_out132 , data_out133 , data_out134 , data_out135 , data_out136 , data_out137 , data_out138 , data_out139 , data_out140 , data_out141 , data_out142 , data_out143 , data_out144 , data_out145 , data_out146 , data_out147 , data_out148 , data_out149 , data_out150 , data_out151 , data_out152 , data_out153 , data_out154 , data_out155 , data_out156 , data_out157 , data_out158 , data_out161 , data_out162 , data_out163 , data_out164 , data_out165 , data_out166 , data_out167 , data_out168 , data_out169 , data_out170 , data_out171 , data_out172 , data_out173 , data_out174 , data_out175 , data_out176 , data_out177 , data_out178 , data_out179 , data_out180 , data_out181 , data_out182 , data_out183 , data_out184 , data_out185 , data_out186 , data_out187 , data_out188 , data_out189 , data_out190 , data_out193 , data_out194 , data_out195 , data_out196 , data_out197 , data_out198 , data_out199 , data_out200 , data_out201 , data_out202 , data_out203 , data_out204 , data_out205 , data_out206 , data_out207 , data_out208 , data_out209 , data_out210 , data_out211 , data_out212 , data_out213 , data_out214 , data_out215 , data_out216 , data_out217 , data_out218 , data_out219 , data_out220 , data_out221 , data_out222 , data_out225 , data_out226 , data_out227 , data_out228 , data_out229 , data_out230 , data_out231 , data_out232 , data_out233 , data_out234 , data_out235 , data_out236 , data_out237 , data_out238 , data_out239 , data_out240 , data_out241 , data_out242 , data_out243 , data_out244 , data_out245 , data_out246 , data_out247 , data_out248 , data_out249 , data_out250 , data_out251 , data_out252 , data_out253 , data_out254 , data_out257 , data_out258 , data_out259 , data_out260 , data_out261 , data_out262 , data_out263 , data_out264 , data_out265 , data_out266 , data_out267 , data_out268 , data_out269 , data_out270 , data_out271 , data_out272 , data_out273 , data_out274 , data_out275 , data_out276 , data_out277 , data_out278 , data_out279 , data_out280 , data_out281 , data_out282 , data_out283 , data_out284 , data_out285 , data_out286 , data_out289 , data_out290 , data_out291 , data_out292 , data_out293 , data_out294 , data_out295 , data_out296 , data_out297 , data_out298 , data_out299 , data_out300 , data_out301 , data_out302 , data_out303 , data_out304 , data_out305 , data_out306 , data_out307 , data_out308 , data_out309 , data_out310 , data_out311 , data_out312 , data_out313 , data_out314 , data_out315 , data_out316 , data_out317 , data_out318 , data_out321 , data_out322 , data_out323 , data_out324 , data_out325 , data_out326 , data_out327 , data_out328 , data_out329 , data_out330 , data_out331 , data_out332 , data_out333 , data_out334 , data_out335 , data_out336 , data_out337 , data_out338 , data_out339 , data_out340 , data_out341 , data_out342 , data_out343 , data_out344 , data_out345 , data_out346 , data_out347 , data_out348 , data_out349 , data_out350 , data_out353 , data_out354 , data_out355 , data_out356 , data_out357 , data_out358 , data_out359 , data_out360 , data_out361 , data_out362 , data_out363 , data_out364 , data_out365 , data_out366 , data_out367 , data_out368 , data_out369 , data_out370 , data_out371 , data_out372 , data_out373 , data_out374 , data_out375 , data_out376 , data_out377 , data_out378 , data_out379 , data_out380 , data_out381 , data_out382 , data_out385 , data_out386 , data_out387 , data_out388 , data_out389 , data_out390 , data_out391 , data_out392 , data_out393 , data_out394 , data_out395 , data_out396 , data_out397 , data_out398 , data_out399 , data_out400 , data_out401 , data_out402 , data_out403 , data_out404 , data_out405 , data_out406 , data_out407 , data_out408 , data_out409 , data_out410 , data_out411 , data_out412 , data_out413 , data_out414 , data_out417 , data_out418 , data_out419 , data_out420 , data_out421 , data_out422 , data_out423 , data_out424 , data_out425 , data_out426 , data_out427 , data_out428 , data_out429 , data_out430 , data_out431 , data_out432 , data_out433 , data_out434 , data_out435 , data_out436 , data_out437 , data_out438 , data_out439 , data_out440 , data_out441 , data_out442 , data_out443 , data_out444 , data_out445 , data_out446 , data_out449 , data_out450 , data_out451 , data_out452 , data_out453 , data_out454 , data_out455 , data_out456 , data_out457 , data_out458 , data_out459 , data_out460 , data_out461 , data_out462 , data_out463 , data_out464 , data_out465 , data_out466 , data_out467 , data_out468 , data_out469 , data_out470 , data_out471 , data_out472 , data_out473 , data_out474 , data_out475 , data_out476 , data_out477 , data_out478 , in_do , out_do );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input [9:0] data_in33;
  wire [9:0] data_in33;
  input [9:0] data_in34;
  wire [9:0] data_in34;
  input [9:0] data_in35;
  wire [9:0] data_in35;
  input [9:0] data_in36;
  wire [9:0] data_in36;
  input [9:0] data_in37;
  wire [9:0] data_in37;
  input [9:0] data_in38;
  wire [9:0] data_in38;
  input [9:0] data_in39;
  wire [9:0] data_in39;
  input [9:0] data_in40;
  wire [9:0] data_in40;
  input [9:0] data_in41;
  wire [9:0] data_in41;
  input [9:0] data_in42;
  wire [9:0] data_in42;
  input [9:0] data_in43;
  wire [9:0] data_in43;
  input [9:0] data_in44;
  wire [9:0] data_in44;
  input [9:0] data_in45;
  wire [9:0] data_in45;
  input [9:0] data_in46;
  wire [9:0] data_in46;
  input [9:0] data_in47;
  wire [9:0] data_in47;
  input [9:0] data_in48;
  wire [9:0] data_in48;
  input [9:0] data_in49;
  wire [9:0] data_in49;
  input [9:0] data_in50;
  wire [9:0] data_in50;
  input [9:0] data_in51;
  wire [9:0] data_in51;
  input [9:0] data_in52;
  wire [9:0] data_in52;
  input [9:0] data_in53;
  wire [9:0] data_in53;
  input [9:0] data_in54;
  wire [9:0] data_in54;
  input [9:0] data_in55;
  wire [9:0] data_in55;
  input [9:0] data_in56;
  wire [9:0] data_in56;
  input [9:0] data_in57;
  wire [9:0] data_in57;
  input [9:0] data_in58;
  wire [9:0] data_in58;
  input [9:0] data_in59;
  wire [9:0] data_in59;
  input [9:0] data_in60;
  wire [9:0] data_in60;
  input [9:0] data_in61;
  wire [9:0] data_in61;
  input [9:0] data_in62;
  wire [9:0] data_in62;
  input [9:0] data_in65;
  wire [9:0] data_in65;
  input [9:0] data_in66;
  wire [9:0] data_in66;
  input [9:0] data_in67;
  wire [9:0] data_in67;
  input [9:0] data_in68;
  wire [9:0] data_in68;
  input [9:0] data_in69;
  wire [9:0] data_in69;
  input [9:0] data_in70;
  wire [9:0] data_in70;
  input [9:0] data_in71;
  wire [9:0] data_in71;
  input [9:0] data_in72;
  wire [9:0] data_in72;
  input [9:0] data_in73;
  wire [9:0] data_in73;
  input [9:0] data_in74;
  wire [9:0] data_in74;
  input [9:0] data_in75;
  wire [9:0] data_in75;
  input [9:0] data_in76;
  wire [9:0] data_in76;
  input [9:0] data_in77;
  wire [9:0] data_in77;
  input [9:0] data_in78;
  wire [9:0] data_in78;
  input [9:0] data_in79;
  wire [9:0] data_in79;
  input [9:0] data_in80;
  wire [9:0] data_in80;
  input [9:0] data_in81;
  wire [9:0] data_in81;
  input [9:0] data_in82;
  wire [9:0] data_in82;
  input [9:0] data_in83;
  wire [9:0] data_in83;
  input [9:0] data_in84;
  wire [9:0] data_in84;
  input [9:0] data_in85;
  wire [9:0] data_in85;
  input [9:0] data_in86;
  wire [9:0] data_in86;
  input [9:0] data_in87;
  wire [9:0] data_in87;
  input [9:0] data_in88;
  wire [9:0] data_in88;
  input [9:0] data_in89;
  wire [9:0] data_in89;
  input [9:0] data_in90;
  wire [9:0] data_in90;
  input [9:0] data_in91;
  wire [9:0] data_in91;
  input [9:0] data_in92;
  wire [9:0] data_in92;
  input [9:0] data_in93;
  wire [9:0] data_in93;
  input [9:0] data_in94;
  wire [9:0] data_in94;
  input [9:0] data_in97;
  wire [9:0] data_in97;
  input [9:0] data_in98;
  wire [9:0] data_in98;
  input [9:0] data_in99;
  wire [9:0] data_in99;
  input [9:0] data_in100;
  wire [9:0] data_in100;
  input [9:0] data_in101;
  wire [9:0] data_in101;
  input [9:0] data_in102;
  wire [9:0] data_in102;
  input [9:0] data_in103;
  wire [9:0] data_in103;
  input [9:0] data_in104;
  wire [9:0] data_in104;
  input [9:0] data_in105;
  wire [9:0] data_in105;
  input [9:0] data_in106;
  wire [9:0] data_in106;
  input [9:0] data_in107;
  wire [9:0] data_in107;
  input [9:0] data_in108;
  wire [9:0] data_in108;
  input [9:0] data_in109;
  wire [9:0] data_in109;
  input [9:0] data_in110;
  wire [9:0] data_in110;
  input [9:0] data_in111;
  wire [9:0] data_in111;
  input [9:0] data_in112;
  wire [9:0] data_in112;
  input [9:0] data_in113;
  wire [9:0] data_in113;
  input [9:0] data_in114;
  wire [9:0] data_in114;
  input [9:0] data_in115;
  wire [9:0] data_in115;
  input [9:0] data_in116;
  wire [9:0] data_in116;
  input [9:0] data_in117;
  wire [9:0] data_in117;
  input [9:0] data_in118;
  wire [9:0] data_in118;
  input [9:0] data_in119;
  wire [9:0] data_in119;
  input [9:0] data_in120;
  wire [9:0] data_in120;
  input [9:0] data_in121;
  wire [9:0] data_in121;
  input [9:0] data_in122;
  wire [9:0] data_in122;
  input [9:0] data_in123;
  wire [9:0] data_in123;
  input [9:0] data_in124;
  wire [9:0] data_in124;
  input [9:0] data_in125;
  wire [9:0] data_in125;
  input [9:0] data_in126;
  wire [9:0] data_in126;
  input [9:0] data_in129;
  wire [9:0] data_in129;
  input [9:0] data_in130;
  wire [9:0] data_in130;
  input [9:0] data_in131;
  wire [9:0] data_in131;
  input [9:0] data_in132;
  wire [9:0] data_in132;
  input [9:0] data_in133;
  wire [9:0] data_in133;
  input [9:0] data_in134;
  wire [9:0] data_in134;
  input [9:0] data_in135;
  wire [9:0] data_in135;
  input [9:0] data_in136;
  wire [9:0] data_in136;
  input [9:0] data_in137;
  wire [9:0] data_in137;
  input [9:0] data_in138;
  wire [9:0] data_in138;
  input [9:0] data_in139;
  wire [9:0] data_in139;
  input [9:0] data_in140;
  wire [9:0] data_in140;
  input [9:0] data_in141;
  wire [9:0] data_in141;
  input [9:0] data_in142;
  wire [9:0] data_in142;
  input [9:0] data_in143;
  wire [9:0] data_in143;
  input [9:0] data_in144;
  wire [9:0] data_in144;
  input [9:0] data_in145;
  wire [9:0] data_in145;
  input [9:0] data_in146;
  wire [9:0] data_in146;
  input [9:0] data_in147;
  wire [9:0] data_in147;
  input [9:0] data_in148;
  wire [9:0] data_in148;
  input [9:0] data_in149;
  wire [9:0] data_in149;
  input [9:0] data_in150;
  wire [9:0] data_in150;
  input [9:0] data_in151;
  wire [9:0] data_in151;
  input [9:0] data_in152;
  wire [9:0] data_in152;
  input [9:0] data_in153;
  wire [9:0] data_in153;
  input [9:0] data_in154;
  wire [9:0] data_in154;
  input [9:0] data_in155;
  wire [9:0] data_in155;
  input [9:0] data_in156;
  wire [9:0] data_in156;
  input [9:0] data_in157;
  wire [9:0] data_in157;
  input [9:0] data_in158;
  wire [9:0] data_in158;
  input [9:0] data_in161;
  wire [9:0] data_in161;
  input [9:0] data_in162;
  wire [9:0] data_in162;
  input [9:0] data_in163;
  wire [9:0] data_in163;
  input [9:0] data_in164;
  wire [9:0] data_in164;
  input [9:0] data_in165;
  wire [9:0] data_in165;
  input [9:0] data_in166;
  wire [9:0] data_in166;
  input [9:0] data_in167;
  wire [9:0] data_in167;
  input [9:0] data_in168;
  wire [9:0] data_in168;
  input [9:0] data_in169;
  wire [9:0] data_in169;
  input [9:0] data_in170;
  wire [9:0] data_in170;
  input [9:0] data_in171;
  wire [9:0] data_in171;
  input [9:0] data_in172;
  wire [9:0] data_in172;
  input [9:0] data_in173;
  wire [9:0] data_in173;
  input [9:0] data_in174;
  wire [9:0] data_in174;
  input [9:0] data_in175;
  wire [9:0] data_in175;
  input [9:0] data_in176;
  wire [9:0] data_in176;
  input [9:0] data_in177;
  wire [9:0] data_in177;
  input [9:0] data_in178;
  wire [9:0] data_in178;
  input [9:0] data_in179;
  wire [9:0] data_in179;
  input [9:0] data_in180;
  wire [9:0] data_in180;
  input [9:0] data_in181;
  wire [9:0] data_in181;
  input [9:0] data_in182;
  wire [9:0] data_in182;
  input [9:0] data_in183;
  wire [9:0] data_in183;
  input [9:0] data_in184;
  wire [9:0] data_in184;
  input [9:0] data_in185;
  wire [9:0] data_in185;
  input [9:0] data_in186;
  wire [9:0] data_in186;
  input [9:0] data_in187;
  wire [9:0] data_in187;
  input [9:0] data_in188;
  wire [9:0] data_in188;
  input [9:0] data_in189;
  wire [9:0] data_in189;
  input [9:0] data_in190;
  wire [9:0] data_in190;
  input [9:0] data_in193;
  wire [9:0] data_in193;
  input [9:0] data_in194;
  wire [9:0] data_in194;
  input [9:0] data_in195;
  wire [9:0] data_in195;
  input [9:0] data_in196;
  wire [9:0] data_in196;
  input [9:0] data_in197;
  wire [9:0] data_in197;
  input [9:0] data_in198;
  wire [9:0] data_in198;
  input [9:0] data_in199;
  wire [9:0] data_in199;
  input [9:0] data_in200;
  wire [9:0] data_in200;
  input [9:0] data_in201;
  wire [9:0] data_in201;
  input [9:0] data_in202;
  wire [9:0] data_in202;
  input [9:0] data_in203;
  wire [9:0] data_in203;
  input [9:0] data_in204;
  wire [9:0] data_in204;
  input [9:0] data_in205;
  wire [9:0] data_in205;
  input [9:0] data_in206;
  wire [9:0] data_in206;
  input [9:0] data_in207;
  wire [9:0] data_in207;
  input [9:0] data_in208;
  wire [9:0] data_in208;
  input [9:0] data_in209;
  wire [9:0] data_in209;
  input [9:0] data_in210;
  wire [9:0] data_in210;
  input [9:0] data_in211;
  wire [9:0] data_in211;
  input [9:0] data_in212;
  wire [9:0] data_in212;
  input [9:0] data_in213;
  wire [9:0] data_in213;
  input [9:0] data_in214;
  wire [9:0] data_in214;
  input [9:0] data_in215;
  wire [9:0] data_in215;
  input [9:0] data_in216;
  wire [9:0] data_in216;
  input [9:0] data_in217;
  wire [9:0] data_in217;
  input [9:0] data_in218;
  wire [9:0] data_in218;
  input [9:0] data_in219;
  wire [9:0] data_in219;
  input [9:0] data_in220;
  wire [9:0] data_in220;
  input [9:0] data_in221;
  wire [9:0] data_in221;
  input [9:0] data_in222;
  wire [9:0] data_in222;
  input [9:0] data_in225;
  wire [9:0] data_in225;
  input [9:0] data_in226;
  wire [9:0] data_in226;
  input [9:0] data_in227;
  wire [9:0] data_in227;
  input [9:0] data_in228;
  wire [9:0] data_in228;
  input [9:0] data_in229;
  wire [9:0] data_in229;
  input [9:0] data_in230;
  wire [9:0] data_in230;
  input [9:0] data_in231;
  wire [9:0] data_in231;
  input [9:0] data_in232;
  wire [9:0] data_in232;
  input [9:0] data_in233;
  wire [9:0] data_in233;
  input [9:0] data_in234;
  wire [9:0] data_in234;
  input [9:0] data_in235;
  wire [9:0] data_in235;
  input [9:0] data_in236;
  wire [9:0] data_in236;
  input [9:0] data_in237;
  wire [9:0] data_in237;
  input [9:0] data_in238;
  wire [9:0] data_in238;
  input [9:0] data_in239;
  wire [9:0] data_in239;
  input [9:0] data_in240;
  wire [9:0] data_in240;
  input [9:0] data_in241;
  wire [9:0] data_in241;
  input [9:0] data_in242;
  wire [9:0] data_in242;
  input [9:0] data_in243;
  wire [9:0] data_in243;
  input [9:0] data_in244;
  wire [9:0] data_in244;
  input [9:0] data_in245;
  wire [9:0] data_in245;
  input [9:0] data_in246;
  wire [9:0] data_in246;
  input [9:0] data_in247;
  wire [9:0] data_in247;
  input [9:0] data_in248;
  wire [9:0] data_in248;
  input [9:0] data_in249;
  wire [9:0] data_in249;
  input [9:0] data_in250;
  wire [9:0] data_in250;
  input [9:0] data_in251;
  wire [9:0] data_in251;
  input [9:0] data_in252;
  wire [9:0] data_in252;
  input [9:0] data_in253;
  wire [9:0] data_in253;
  input [9:0] data_in254;
  wire [9:0] data_in254;
  input [9:0] data_in257;
  wire [9:0] data_in257;
  input [9:0] data_in258;
  wire [9:0] data_in258;
  input [9:0] data_in259;
  wire [9:0] data_in259;
  input [9:0] data_in260;
  wire [9:0] data_in260;
  input [9:0] data_in261;
  wire [9:0] data_in261;
  input [9:0] data_in262;
  wire [9:0] data_in262;
  input [9:0] data_in263;
  wire [9:0] data_in263;
  input [9:0] data_in264;
  wire [9:0] data_in264;
  input [9:0] data_in265;
  wire [9:0] data_in265;
  input [9:0] data_in266;
  wire [9:0] data_in266;
  input [9:0] data_in267;
  wire [9:0] data_in267;
  input [9:0] data_in268;
  wire [9:0] data_in268;
  input [9:0] data_in269;
  wire [9:0] data_in269;
  input [9:0] data_in270;
  wire [9:0] data_in270;
  input [9:0] data_in271;
  wire [9:0] data_in271;
  input [9:0] data_in272;
  wire [9:0] data_in272;
  input [9:0] data_in273;
  wire [9:0] data_in273;
  input [9:0] data_in274;
  wire [9:0] data_in274;
  input [9:0] data_in275;
  wire [9:0] data_in275;
  input [9:0] data_in276;
  wire [9:0] data_in276;
  input [9:0] data_in277;
  wire [9:0] data_in277;
  input [9:0] data_in278;
  wire [9:0] data_in278;
  input [9:0] data_in279;
  wire [9:0] data_in279;
  input [9:0] data_in280;
  wire [9:0] data_in280;
  input [9:0] data_in281;
  wire [9:0] data_in281;
  input [9:0] data_in282;
  wire [9:0] data_in282;
  input [9:0] data_in283;
  wire [9:0] data_in283;
  input [9:0] data_in284;
  wire [9:0] data_in284;
  input [9:0] data_in285;
  wire [9:0] data_in285;
  input [9:0] data_in286;
  wire [9:0] data_in286;
  input [9:0] data_in289;
  wire [9:0] data_in289;
  input [9:0] data_in290;
  wire [9:0] data_in290;
  input [9:0] data_in291;
  wire [9:0] data_in291;
  input [9:0] data_in292;
  wire [9:0] data_in292;
  input [9:0] data_in293;
  wire [9:0] data_in293;
  input [9:0] data_in294;
  wire [9:0] data_in294;
  input [9:0] data_in295;
  wire [9:0] data_in295;
  input [9:0] data_in296;
  wire [9:0] data_in296;
  input [9:0] data_in297;
  wire [9:0] data_in297;
  input [9:0] data_in298;
  wire [9:0] data_in298;
  input [9:0] data_in299;
  wire [9:0] data_in299;
  input [9:0] data_in300;
  wire [9:0] data_in300;
  input [9:0] data_in301;
  wire [9:0] data_in301;
  input [9:0] data_in302;
  wire [9:0] data_in302;
  input [9:0] data_in303;
  wire [9:0] data_in303;
  input [9:0] data_in304;
  wire [9:0] data_in304;
  input [9:0] data_in305;
  wire [9:0] data_in305;
  input [9:0] data_in306;
  wire [9:0] data_in306;
  input [9:0] data_in307;
  wire [9:0] data_in307;
  input [9:0] data_in308;
  wire [9:0] data_in308;
  input [9:0] data_in309;
  wire [9:0] data_in309;
  input [9:0] data_in310;
  wire [9:0] data_in310;
  input [9:0] data_in311;
  wire [9:0] data_in311;
  input [9:0] data_in312;
  wire [9:0] data_in312;
  input [9:0] data_in313;
  wire [9:0] data_in313;
  input [9:0] data_in314;
  wire [9:0] data_in314;
  input [9:0] data_in315;
  wire [9:0] data_in315;
  input [9:0] data_in316;
  wire [9:0] data_in316;
  input [9:0] data_in317;
  wire [9:0] data_in317;
  input [9:0] data_in318;
  wire [9:0] data_in318;
  input [9:0] data_in321;
  wire [9:0] data_in321;
  input [9:0] data_in322;
  wire [9:0] data_in322;
  input [9:0] data_in323;
  wire [9:0] data_in323;
  input [9:0] data_in324;
  wire [9:0] data_in324;
  input [9:0] data_in325;
  wire [9:0] data_in325;
  input [9:0] data_in326;
  wire [9:0] data_in326;
  input [9:0] data_in327;
  wire [9:0] data_in327;
  input [9:0] data_in328;
  wire [9:0] data_in328;
  input [9:0] data_in329;
  wire [9:0] data_in329;
  input [9:0] data_in330;
  wire [9:0] data_in330;
  input [9:0] data_in331;
  wire [9:0] data_in331;
  input [9:0] data_in332;
  wire [9:0] data_in332;
  input [9:0] data_in333;
  wire [9:0] data_in333;
  input [9:0] data_in334;
  wire [9:0] data_in334;
  input [9:0] data_in335;
  wire [9:0] data_in335;
  input [9:0] data_in336;
  wire [9:0] data_in336;
  input [9:0] data_in337;
  wire [9:0] data_in337;
  input [9:0] data_in338;
  wire [9:0] data_in338;
  input [9:0] data_in339;
  wire [9:0] data_in339;
  input [9:0] data_in340;
  wire [9:0] data_in340;
  input [9:0] data_in341;
  wire [9:0] data_in341;
  input [9:0] data_in342;
  wire [9:0] data_in342;
  input [9:0] data_in343;
  wire [9:0] data_in343;
  input [9:0] data_in344;
  wire [9:0] data_in344;
  input [9:0] data_in345;
  wire [9:0] data_in345;
  input [9:0] data_in346;
  wire [9:0] data_in346;
  input [9:0] data_in347;
  wire [9:0] data_in347;
  input [9:0] data_in348;
  wire [9:0] data_in348;
  input [9:0] data_in349;
  wire [9:0] data_in349;
  input [9:0] data_in350;
  wire [9:0] data_in350;
  input [9:0] data_in353;
  wire [9:0] data_in353;
  input [9:0] data_in354;
  wire [9:0] data_in354;
  input [9:0] data_in355;
  wire [9:0] data_in355;
  input [9:0] data_in356;
  wire [9:0] data_in356;
  input [9:0] data_in357;
  wire [9:0] data_in357;
  input [9:0] data_in358;
  wire [9:0] data_in358;
  input [9:0] data_in359;
  wire [9:0] data_in359;
  input [9:0] data_in360;
  wire [9:0] data_in360;
  input [9:0] data_in361;
  wire [9:0] data_in361;
  input [9:0] data_in362;
  wire [9:0] data_in362;
  input [9:0] data_in363;
  wire [9:0] data_in363;
  input [9:0] data_in364;
  wire [9:0] data_in364;
  input [9:0] data_in365;
  wire [9:0] data_in365;
  input [9:0] data_in366;
  wire [9:0] data_in366;
  input [9:0] data_in367;
  wire [9:0] data_in367;
  input [9:0] data_in368;
  wire [9:0] data_in368;
  input [9:0] data_in369;
  wire [9:0] data_in369;
  input [9:0] data_in370;
  wire [9:0] data_in370;
  input [9:0] data_in371;
  wire [9:0] data_in371;
  input [9:0] data_in372;
  wire [9:0] data_in372;
  input [9:0] data_in373;
  wire [9:0] data_in373;
  input [9:0] data_in374;
  wire [9:0] data_in374;
  input [9:0] data_in375;
  wire [9:0] data_in375;
  input [9:0] data_in376;
  wire [9:0] data_in376;
  input [9:0] data_in377;
  wire [9:0] data_in377;
  input [9:0] data_in378;
  wire [9:0] data_in378;
  input [9:0] data_in379;
  wire [9:0] data_in379;
  input [9:0] data_in380;
  wire [9:0] data_in380;
  input [9:0] data_in381;
  wire [9:0] data_in381;
  input [9:0] data_in382;
  wire [9:0] data_in382;
  input [9:0] data_in385;
  wire [9:0] data_in385;
  input [9:0] data_in386;
  wire [9:0] data_in386;
  input [9:0] data_in387;
  wire [9:0] data_in387;
  input [9:0] data_in388;
  wire [9:0] data_in388;
  input [9:0] data_in389;
  wire [9:0] data_in389;
  input [9:0] data_in390;
  wire [9:0] data_in390;
  input [9:0] data_in391;
  wire [9:0] data_in391;
  input [9:0] data_in392;
  wire [9:0] data_in392;
  input [9:0] data_in393;
  wire [9:0] data_in393;
  input [9:0] data_in394;
  wire [9:0] data_in394;
  input [9:0] data_in395;
  wire [9:0] data_in395;
  input [9:0] data_in396;
  wire [9:0] data_in396;
  input [9:0] data_in397;
  wire [9:0] data_in397;
  input [9:0] data_in398;
  wire [9:0] data_in398;
  input [9:0] data_in399;
  wire [9:0] data_in399;
  input [9:0] data_in400;
  wire [9:0] data_in400;
  input [9:0] data_in401;
  wire [9:0] data_in401;
  input [9:0] data_in402;
  wire [9:0] data_in402;
  input [9:0] data_in403;
  wire [9:0] data_in403;
  input [9:0] data_in404;
  wire [9:0] data_in404;
  input [9:0] data_in405;
  wire [9:0] data_in405;
  input [9:0] data_in406;
  wire [9:0] data_in406;
  input [9:0] data_in407;
  wire [9:0] data_in407;
  input [9:0] data_in408;
  wire [9:0] data_in408;
  input [9:0] data_in409;
  wire [9:0] data_in409;
  input [9:0] data_in410;
  wire [9:0] data_in410;
  input [9:0] data_in411;
  wire [9:0] data_in411;
  input [9:0] data_in412;
  wire [9:0] data_in412;
  input [9:0] data_in413;
  wire [9:0] data_in413;
  input [9:0] data_in414;
  wire [9:0] data_in414;
  input [9:0] data_in417;
  wire [9:0] data_in417;
  input [9:0] data_in418;
  wire [9:0] data_in418;
  input [9:0] data_in419;
  wire [9:0] data_in419;
  input [9:0] data_in420;
  wire [9:0] data_in420;
  input [9:0] data_in421;
  wire [9:0] data_in421;
  input [9:0] data_in422;
  wire [9:0] data_in422;
  input [9:0] data_in423;
  wire [9:0] data_in423;
  input [9:0] data_in424;
  wire [9:0] data_in424;
  input [9:0] data_in425;
  wire [9:0] data_in425;
  input [9:0] data_in426;
  wire [9:0] data_in426;
  input [9:0] data_in427;
  wire [9:0] data_in427;
  input [9:0] data_in428;
  wire [9:0] data_in428;
  input [9:0] data_in429;
  wire [9:0] data_in429;
  input [9:0] data_in430;
  wire [9:0] data_in430;
  input [9:0] data_in431;
  wire [9:0] data_in431;
  input [9:0] data_in432;
  wire [9:0] data_in432;
  input [9:0] data_in433;
  wire [9:0] data_in433;
  input [9:0] data_in434;
  wire [9:0] data_in434;
  input [9:0] data_in435;
  wire [9:0] data_in435;
  input [9:0] data_in436;
  wire [9:0] data_in436;
  input [9:0] data_in437;
  wire [9:0] data_in437;
  input [9:0] data_in438;
  wire [9:0] data_in438;
  input [9:0] data_in439;
  wire [9:0] data_in439;
  input [9:0] data_in440;
  wire [9:0] data_in440;
  input [9:0] data_in441;
  wire [9:0] data_in441;
  input [9:0] data_in442;
  wire [9:0] data_in442;
  input [9:0] data_in443;
  wire [9:0] data_in443;
  input [9:0] data_in444;
  wire [9:0] data_in444;
  input [9:0] data_in445;
  wire [9:0] data_in445;
  input [9:0] data_in446;
  wire [9:0] data_in446;
  input [9:0] data_in449;
  wire [9:0] data_in449;
  input [9:0] data_in450;
  wire [9:0] data_in450;
  input [9:0] data_in451;
  wire [9:0] data_in451;
  input [9:0] data_in452;
  wire [9:0] data_in452;
  input [9:0] data_in453;
  wire [9:0] data_in453;
  input [9:0] data_in454;
  wire [9:0] data_in454;
  input [9:0] data_in455;
  wire [9:0] data_in455;
  input [9:0] data_in456;
  wire [9:0] data_in456;
  input [9:0] data_in457;
  wire [9:0] data_in457;
  input [9:0] data_in458;
  wire [9:0] data_in458;
  input [9:0] data_in459;
  wire [9:0] data_in459;
  input [9:0] data_in460;
  wire [9:0] data_in460;
  input [9:0] data_in461;
  wire [9:0] data_in461;
  input [9:0] data_in462;
  wire [9:0] data_in462;
  input [9:0] data_in463;
  wire [9:0] data_in463;
  input [9:0] data_in464;
  wire [9:0] data_in464;
  input [9:0] data_in465;
  wire [9:0] data_in465;
  input [9:0] data_in466;
  wire [9:0] data_in466;
  input [9:0] data_in467;
  wire [9:0] data_in467;
  input [9:0] data_in468;
  wire [9:0] data_in468;
  input [9:0] data_in469;
  wire [9:0] data_in469;
  input [9:0] data_in470;
  wire [9:0] data_in470;
  input [9:0] data_in471;
  wire [9:0] data_in471;
  input [9:0] data_in472;
  wire [9:0] data_in472;
  input [9:0] data_in473;
  wire [9:0] data_in473;
  input [9:0] data_in474;
  wire [9:0] data_in474;
  input [9:0] data_in475;
  wire [9:0] data_in475;
  input [9:0] data_in476;
  wire [9:0] data_in476;
  input [9:0] data_in477;
  wire [9:0] data_in477;
  input [9:0] data_in478;
  wire [9:0] data_in478;
  input [9:0] start;
  wire [9:0] start;
  input [9:0] goal;
  wire [9:0] goal;
  output [9:0] data_out33;
  wire [9:0] data_out33;
  output [9:0] data_out34;
  wire [9:0] data_out34;
  output [9:0] data_out35;
  wire [9:0] data_out35;
  output [9:0] data_out36;
  wire [9:0] data_out36;
  output [9:0] data_out37;
  wire [9:0] data_out37;
  output [9:0] data_out38;
  wire [9:0] data_out38;
  output [9:0] data_out39;
  wire [9:0] data_out39;
  output [9:0] data_out40;
  wire [9:0] data_out40;
  output [9:0] data_out41;
  wire [9:0] data_out41;
  output [9:0] data_out42;
  wire [9:0] data_out42;
  output [9:0] data_out43;
  wire [9:0] data_out43;
  output [9:0] data_out44;
  wire [9:0] data_out44;
  output [9:0] data_out45;
  wire [9:0] data_out45;
  output [9:0] data_out46;
  wire [9:0] data_out46;
  output [9:0] data_out47;
  wire [9:0] data_out47;
  output [9:0] data_out48;
  wire [9:0] data_out48;
  output [9:0] data_out49;
  wire [9:0] data_out49;
  output [9:0] data_out50;
  wire [9:0] data_out50;
  output [9:0] data_out51;
  wire [9:0] data_out51;
  output [9:0] data_out52;
  wire [9:0] data_out52;
  output [9:0] data_out53;
  wire [9:0] data_out53;
  output [9:0] data_out54;
  wire [9:0] data_out54;
  output [9:0] data_out55;
  wire [9:0] data_out55;
  output [9:0] data_out56;
  wire [9:0] data_out56;
  output [9:0] data_out57;
  wire [9:0] data_out57;
  output [9:0] data_out58;
  wire [9:0] data_out58;
  output [9:0] data_out59;
  wire [9:0] data_out59;
  output [9:0] data_out60;
  wire [9:0] data_out60;
  output [9:0] data_out61;
  wire [9:0] data_out61;
  output [9:0] data_out62;
  wire [9:0] data_out62;
  output [9:0] data_out65;
  wire [9:0] data_out65;
  output [9:0] data_out66;
  wire [9:0] data_out66;
  output [9:0] data_out67;
  wire [9:0] data_out67;
  output [9:0] data_out68;
  wire [9:0] data_out68;
  output [9:0] data_out69;
  wire [9:0] data_out69;
  output [9:0] data_out70;
  wire [9:0] data_out70;
  output [9:0] data_out71;
  wire [9:0] data_out71;
  output [9:0] data_out72;
  wire [9:0] data_out72;
  output [9:0] data_out73;
  wire [9:0] data_out73;
  output [9:0] data_out74;
  wire [9:0] data_out74;
  output [9:0] data_out75;
  wire [9:0] data_out75;
  output [9:0] data_out76;
  wire [9:0] data_out76;
  output [9:0] data_out77;
  wire [9:0] data_out77;
  output [9:0] data_out78;
  wire [9:0] data_out78;
  output [9:0] data_out79;
  wire [9:0] data_out79;
  output [9:0] data_out80;
  wire [9:0] data_out80;
  output [9:0] data_out81;
  wire [9:0] data_out81;
  output [9:0] data_out82;
  wire [9:0] data_out82;
  output [9:0] data_out83;
  wire [9:0] data_out83;
  output [9:0] data_out84;
  wire [9:0] data_out84;
  output [9:0] data_out85;
  wire [9:0] data_out85;
  output [9:0] data_out86;
  wire [9:0] data_out86;
  output [9:0] data_out87;
  wire [9:0] data_out87;
  output [9:0] data_out88;
  wire [9:0] data_out88;
  output [9:0] data_out89;
  wire [9:0] data_out89;
  output [9:0] data_out90;
  wire [9:0] data_out90;
  output [9:0] data_out91;
  wire [9:0] data_out91;
  output [9:0] data_out92;
  wire [9:0] data_out92;
  output [9:0] data_out93;
  wire [9:0] data_out93;
  output [9:0] data_out94;
  wire [9:0] data_out94;
  output [9:0] data_out97;
  wire [9:0] data_out97;
  output [9:0] data_out98;
  wire [9:0] data_out98;
  output [9:0] data_out99;
  wire [9:0] data_out99;
  output [9:0] data_out100;
  wire [9:0] data_out100;
  output [9:0] data_out101;
  wire [9:0] data_out101;
  output [9:0] data_out102;
  wire [9:0] data_out102;
  output [9:0] data_out103;
  wire [9:0] data_out103;
  output [9:0] data_out104;
  wire [9:0] data_out104;
  output [9:0] data_out105;
  wire [9:0] data_out105;
  output [9:0] data_out106;
  wire [9:0] data_out106;
  output [9:0] data_out107;
  wire [9:0] data_out107;
  output [9:0] data_out108;
  wire [9:0] data_out108;
  output [9:0] data_out109;
  wire [9:0] data_out109;
  output [9:0] data_out110;
  wire [9:0] data_out110;
  output [9:0] data_out111;
  wire [9:0] data_out111;
  output [9:0] data_out112;
  wire [9:0] data_out112;
  output [9:0] data_out113;
  wire [9:0] data_out113;
  output [9:0] data_out114;
  wire [9:0] data_out114;
  output [9:0] data_out115;
  wire [9:0] data_out115;
  output [9:0] data_out116;
  wire [9:0] data_out116;
  output [9:0] data_out117;
  wire [9:0] data_out117;
  output [9:0] data_out118;
  wire [9:0] data_out118;
  output [9:0] data_out119;
  wire [9:0] data_out119;
  output [9:0] data_out120;
  wire [9:0] data_out120;
  output [9:0] data_out121;
  wire [9:0] data_out121;
  output [9:0] data_out122;
  wire [9:0] data_out122;
  output [9:0] data_out123;
  wire [9:0] data_out123;
  output [9:0] data_out124;
  wire [9:0] data_out124;
  output [9:0] data_out125;
  wire [9:0] data_out125;
  output [9:0] data_out126;
  wire [9:0] data_out126;
  output [9:0] data_out129;
  wire [9:0] data_out129;
  output [9:0] data_out130;
  wire [9:0] data_out130;
  output [9:0] data_out131;
  wire [9:0] data_out131;
  output [9:0] data_out132;
  wire [9:0] data_out132;
  output [9:0] data_out133;
  wire [9:0] data_out133;
  output [9:0] data_out134;
  wire [9:0] data_out134;
  output [9:0] data_out135;
  wire [9:0] data_out135;
  output [9:0] data_out136;
  wire [9:0] data_out136;
  output [9:0] data_out137;
  wire [9:0] data_out137;
  output [9:0] data_out138;
  wire [9:0] data_out138;
  output [9:0] data_out139;
  wire [9:0] data_out139;
  output [9:0] data_out140;
  wire [9:0] data_out140;
  output [9:0] data_out141;
  wire [9:0] data_out141;
  output [9:0] data_out142;
  wire [9:0] data_out142;
  output [9:0] data_out143;
  wire [9:0] data_out143;
  output [9:0] data_out144;
  wire [9:0] data_out144;
  output [9:0] data_out145;
  wire [9:0] data_out145;
  output [9:0] data_out146;
  wire [9:0] data_out146;
  output [9:0] data_out147;
  wire [9:0] data_out147;
  output [9:0] data_out148;
  wire [9:0] data_out148;
  output [9:0] data_out149;
  wire [9:0] data_out149;
  output [9:0] data_out150;
  wire [9:0] data_out150;
  output [9:0] data_out151;
  wire [9:0] data_out151;
  output [9:0] data_out152;
  wire [9:0] data_out152;
  output [9:0] data_out153;
  wire [9:0] data_out153;
  output [9:0] data_out154;
  wire [9:0] data_out154;
  output [9:0] data_out155;
  wire [9:0] data_out155;
  output [9:0] data_out156;
  wire [9:0] data_out156;
  output [9:0] data_out157;
  wire [9:0] data_out157;
  output [9:0] data_out158;
  wire [9:0] data_out158;
  output [9:0] data_out161;
  wire [9:0] data_out161;
  output [9:0] data_out162;
  wire [9:0] data_out162;
  output [9:0] data_out163;
  wire [9:0] data_out163;
  output [9:0] data_out164;
  wire [9:0] data_out164;
  output [9:0] data_out165;
  wire [9:0] data_out165;
  output [9:0] data_out166;
  wire [9:0] data_out166;
  output [9:0] data_out167;
  wire [9:0] data_out167;
  output [9:0] data_out168;
  wire [9:0] data_out168;
  output [9:0] data_out169;
  wire [9:0] data_out169;
  output [9:0] data_out170;
  wire [9:0] data_out170;
  output [9:0] data_out171;
  wire [9:0] data_out171;
  output [9:0] data_out172;
  wire [9:0] data_out172;
  output [9:0] data_out173;
  wire [9:0] data_out173;
  output [9:0] data_out174;
  wire [9:0] data_out174;
  output [9:0] data_out175;
  wire [9:0] data_out175;
  output [9:0] data_out176;
  wire [9:0] data_out176;
  output [9:0] data_out177;
  wire [9:0] data_out177;
  output [9:0] data_out178;
  wire [9:0] data_out178;
  output [9:0] data_out179;
  wire [9:0] data_out179;
  output [9:0] data_out180;
  wire [9:0] data_out180;
  output [9:0] data_out181;
  wire [9:0] data_out181;
  output [9:0] data_out182;
  wire [9:0] data_out182;
  output [9:0] data_out183;
  wire [9:0] data_out183;
  output [9:0] data_out184;
  wire [9:0] data_out184;
  output [9:0] data_out185;
  wire [9:0] data_out185;
  output [9:0] data_out186;
  wire [9:0] data_out186;
  output [9:0] data_out187;
  wire [9:0] data_out187;
  output [9:0] data_out188;
  wire [9:0] data_out188;
  output [9:0] data_out189;
  wire [9:0] data_out189;
  output [9:0] data_out190;
  wire [9:0] data_out190;
  output [9:0] data_out193;
  wire [9:0] data_out193;
  output [9:0] data_out194;
  wire [9:0] data_out194;
  output [9:0] data_out195;
  wire [9:0] data_out195;
  output [9:0] data_out196;
  wire [9:0] data_out196;
  output [9:0] data_out197;
  wire [9:0] data_out197;
  output [9:0] data_out198;
  wire [9:0] data_out198;
  output [9:0] data_out199;
  wire [9:0] data_out199;
  output [9:0] data_out200;
  wire [9:0] data_out200;
  output [9:0] data_out201;
  wire [9:0] data_out201;
  output [9:0] data_out202;
  wire [9:0] data_out202;
  output [9:0] data_out203;
  wire [9:0] data_out203;
  output [9:0] data_out204;
  wire [9:0] data_out204;
  output [9:0] data_out205;
  wire [9:0] data_out205;
  output [9:0] data_out206;
  wire [9:0] data_out206;
  output [9:0] data_out207;
  wire [9:0] data_out207;
  output [9:0] data_out208;
  wire [9:0] data_out208;
  output [9:0] data_out209;
  wire [9:0] data_out209;
  output [9:0] data_out210;
  wire [9:0] data_out210;
  output [9:0] data_out211;
  wire [9:0] data_out211;
  output [9:0] data_out212;
  wire [9:0] data_out212;
  output [9:0] data_out213;
  wire [9:0] data_out213;
  output [9:0] data_out214;
  wire [9:0] data_out214;
  output [9:0] data_out215;
  wire [9:0] data_out215;
  output [9:0] data_out216;
  wire [9:0] data_out216;
  output [9:0] data_out217;
  wire [9:0] data_out217;
  output [9:0] data_out218;
  wire [9:0] data_out218;
  output [9:0] data_out219;
  wire [9:0] data_out219;
  output [9:0] data_out220;
  wire [9:0] data_out220;
  output [9:0] data_out221;
  wire [9:0] data_out221;
  output [9:0] data_out222;
  wire [9:0] data_out222;
  output [9:0] data_out225;
  wire [9:0] data_out225;
  output [9:0] data_out226;
  wire [9:0] data_out226;
  output [9:0] data_out227;
  wire [9:0] data_out227;
  output [9:0] data_out228;
  wire [9:0] data_out228;
  output [9:0] data_out229;
  wire [9:0] data_out229;
  output [9:0] data_out230;
  wire [9:0] data_out230;
  output [9:0] data_out231;
  wire [9:0] data_out231;
  output [9:0] data_out232;
  wire [9:0] data_out232;
  output [9:0] data_out233;
  wire [9:0] data_out233;
  output [9:0] data_out234;
  wire [9:0] data_out234;
  output [9:0] data_out235;
  wire [9:0] data_out235;
  output [9:0] data_out236;
  wire [9:0] data_out236;
  output [9:0] data_out237;
  wire [9:0] data_out237;
  output [9:0] data_out238;
  wire [9:0] data_out238;
  output [9:0] data_out239;
  wire [9:0] data_out239;
  output [9:0] data_out240;
  wire [9:0] data_out240;
  output [9:0] data_out241;
  wire [9:0] data_out241;
  output [9:0] data_out242;
  wire [9:0] data_out242;
  output [9:0] data_out243;
  wire [9:0] data_out243;
  output [9:0] data_out244;
  wire [9:0] data_out244;
  output [9:0] data_out245;
  wire [9:0] data_out245;
  output [9:0] data_out246;
  wire [9:0] data_out246;
  output [9:0] data_out247;
  wire [9:0] data_out247;
  output [9:0] data_out248;
  wire [9:0] data_out248;
  output [9:0] data_out249;
  wire [9:0] data_out249;
  output [9:0] data_out250;
  wire [9:0] data_out250;
  output [9:0] data_out251;
  wire [9:0] data_out251;
  output [9:0] data_out252;
  wire [9:0] data_out252;
  output [9:0] data_out253;
  wire [9:0] data_out253;
  output [9:0] data_out254;
  wire [9:0] data_out254;
  output [9:0] data_out257;
  wire [9:0] data_out257;
  output [9:0] data_out258;
  wire [9:0] data_out258;
  output [9:0] data_out259;
  wire [9:0] data_out259;
  output [9:0] data_out260;
  wire [9:0] data_out260;
  output [9:0] data_out261;
  wire [9:0] data_out261;
  output [9:0] data_out262;
  wire [9:0] data_out262;
  output [9:0] data_out263;
  wire [9:0] data_out263;
  output [9:0] data_out264;
  wire [9:0] data_out264;
  output [9:0] data_out265;
  wire [9:0] data_out265;
  output [9:0] data_out266;
  wire [9:0] data_out266;
  output [9:0] data_out267;
  wire [9:0] data_out267;
  output [9:0] data_out268;
  wire [9:0] data_out268;
  output [9:0] data_out269;
  wire [9:0] data_out269;
  output [9:0] data_out270;
  wire [9:0] data_out270;
  output [9:0] data_out271;
  wire [9:0] data_out271;
  output [9:0] data_out272;
  wire [9:0] data_out272;
  output [9:0] data_out273;
  wire [9:0] data_out273;
  output [9:0] data_out274;
  wire [9:0] data_out274;
  output [9:0] data_out275;
  wire [9:0] data_out275;
  output [9:0] data_out276;
  wire [9:0] data_out276;
  output [9:0] data_out277;
  wire [9:0] data_out277;
  output [9:0] data_out278;
  wire [9:0] data_out278;
  output [9:0] data_out279;
  wire [9:0] data_out279;
  output [9:0] data_out280;
  wire [9:0] data_out280;
  output [9:0] data_out281;
  wire [9:0] data_out281;
  output [9:0] data_out282;
  wire [9:0] data_out282;
  output [9:0] data_out283;
  wire [9:0] data_out283;
  output [9:0] data_out284;
  wire [9:0] data_out284;
  output [9:0] data_out285;
  wire [9:0] data_out285;
  output [9:0] data_out286;
  wire [9:0] data_out286;
  output [9:0] data_out289;
  wire [9:0] data_out289;
  output [9:0] data_out290;
  wire [9:0] data_out290;
  output [9:0] data_out291;
  wire [9:0] data_out291;
  output [9:0] data_out292;
  wire [9:0] data_out292;
  output [9:0] data_out293;
  wire [9:0] data_out293;
  output [9:0] data_out294;
  wire [9:0] data_out294;
  output [9:0] data_out295;
  wire [9:0] data_out295;
  output [9:0] data_out296;
  wire [9:0] data_out296;
  output [9:0] data_out297;
  wire [9:0] data_out297;
  output [9:0] data_out298;
  wire [9:0] data_out298;
  output [9:0] data_out299;
  wire [9:0] data_out299;
  output [9:0] data_out300;
  wire [9:0] data_out300;
  output [9:0] data_out301;
  wire [9:0] data_out301;
  output [9:0] data_out302;
  wire [9:0] data_out302;
  output [9:0] data_out303;
  wire [9:0] data_out303;
  output [9:0] data_out304;
  wire [9:0] data_out304;
  output [9:0] data_out305;
  wire [9:0] data_out305;
  output [9:0] data_out306;
  wire [9:0] data_out306;
  output [9:0] data_out307;
  wire [9:0] data_out307;
  output [9:0] data_out308;
  wire [9:0] data_out308;
  output [9:0] data_out309;
  wire [9:0] data_out309;
  output [9:0] data_out310;
  wire [9:0] data_out310;
  output [9:0] data_out311;
  wire [9:0] data_out311;
  output [9:0] data_out312;
  wire [9:0] data_out312;
  output [9:0] data_out313;
  wire [9:0] data_out313;
  output [9:0] data_out314;
  wire [9:0] data_out314;
  output [9:0] data_out315;
  wire [9:0] data_out315;
  output [9:0] data_out316;
  wire [9:0] data_out316;
  output [9:0] data_out317;
  wire [9:0] data_out317;
  output [9:0] data_out318;
  wire [9:0] data_out318;
  output [9:0] data_out321;
  wire [9:0] data_out321;
  output [9:0] data_out322;
  wire [9:0] data_out322;
  output [9:0] data_out323;
  wire [9:0] data_out323;
  output [9:0] data_out324;
  wire [9:0] data_out324;
  output [9:0] data_out325;
  wire [9:0] data_out325;
  output [9:0] data_out326;
  wire [9:0] data_out326;
  output [9:0] data_out327;
  wire [9:0] data_out327;
  output [9:0] data_out328;
  wire [9:0] data_out328;
  output [9:0] data_out329;
  wire [9:0] data_out329;
  output [9:0] data_out330;
  wire [9:0] data_out330;
  output [9:0] data_out331;
  wire [9:0] data_out331;
  output [9:0] data_out332;
  wire [9:0] data_out332;
  output [9:0] data_out333;
  wire [9:0] data_out333;
  output [9:0] data_out334;
  wire [9:0] data_out334;
  output [9:0] data_out335;
  wire [9:0] data_out335;
  output [9:0] data_out336;
  wire [9:0] data_out336;
  output [9:0] data_out337;
  wire [9:0] data_out337;
  output [9:0] data_out338;
  wire [9:0] data_out338;
  output [9:0] data_out339;
  wire [9:0] data_out339;
  output [9:0] data_out340;
  wire [9:0] data_out340;
  output [9:0] data_out341;
  wire [9:0] data_out341;
  output [9:0] data_out342;
  wire [9:0] data_out342;
  output [9:0] data_out343;
  wire [9:0] data_out343;
  output [9:0] data_out344;
  wire [9:0] data_out344;
  output [9:0] data_out345;
  wire [9:0] data_out345;
  output [9:0] data_out346;
  wire [9:0] data_out346;
  output [9:0] data_out347;
  wire [9:0] data_out347;
  output [9:0] data_out348;
  wire [9:0] data_out348;
  output [9:0] data_out349;
  wire [9:0] data_out349;
  output [9:0] data_out350;
  wire [9:0] data_out350;
  output [9:0] data_out353;
  wire [9:0] data_out353;
  output [9:0] data_out354;
  wire [9:0] data_out354;
  output [9:0] data_out355;
  wire [9:0] data_out355;
  output [9:0] data_out356;
  wire [9:0] data_out356;
  output [9:0] data_out357;
  wire [9:0] data_out357;
  output [9:0] data_out358;
  wire [9:0] data_out358;
  output [9:0] data_out359;
  wire [9:0] data_out359;
  output [9:0] data_out360;
  wire [9:0] data_out360;
  output [9:0] data_out361;
  wire [9:0] data_out361;
  output [9:0] data_out362;
  wire [9:0] data_out362;
  output [9:0] data_out363;
  wire [9:0] data_out363;
  output [9:0] data_out364;
  wire [9:0] data_out364;
  output [9:0] data_out365;
  wire [9:0] data_out365;
  output [9:0] data_out366;
  wire [9:0] data_out366;
  output [9:0] data_out367;
  wire [9:0] data_out367;
  output [9:0] data_out368;
  wire [9:0] data_out368;
  output [9:0] data_out369;
  wire [9:0] data_out369;
  output [9:0] data_out370;
  wire [9:0] data_out370;
  output [9:0] data_out371;
  wire [9:0] data_out371;
  output [9:0] data_out372;
  wire [9:0] data_out372;
  output [9:0] data_out373;
  wire [9:0] data_out373;
  output [9:0] data_out374;
  wire [9:0] data_out374;
  output [9:0] data_out375;
  wire [9:0] data_out375;
  output [9:0] data_out376;
  wire [9:0] data_out376;
  output [9:0] data_out377;
  wire [9:0] data_out377;
  output [9:0] data_out378;
  wire [9:0] data_out378;
  output [9:0] data_out379;
  wire [9:0] data_out379;
  output [9:0] data_out380;
  wire [9:0] data_out380;
  output [9:0] data_out381;
  wire [9:0] data_out381;
  output [9:0] data_out382;
  wire [9:0] data_out382;
  output [9:0] data_out385;
  wire [9:0] data_out385;
  output [9:0] data_out386;
  wire [9:0] data_out386;
  output [9:0] data_out387;
  wire [9:0] data_out387;
  output [9:0] data_out388;
  wire [9:0] data_out388;
  output [9:0] data_out389;
  wire [9:0] data_out389;
  output [9:0] data_out390;
  wire [9:0] data_out390;
  output [9:0] data_out391;
  wire [9:0] data_out391;
  output [9:0] data_out392;
  wire [9:0] data_out392;
  output [9:0] data_out393;
  wire [9:0] data_out393;
  output [9:0] data_out394;
  wire [9:0] data_out394;
  output [9:0] data_out395;
  wire [9:0] data_out395;
  output [9:0] data_out396;
  wire [9:0] data_out396;
  output [9:0] data_out397;
  wire [9:0] data_out397;
  output [9:0] data_out398;
  wire [9:0] data_out398;
  output [9:0] data_out399;
  wire [9:0] data_out399;
  output [9:0] data_out400;
  wire [9:0] data_out400;
  output [9:0] data_out401;
  wire [9:0] data_out401;
  output [9:0] data_out402;
  wire [9:0] data_out402;
  output [9:0] data_out403;
  wire [9:0] data_out403;
  output [9:0] data_out404;
  wire [9:0] data_out404;
  output [9:0] data_out405;
  wire [9:0] data_out405;
  output [9:0] data_out406;
  wire [9:0] data_out406;
  output [9:0] data_out407;
  wire [9:0] data_out407;
  output [9:0] data_out408;
  wire [9:0] data_out408;
  output [9:0] data_out409;
  wire [9:0] data_out409;
  output [9:0] data_out410;
  wire [9:0] data_out410;
  output [9:0] data_out411;
  wire [9:0] data_out411;
  output [9:0] data_out412;
  wire [9:0] data_out412;
  output [9:0] data_out413;
  wire [9:0] data_out413;
  output [9:0] data_out414;
  wire [9:0] data_out414;
  output [9:0] data_out417;
  wire [9:0] data_out417;
  output [9:0] data_out418;
  wire [9:0] data_out418;
  output [9:0] data_out419;
  wire [9:0] data_out419;
  output [9:0] data_out420;
  wire [9:0] data_out420;
  output [9:0] data_out421;
  wire [9:0] data_out421;
  output [9:0] data_out422;
  wire [9:0] data_out422;
  output [9:0] data_out423;
  wire [9:0] data_out423;
  output [9:0] data_out424;
  wire [9:0] data_out424;
  output [9:0] data_out425;
  wire [9:0] data_out425;
  output [9:0] data_out426;
  wire [9:0] data_out426;
  output [9:0] data_out427;
  wire [9:0] data_out427;
  output [9:0] data_out428;
  wire [9:0] data_out428;
  output [9:0] data_out429;
  wire [9:0] data_out429;
  output [9:0] data_out430;
  wire [9:0] data_out430;
  output [9:0] data_out431;
  wire [9:0] data_out431;
  output [9:0] data_out432;
  wire [9:0] data_out432;
  output [9:0] data_out433;
  wire [9:0] data_out433;
  output [9:0] data_out434;
  wire [9:0] data_out434;
  output [9:0] data_out435;
  wire [9:0] data_out435;
  output [9:0] data_out436;
  wire [9:0] data_out436;
  output [9:0] data_out437;
  wire [9:0] data_out437;
  output [9:0] data_out438;
  wire [9:0] data_out438;
  output [9:0] data_out439;
  wire [9:0] data_out439;
  output [9:0] data_out440;
  wire [9:0] data_out440;
  output [9:0] data_out441;
  wire [9:0] data_out441;
  output [9:0] data_out442;
  wire [9:0] data_out442;
  output [9:0] data_out443;
  wire [9:0] data_out443;
  output [9:0] data_out444;
  wire [9:0] data_out444;
  output [9:0] data_out445;
  wire [9:0] data_out445;
  output [9:0] data_out446;
  wire [9:0] data_out446;
  output [9:0] data_out449;
  wire [9:0] data_out449;
  output [9:0] data_out450;
  wire [9:0] data_out450;
  output [9:0] data_out451;
  wire [9:0] data_out451;
  output [9:0] data_out452;
  wire [9:0] data_out452;
  output [9:0] data_out453;
  wire [9:0] data_out453;
  output [9:0] data_out454;
  wire [9:0] data_out454;
  output [9:0] data_out455;
  wire [9:0] data_out455;
  output [9:0] data_out456;
  wire [9:0] data_out456;
  output [9:0] data_out457;
  wire [9:0] data_out457;
  output [9:0] data_out458;
  wire [9:0] data_out458;
  output [9:0] data_out459;
  wire [9:0] data_out459;
  output [9:0] data_out460;
  wire [9:0] data_out460;
  output [9:0] data_out461;
  wire [9:0] data_out461;
  output [9:0] data_out462;
  wire [9:0] data_out462;
  output [9:0] data_out463;
  wire [9:0] data_out463;
  output [9:0] data_out464;
  wire [9:0] data_out464;
  output [9:0] data_out465;
  wire [9:0] data_out465;
  output [9:0] data_out466;
  wire [9:0] data_out466;
  output [9:0] data_out467;
  wire [9:0] data_out467;
  output [9:0] data_out468;
  wire [9:0] data_out468;
  output [9:0] data_out469;
  wire [9:0] data_out469;
  output [9:0] data_out470;
  wire [9:0] data_out470;
  output [9:0] data_out471;
  wire [9:0] data_out471;
  output [9:0] data_out472;
  wire [9:0] data_out472;
  output [9:0] data_out473;
  wire [9:0] data_out473;
  output [9:0] data_out474;
  wire [9:0] data_out474;
  output [9:0] data_out475;
  wire [9:0] data_out475;
  output [9:0] data_out476;
  wire [9:0] data_out476;
  output [9:0] data_out477;
  wire [9:0] data_out477;
  output [9:0] data_out478;
  wire [9:0] data_out478;
  input in_do;
  wire in_do;
  output out_do;
  wire out_do;
  wire dig_exit;
  reg [1:0] kanwa_exit;
  reg [9:0] start_reg;
  reg [9:0] goal_reg;
  reg even;
  wire even_w1;
  wire [9:0] start_wire;
  wire [9:0] goal_wire;
  wire wall_w;
  wire [9:0] data_wire33;
  wire [9:0] data_wire34;
  wire [9:0] data_wire35;
  wire [9:0] data_wire36;
  wire [9:0] data_wire37;
  wire [9:0] data_wire38;
  wire [9:0] data_wire39;
  wire [9:0] data_wire40;
  wire [9:0] data_wire41;
  wire [9:0] data_wire42;
  wire [9:0] data_wire43;
  wire [9:0] data_wire44;
  wire [9:0] data_wire45;
  wire [9:0] data_wire46;
  wire [9:0] data_wire47;
  wire [9:0] data_wire48;
  wire [9:0] data_wire49;
  wire [9:0] data_wire50;
  wire [9:0] data_wire51;
  wire [9:0] data_wire52;
  wire [9:0] data_wire53;
  wire [9:0] data_wire54;
  wire [9:0] data_wire55;
  wire [9:0] data_wire56;
  wire [9:0] data_wire57;
  wire [9:0] data_wire58;
  wire [9:0] data_wire59;
  wire [9:0] data_wire60;
  wire [9:0] data_wire61;
  wire [9:0] data_wire62;
  wire [9:0] data_wire65;
  wire [9:0] data_wire66;
  wire [9:0] data_wire67;
  wire [9:0] data_wire68;
  wire [9:0] data_wire69;
  wire [9:0] data_wire70;
  wire [9:0] data_wire71;
  wire [9:0] data_wire72;
  wire [9:0] data_wire73;
  wire [9:0] data_wire74;
  wire [9:0] data_wire75;
  wire [9:0] data_wire76;
  wire [9:0] data_wire77;
  wire [9:0] data_wire78;
  wire [9:0] data_wire79;
  wire [9:0] data_wire80;
  wire [9:0] data_wire81;
  wire [9:0] data_wire82;
  wire [9:0] data_wire83;
  wire [9:0] data_wire84;
  wire [9:0] data_wire85;
  wire [9:0] data_wire86;
  wire [9:0] data_wire87;
  wire [9:0] data_wire88;
  wire [9:0] data_wire89;
  wire [9:0] data_wire90;
  wire [9:0] data_wire91;
  wire [9:0] data_wire92;
  wire [9:0] data_wire93;
  wire [9:0] data_wire94;
  wire [9:0] data_wire97;
  wire [9:0] data_wire98;
  wire [9:0] data_wire99;
  wire [9:0] data_wire100;
  wire [9:0] data_wire101;
  wire [9:0] data_wire102;
  wire [9:0] data_wire103;
  wire [9:0] data_wire104;
  wire [9:0] data_wire105;
  wire [9:0] data_wire106;
  wire [9:0] data_wire107;
  wire [9:0] data_wire108;
  wire [9:0] data_wire109;
  wire [9:0] data_wire110;
  wire [9:0] data_wire111;
  wire [9:0] data_wire112;
  wire [9:0] data_wire113;
  wire [9:0] data_wire114;
  wire [9:0] data_wire115;
  wire [9:0] data_wire116;
  wire [9:0] data_wire117;
  wire [9:0] data_wire118;
  wire [9:0] data_wire119;
  wire [9:0] data_wire120;
  wire [9:0] data_wire121;
  wire [9:0] data_wire122;
  wire [9:0] data_wire123;
  wire [9:0] data_wire124;
  wire [9:0] data_wire125;
  wire [9:0] data_wire126;
  wire [9:0] data_wire129;
  wire [9:0] data_wire130;
  wire [9:0] data_wire131;
  wire [9:0] data_wire132;
  wire [9:0] data_wire133;
  wire [9:0] data_wire134;
  wire [9:0] data_wire135;
  wire [9:0] data_wire136;
  wire [9:0] data_wire137;
  wire [9:0] data_wire138;
  wire [9:0] data_wire139;
  wire [9:0] data_wire140;
  wire [9:0] data_wire141;
  wire [9:0] data_wire142;
  wire [9:0] data_wire143;
  wire [9:0] data_wire144;
  wire [9:0] data_wire145;
  wire [9:0] data_wire146;
  wire [9:0] data_wire147;
  wire [9:0] data_wire148;
  wire [9:0] data_wire149;
  wire [9:0] data_wire150;
  wire [9:0] data_wire151;
  wire [9:0] data_wire152;
  wire [9:0] data_wire153;
  wire [9:0] data_wire154;
  wire [9:0] data_wire155;
  wire [9:0] data_wire156;
  wire [9:0] data_wire157;
  wire [9:0] data_wire158;
  wire [9:0] data_wire161;
  wire [9:0] data_wire162;
  wire [9:0] data_wire163;
  wire [9:0] data_wire164;
  wire [9:0] data_wire165;
  wire [9:0] data_wire166;
  wire [9:0] data_wire167;
  wire [9:0] data_wire168;
  wire [9:0] data_wire169;
  wire [9:0] data_wire170;
  wire [9:0] data_wire171;
  wire [9:0] data_wire172;
  wire [9:0] data_wire173;
  wire [9:0] data_wire174;
  wire [9:0] data_wire175;
  wire [9:0] data_wire176;
  wire [9:0] data_wire177;
  wire [9:0] data_wire178;
  wire [9:0] data_wire179;
  wire [9:0] data_wire180;
  wire [9:0] data_wire181;
  wire [9:0] data_wire182;
  wire [9:0] data_wire183;
  wire [9:0] data_wire184;
  wire [9:0] data_wire185;
  wire [9:0] data_wire186;
  wire [9:0] data_wire187;
  wire [9:0] data_wire188;
  wire [9:0] data_wire189;
  wire [9:0] data_wire190;
  wire [9:0] data_wire193;
  wire [9:0] data_wire194;
  wire [9:0] data_wire195;
  wire [9:0] data_wire196;
  wire [9:0] data_wire197;
  wire [9:0] data_wire198;
  wire [9:0] data_wire199;
  wire [9:0] data_wire200;
  wire [9:0] data_wire201;
  wire [9:0] data_wire202;
  wire [9:0] data_wire203;
  wire [9:0] data_wire204;
  wire [9:0] data_wire205;
  wire [9:0] data_wire206;
  wire [9:0] data_wire207;
  wire [9:0] data_wire208;
  wire [9:0] data_wire209;
  wire [9:0] data_wire210;
  wire [9:0] data_wire211;
  wire [9:0] data_wire212;
  wire [9:0] data_wire213;
  wire [9:0] data_wire214;
  wire [9:0] data_wire215;
  wire [9:0] data_wire216;
  wire [9:0] data_wire217;
  wire [9:0] data_wire218;
  wire [9:0] data_wire219;
  wire [9:0] data_wire220;
  wire [9:0] data_wire221;
  wire [9:0] data_wire222;
  wire [9:0] data_wire225;
  wire [9:0] data_wire226;
  wire [9:0] data_wire227;
  wire [9:0] data_wire228;
  wire [9:0] data_wire229;
  wire [9:0] data_wire230;
  wire [9:0] data_wire231;
  wire [9:0] data_wire232;
  wire [9:0] data_wire233;
  wire [9:0] data_wire234;
  wire [9:0] data_wire235;
  wire [9:0] data_wire236;
  wire [9:0] data_wire237;
  wire [9:0] data_wire238;
  wire [9:0] data_wire239;
  wire [9:0] data_wire240;
  wire [9:0] data_wire241;
  wire [9:0] data_wire242;
  wire [9:0] data_wire243;
  wire [9:0] data_wire244;
  wire [9:0] data_wire245;
  wire [9:0] data_wire246;
  wire [9:0] data_wire247;
  wire [9:0] data_wire248;
  wire [9:0] data_wire249;
  wire [9:0] data_wire250;
  wire [9:0] data_wire251;
  wire [9:0] data_wire252;
  wire [9:0] data_wire253;
  wire [9:0] data_wire254;
  wire [9:0] data_wire257;
  wire [9:0] data_wire258;
  wire [9:0] data_wire259;
  wire [9:0] data_wire260;
  wire [9:0] data_wire261;
  wire [9:0] data_wire262;
  wire [9:0] data_wire263;
  wire [9:0] data_wire264;
  wire [9:0] data_wire265;
  wire [9:0] data_wire266;
  wire [9:0] data_wire267;
  wire [9:0] data_wire268;
  wire [9:0] data_wire269;
  wire [9:0] data_wire270;
  wire [9:0] data_wire271;
  wire [9:0] data_wire272;
  wire [9:0] data_wire273;
  wire [9:0] data_wire274;
  wire [9:0] data_wire275;
  wire [9:0] data_wire276;
  wire [9:0] data_wire277;
  wire [9:0] data_wire278;
  wire [9:0] data_wire279;
  wire [9:0] data_wire280;
  wire [9:0] data_wire281;
  wire [9:0] data_wire282;
  wire [9:0] data_wire283;
  wire [9:0] data_wire284;
  wire [9:0] data_wire285;
  wire [9:0] data_wire286;
  wire [9:0] data_wire289;
  wire [9:0] data_wire290;
  wire [9:0] data_wire291;
  wire [9:0] data_wire292;
  wire [9:0] data_wire293;
  wire [9:0] data_wire294;
  wire [9:0] data_wire295;
  wire [9:0] data_wire296;
  wire [9:0] data_wire297;
  wire [9:0] data_wire298;
  wire [9:0] data_wire299;
  wire [9:0] data_wire300;
  wire [9:0] data_wire301;
  wire [9:0] data_wire302;
  wire [9:0] data_wire303;
  wire [9:0] data_wire304;
  wire [9:0] data_wire305;
  wire [9:0] data_wire306;
  wire [9:0] data_wire307;
  wire [9:0] data_wire308;
  wire [9:0] data_wire309;
  wire [9:0] data_wire310;
  wire [9:0] data_wire311;
  wire [9:0] data_wire312;
  wire [9:0] data_wire313;
  wire [9:0] data_wire314;
  wire [9:0] data_wire315;
  wire [9:0] data_wire316;
  wire [9:0] data_wire317;
  wire [9:0] data_wire318;
  wire [9:0] data_wire321;
  wire [9:0] data_wire322;
  wire [9:0] data_wire323;
  wire [9:0] data_wire324;
  wire [9:0] data_wire325;
  wire [9:0] data_wire326;
  wire [9:0] data_wire327;
  wire [9:0] data_wire328;
  wire [9:0] data_wire329;
  wire [9:0] data_wire330;
  wire [9:0] data_wire331;
  wire [9:0] data_wire332;
  wire [9:0] data_wire333;
  wire [9:0] data_wire334;
  wire [9:0] data_wire335;
  wire [9:0] data_wire336;
  wire [9:0] data_wire337;
  wire [9:0] data_wire338;
  wire [9:0] data_wire339;
  wire [9:0] data_wire340;
  wire [9:0] data_wire341;
  wire [9:0] data_wire342;
  wire [9:0] data_wire343;
  wire [9:0] data_wire344;
  wire [9:0] data_wire345;
  wire [9:0] data_wire346;
  wire [9:0] data_wire347;
  wire [9:0] data_wire348;
  wire [9:0] data_wire349;
  wire [9:0] data_wire350;
  wire [9:0] data_wire353;
  wire [9:0] data_wire354;
  wire [9:0] data_wire355;
  wire [9:0] data_wire356;
  wire [9:0] data_wire357;
  wire [9:0] data_wire358;
  wire [9:0] data_wire359;
  wire [9:0] data_wire360;
  wire [9:0] data_wire361;
  wire [9:0] data_wire362;
  wire [9:0] data_wire363;
  wire [9:0] data_wire364;
  wire [9:0] data_wire365;
  wire [9:0] data_wire366;
  wire [9:0] data_wire367;
  wire [9:0] data_wire368;
  wire [9:0] data_wire369;
  wire [9:0] data_wire370;
  wire [9:0] data_wire371;
  wire [9:0] data_wire372;
  wire [9:0] data_wire373;
  wire [9:0] data_wire374;
  wire [9:0] data_wire375;
  wire [9:0] data_wire376;
  wire [9:0] data_wire377;
  wire [9:0] data_wire378;
  wire [9:0] data_wire379;
  wire [9:0] data_wire380;
  wire [9:0] data_wire381;
  wire [9:0] data_wire382;
  wire [9:0] data_wire385;
  wire [9:0] data_wire386;
  wire [9:0] data_wire387;
  wire [9:0] data_wire388;
  wire [9:0] data_wire389;
  wire [9:0] data_wire390;
  wire [9:0] data_wire391;
  wire [9:0] data_wire392;
  wire [9:0] data_wire393;
  wire [9:0] data_wire394;
  wire [9:0] data_wire395;
  wire [9:0] data_wire396;
  wire [9:0] data_wire397;
  wire [9:0] data_wire398;
  wire [9:0] data_wire399;
  wire [9:0] data_wire400;
  wire [9:0] data_wire401;
  wire [9:0] data_wire402;
  wire [9:0] data_wire403;
  wire [9:0] data_wire404;
  wire [9:0] data_wire405;
  wire [9:0] data_wire406;
  wire [9:0] data_wire407;
  wire [9:0] data_wire408;
  wire [9:0] data_wire409;
  wire [9:0] data_wire410;
  wire [9:0] data_wire411;
  wire [9:0] data_wire412;
  wire [9:0] data_wire413;
  wire [9:0] data_wire414;
  wire [9:0] data_wire417;
  wire [9:0] data_wire418;
  wire [9:0] data_wire419;
  wire [9:0] data_wire420;
  wire [9:0] data_wire421;
  wire [9:0] data_wire422;
  wire [9:0] data_wire423;
  wire [9:0] data_wire424;
  wire [9:0] data_wire425;
  wire [9:0] data_wire426;
  wire [9:0] data_wire427;
  wire [9:0] data_wire428;
  wire [9:0] data_wire429;
  wire [9:0] data_wire430;
  wire [9:0] data_wire431;
  wire [9:0] data_wire432;
  wire [9:0] data_wire433;
  wire [9:0] data_wire434;
  wire [9:0] data_wire435;
  wire [9:0] data_wire436;
  wire [9:0] data_wire437;
  wire [9:0] data_wire438;
  wire [9:0] data_wire439;
  wire [9:0] data_wire440;
  wire [9:0] data_wire441;
  wire [9:0] data_wire442;
  wire [9:0] data_wire443;
  wire [9:0] data_wire444;
  wire [9:0] data_wire445;
  wire [9:0] data_wire446;
  wire [9:0] data_wire449;
  wire [9:0] data_wire450;
  wire [9:0] data_wire451;
  wire [9:0] data_wire452;
  wire [9:0] data_wire453;
  wire [9:0] data_wire454;
  wire [9:0] data_wire455;
  wire [9:0] data_wire456;
  wire [9:0] data_wire457;
  wire [9:0] data_wire458;
  wire [9:0] data_wire459;
  wire [9:0] data_wire460;
  wire [9:0] data_wire461;
  wire [9:0] data_wire462;
  wire [9:0] data_wire463;
  wire [9:0] data_wire464;
  wire [9:0] data_wire465;
  wire [9:0] data_wire466;
  wire [9:0] data_wire467;
  wire [9:0] data_wire468;
  wire [9:0] data_wire469;
  wire [9:0] data_wire470;
  wire [9:0] data_wire471;
  wire [9:0] data_wire472;
  wire [9:0] data_wire473;
  wire [9:0] data_wire474;
  wire [9:0] data_wire475;
  wire [9:0] data_wire476;
  wire [9:0] data_wire477;
  wire [9:0] data_wire478;
  wire [9:0] data_out_org33;
  wire [9:0] data_out_org34;
  wire [9:0] data_out_org35;
  wire [9:0] data_out_org36;
  wire [9:0] data_out_org37;
  wire [9:0] data_out_org38;
  wire [9:0] data_out_org39;
  wire [9:0] data_out_org40;
  wire [9:0] data_out_org41;
  wire [9:0] data_out_org42;
  wire [9:0] data_out_org43;
  wire [9:0] data_out_org44;
  wire [9:0] data_out_org45;
  wire [9:0] data_out_org46;
  wire [9:0] data_out_org47;
  wire [9:0] data_out_org48;
  wire [9:0] data_out_org49;
  wire [9:0] data_out_org50;
  wire [9:0] data_out_org51;
  wire [9:0] data_out_org52;
  wire [9:0] data_out_org53;
  wire [9:0] data_out_org54;
  wire [9:0] data_out_org55;
  wire [9:0] data_out_org56;
  wire [9:0] data_out_org57;
  wire [9:0] data_out_org58;
  wire [9:0] data_out_org59;
  wire [9:0] data_out_org60;
  wire [9:0] data_out_org61;
  wire [9:0] data_out_org62;
  wire [9:0] data_out_org65;
  wire [9:0] data_out_org66;
  wire [9:0] data_out_org67;
  wire [9:0] data_out_org68;
  wire [9:0] data_out_org69;
  wire [9:0] data_out_org70;
  wire [9:0] data_out_org71;
  wire [9:0] data_out_org72;
  wire [9:0] data_out_org73;
  wire [9:0] data_out_org74;
  wire [9:0] data_out_org75;
  wire [9:0] data_out_org76;
  wire [9:0] data_out_org77;
  wire [9:0] data_out_org78;
  wire [9:0] data_out_org79;
  wire [9:0] data_out_org80;
  wire [9:0] data_out_org81;
  wire [9:0] data_out_org82;
  wire [9:0] data_out_org83;
  wire [9:0] data_out_org84;
  wire [9:0] data_out_org85;
  wire [9:0] data_out_org86;
  wire [9:0] data_out_org87;
  wire [9:0] data_out_org88;
  wire [9:0] data_out_org89;
  wire [9:0] data_out_org90;
  wire [9:0] data_out_org91;
  wire [9:0] data_out_org92;
  wire [9:0] data_out_org93;
  wire [9:0] data_out_org94;
  wire [9:0] data_out_org97;
  wire [9:0] data_out_org98;
  wire [9:0] data_out_org99;
  wire [9:0] data_out_org100;
  wire [9:0] data_out_org101;
  wire [9:0] data_out_org102;
  wire [9:0] data_out_org103;
  wire [9:0] data_out_org104;
  wire [9:0] data_out_org105;
  wire [9:0] data_out_org106;
  wire [9:0] data_out_org107;
  wire [9:0] data_out_org108;
  wire [9:0] data_out_org109;
  wire [9:0] data_out_org110;
  wire [9:0] data_out_org111;
  wire [9:0] data_out_org112;
  wire [9:0] data_out_org113;
  wire [9:0] data_out_org114;
  wire [9:0] data_out_org115;
  wire [9:0] data_out_org116;
  wire [9:0] data_out_org117;
  wire [9:0] data_out_org118;
  wire [9:0] data_out_org119;
  wire [9:0] data_out_org120;
  wire [9:0] data_out_org121;
  wire [9:0] data_out_org122;
  wire [9:0] data_out_org123;
  wire [9:0] data_out_org124;
  wire [9:0] data_out_org125;
  wire [9:0] data_out_org126;
  wire [9:0] data_out_org129;
  wire [9:0] data_out_org130;
  wire [9:0] data_out_org131;
  wire [9:0] data_out_org132;
  wire [9:0] data_out_org133;
  wire [9:0] data_out_org134;
  wire [9:0] data_out_org135;
  wire [9:0] data_out_org136;
  wire [9:0] data_out_org137;
  wire [9:0] data_out_org138;
  wire [9:0] data_out_org139;
  wire [9:0] data_out_org140;
  wire [9:0] data_out_org141;
  wire [9:0] data_out_org142;
  wire [9:0] data_out_org143;
  wire [9:0] data_out_org144;
  wire [9:0] data_out_org145;
  wire [9:0] data_out_org146;
  wire [9:0] data_out_org147;
  wire [9:0] data_out_org148;
  wire [9:0] data_out_org149;
  wire [9:0] data_out_org150;
  wire [9:0] data_out_org151;
  wire [9:0] data_out_org152;
  wire [9:0] data_out_org153;
  wire [9:0] data_out_org154;
  wire [9:0] data_out_org155;
  wire [9:0] data_out_org156;
  wire [9:0] data_out_org157;
  wire [9:0] data_out_org158;
  wire [9:0] data_out_org161;
  wire [9:0] data_out_org162;
  wire [9:0] data_out_org163;
  wire [9:0] data_out_org164;
  wire [9:0] data_out_org165;
  wire [9:0] data_out_org166;
  wire [9:0] data_out_org167;
  wire [9:0] data_out_org168;
  wire [9:0] data_out_org169;
  wire [9:0] data_out_org170;
  wire [9:0] data_out_org171;
  wire [9:0] data_out_org172;
  wire [9:0] data_out_org173;
  wire [9:0] data_out_org174;
  wire [9:0] data_out_org175;
  wire [9:0] data_out_org176;
  wire [9:0] data_out_org177;
  wire [9:0] data_out_org178;
  wire [9:0] data_out_org179;
  wire [9:0] data_out_org180;
  wire [9:0] data_out_org181;
  wire [9:0] data_out_org182;
  wire [9:0] data_out_org183;
  wire [9:0] data_out_org184;
  wire [9:0] data_out_org185;
  wire [9:0] data_out_org186;
  wire [9:0] data_out_org187;
  wire [9:0] data_out_org188;
  wire [9:0] data_out_org189;
  wire [9:0] data_out_org190;
  wire [9:0] data_out_org193;
  wire [9:0] data_out_org194;
  wire [9:0] data_out_org195;
  wire [9:0] data_out_org196;
  wire [9:0] data_out_org197;
  wire [9:0] data_out_org198;
  wire [9:0] data_out_org199;
  wire [9:0] data_out_org200;
  wire [9:0] data_out_org201;
  wire [9:0] data_out_org202;
  wire [9:0] data_out_org203;
  wire [9:0] data_out_org204;
  wire [9:0] data_out_org205;
  wire [9:0] data_out_org206;
  wire [9:0] data_out_org207;
  wire [9:0] data_out_org208;
  wire [9:0] data_out_org209;
  wire [9:0] data_out_org210;
  wire [9:0] data_out_org211;
  wire [9:0] data_out_org212;
  wire [9:0] data_out_org213;
  wire [9:0] data_out_org214;
  wire [9:0] data_out_org215;
  wire [9:0] data_out_org216;
  wire [9:0] data_out_org217;
  wire [9:0] data_out_org218;
  wire [9:0] data_out_org219;
  wire [9:0] data_out_org220;
  wire [9:0] data_out_org221;
  wire [9:0] data_out_org222;
  wire [9:0] data_out_org225;
  wire [9:0] data_out_org226;
  wire [9:0] data_out_org227;
  wire [9:0] data_out_org228;
  wire [9:0] data_out_org229;
  wire [9:0] data_out_org230;
  wire [9:0] data_out_org231;
  wire [9:0] data_out_org232;
  wire [9:0] data_out_org233;
  wire [9:0] data_out_org234;
  wire [9:0] data_out_org235;
  wire [9:0] data_out_org236;
  wire [9:0] data_out_org237;
  wire [9:0] data_out_org238;
  wire [9:0] data_out_org239;
  wire [9:0] data_out_org240;
  wire [9:0] data_out_org241;
  wire [9:0] data_out_org242;
  wire [9:0] data_out_org243;
  wire [9:0] data_out_org244;
  wire [9:0] data_out_org245;
  wire [9:0] data_out_org246;
  wire [9:0] data_out_org247;
  wire [9:0] data_out_org248;
  wire [9:0] data_out_org249;
  wire [9:0] data_out_org250;
  wire [9:0] data_out_org251;
  wire [9:0] data_out_org252;
  wire [9:0] data_out_org253;
  wire [9:0] data_out_org254;
  wire [9:0] data_out_org257;
  wire [9:0] data_out_org258;
  wire [9:0] data_out_org259;
  wire [9:0] data_out_org260;
  wire [9:0] data_out_org261;
  wire [9:0] data_out_org262;
  wire [9:0] data_out_org263;
  wire [9:0] data_out_org264;
  wire [9:0] data_out_org265;
  wire [9:0] data_out_org266;
  wire [9:0] data_out_org267;
  wire [9:0] data_out_org268;
  wire [9:0] data_out_org269;
  wire [9:0] data_out_org270;
  wire [9:0] data_out_org271;
  wire [9:0] data_out_org272;
  wire [9:0] data_out_org273;
  wire [9:0] data_out_org274;
  wire [9:0] data_out_org275;
  wire [9:0] data_out_org276;
  wire [9:0] data_out_org277;
  wire [9:0] data_out_org278;
  wire [9:0] data_out_org279;
  wire [9:0] data_out_org280;
  wire [9:0] data_out_org281;
  wire [9:0] data_out_org282;
  wire [9:0] data_out_org283;
  wire [9:0] data_out_org284;
  wire [9:0] data_out_org285;
  wire [9:0] data_out_org286;
  wire [9:0] data_out_org289;
  wire [9:0] data_out_org290;
  wire [9:0] data_out_org291;
  wire [9:0] data_out_org292;
  wire [9:0] data_out_org293;
  wire [9:0] data_out_org294;
  wire [9:0] data_out_org295;
  wire [9:0] data_out_org296;
  wire [9:0] data_out_org297;
  wire [9:0] data_out_org298;
  wire [9:0] data_out_org299;
  wire [9:0] data_out_org300;
  wire [9:0] data_out_org301;
  wire [9:0] data_out_org302;
  wire [9:0] data_out_org303;
  wire [9:0] data_out_org304;
  wire [9:0] data_out_org305;
  wire [9:0] data_out_org306;
  wire [9:0] data_out_org307;
  wire [9:0] data_out_org308;
  wire [9:0] data_out_org309;
  wire [9:0] data_out_org310;
  wire [9:0] data_out_org311;
  wire [9:0] data_out_org312;
  wire [9:0] data_out_org313;
  wire [9:0] data_out_org314;
  wire [9:0] data_out_org315;
  wire [9:0] data_out_org316;
  wire [9:0] data_out_org317;
  wire [9:0] data_out_org318;
  wire [9:0] data_out_org321;
  wire [9:0] data_out_org322;
  wire [9:0] data_out_org323;
  wire [9:0] data_out_org324;
  wire [9:0] data_out_org325;
  wire [9:0] data_out_org326;
  wire [9:0] data_out_org327;
  wire [9:0] data_out_org328;
  wire [9:0] data_out_org329;
  wire [9:0] data_out_org330;
  wire [9:0] data_out_org331;
  wire [9:0] data_out_org332;
  wire [9:0] data_out_org333;
  wire [9:0] data_out_org334;
  wire [9:0] data_out_org335;
  wire [9:0] data_out_org336;
  wire [9:0] data_out_org337;
  wire [9:0] data_out_org338;
  wire [9:0] data_out_org339;
  wire [9:0] data_out_org340;
  wire [9:0] data_out_org341;
  wire [9:0] data_out_org342;
  wire [9:0] data_out_org343;
  wire [9:0] data_out_org344;
  wire [9:0] data_out_org345;
  wire [9:0] data_out_org346;
  wire [9:0] data_out_org347;
  wire [9:0] data_out_org348;
  wire [9:0] data_out_org349;
  wire [9:0] data_out_org350;
  wire [9:0] data_out_org353;
  wire [9:0] data_out_org354;
  wire [9:0] data_out_org355;
  wire [9:0] data_out_org356;
  wire [9:0] data_out_org357;
  wire [9:0] data_out_org358;
  wire [9:0] data_out_org359;
  wire [9:0] data_out_org360;
  wire [9:0] data_out_org361;
  wire [9:0] data_out_org362;
  wire [9:0] data_out_org363;
  wire [9:0] data_out_org364;
  wire [9:0] data_out_org365;
  wire [9:0] data_out_org366;
  wire [9:0] data_out_org367;
  wire [9:0] data_out_org368;
  wire [9:0] data_out_org369;
  wire [9:0] data_out_org370;
  wire [9:0] data_out_org371;
  wire [9:0] data_out_org372;
  wire [9:0] data_out_org373;
  wire [9:0] data_out_org374;
  wire [9:0] data_out_org375;
  wire [9:0] data_out_org376;
  wire [9:0] data_out_org377;
  wire [9:0] data_out_org378;
  wire [9:0] data_out_org379;
  wire [9:0] data_out_org380;
  wire [9:0] data_out_org381;
  wire [9:0] data_out_org382;
  wire [9:0] data_out_org385;
  wire [9:0] data_out_org386;
  wire [9:0] data_out_org387;
  wire [9:0] data_out_org388;
  wire [9:0] data_out_org389;
  wire [9:0] data_out_org390;
  wire [9:0] data_out_org391;
  wire [9:0] data_out_org392;
  wire [9:0] data_out_org393;
  wire [9:0] data_out_org394;
  wire [9:0] data_out_org395;
  wire [9:0] data_out_org396;
  wire [9:0] data_out_org397;
  wire [9:0] data_out_org398;
  wire [9:0] data_out_org399;
  wire [9:0] data_out_org400;
  wire [9:0] data_out_org401;
  wire [9:0] data_out_org402;
  wire [9:0] data_out_org403;
  wire [9:0] data_out_org404;
  wire [9:0] data_out_org405;
  wire [9:0] data_out_org406;
  wire [9:0] data_out_org407;
  wire [9:0] data_out_org408;
  wire [9:0] data_out_org409;
  wire [9:0] data_out_org410;
  wire [9:0] data_out_org411;
  wire [9:0] data_out_org412;
  wire [9:0] data_out_org413;
  wire [9:0] data_out_org414;
  wire [9:0] data_out_org417;
  wire [9:0] data_out_org418;
  wire [9:0] data_out_org419;
  wire [9:0] data_out_org420;
  wire [9:0] data_out_org421;
  wire [9:0] data_out_org422;
  wire [9:0] data_out_org423;
  wire [9:0] data_out_org424;
  wire [9:0] data_out_org425;
  wire [9:0] data_out_org426;
  wire [9:0] data_out_org427;
  wire [9:0] data_out_org428;
  wire [9:0] data_out_org429;
  wire [9:0] data_out_org430;
  wire [9:0] data_out_org431;
  wire [9:0] data_out_org432;
  wire [9:0] data_out_org433;
  wire [9:0] data_out_org434;
  wire [9:0] data_out_org435;
  wire [9:0] data_out_org436;
  wire [9:0] data_out_org437;
  wire [9:0] data_out_org438;
  wire [9:0] data_out_org439;
  wire [9:0] data_out_org440;
  wire [9:0] data_out_org441;
  wire [9:0] data_out_org442;
  wire [9:0] data_out_org443;
  wire [9:0] data_out_org444;
  wire [9:0] data_out_org445;
  wire [9:0] data_out_org446;
  wire [9:0] data_out_org449;
  wire [9:0] data_out_org450;
  wire [9:0] data_out_org451;
  wire [9:0] data_out_org452;
  wire [9:0] data_out_org453;
  wire [9:0] data_out_org454;
  wire [9:0] data_out_org455;
  wire [9:0] data_out_org456;
  wire [9:0] data_out_org457;
  wire [9:0] data_out_org458;
  wire [9:0] data_out_org459;
  wire [9:0] data_out_org460;
  wire [9:0] data_out_org461;
  wire [9:0] data_out_org462;
  wire [9:0] data_out_org463;
  wire [9:0] data_out_org464;
  wire [9:0] data_out_org465;
  wire [9:0] data_out_org466;
  wire [9:0] data_out_org467;
  wire [9:0] data_out_org468;
  wire [9:0] data_out_org469;
  wire [9:0] data_out_org470;
  wire [9:0] data_out_org471;
  wire [9:0] data_out_org472;
  wire [9:0] data_out_org473;
  wire [9:0] data_out_org474;
  wire [9:0] data_out_org475;
  wire [9:0] data_out_org476;
  wire [9:0] data_out_org477;
  wire [9:0] data_out_org478;
  wire [1:0] sg33;
  wire [1:0] sg34;
  wire [1:0] sg35;
  wire [1:0] sg36;
  wire [1:0] sg37;
  wire [1:0] sg38;
  wire [1:0] sg39;
  wire [1:0] sg40;
  wire [1:0] sg41;
  wire [1:0] sg42;
  wire [1:0] sg43;
  wire [1:0] sg44;
  wire [1:0] sg45;
  wire [1:0] sg46;
  wire [1:0] sg47;
  wire [1:0] sg48;
  wire [1:0] sg49;
  wire [1:0] sg50;
  wire [1:0] sg51;
  wire [1:0] sg52;
  wire [1:0] sg53;
  wire [1:0] sg54;
  wire [1:0] sg55;
  wire [1:0] sg56;
  wire [1:0] sg57;
  wire [1:0] sg58;
  wire [1:0] sg59;
  wire [1:0] sg60;
  wire [1:0] sg61;
  wire [9:0] sg62;
  wire [1:0] sg65;
  wire [1:0] sg66;
  wire [1:0] sg67;
  wire [1:0] sg68;
  wire [1:0] sg69;
  wire [1:0] sg70;
  wire [1:0] sg71;
  wire [1:0] sg72;
  wire [1:0] sg73;
  wire [1:0] sg74;
  wire [1:0] sg75;
  wire [1:0] sg76;
  wire [1:0] sg77;
  wire [1:0] sg78;
  wire [1:0] sg79;
  wire [1:0] sg80;
  wire [1:0] sg81;
  wire [1:0] sg82;
  wire [1:0] sg83;
  wire [1:0] sg84;
  wire [1:0] sg85;
  wire [1:0] sg86;
  wire [1:0] sg87;
  wire [1:0] sg88;
  wire [1:0] sg89;
  wire [1:0] sg90;
  wire [1:0] sg91;
  wire [1:0] sg92;
  wire [1:0] sg93;
  wire [9:0] sg94;
  wire [1:0] sg97;
  wire [1:0] sg98;
  wire [1:0] sg99;
  wire [1:0] sg100;
  wire [1:0] sg101;
  wire [1:0] sg102;
  wire [1:0] sg103;
  wire [1:0] sg104;
  wire [1:0] sg105;
  wire [1:0] sg106;
  wire [1:0] sg107;
  wire [1:0] sg108;
  wire [1:0] sg109;
  wire [1:0] sg110;
  wire [1:0] sg111;
  wire [1:0] sg112;
  wire [1:0] sg113;
  wire [1:0] sg114;
  wire [1:0] sg115;
  wire [1:0] sg116;
  wire [1:0] sg117;
  wire [1:0] sg118;
  wire [1:0] sg119;
  wire [1:0] sg120;
  wire [1:0] sg121;
  wire [1:0] sg122;
  wire [1:0] sg123;
  wire [1:0] sg124;
  wire [1:0] sg125;
  wire [9:0] sg126;
  wire [1:0] sg129;
  wire [1:0] sg130;
  wire [1:0] sg131;
  wire [1:0] sg132;
  wire [1:0] sg133;
  wire [1:0] sg134;
  wire [1:0] sg135;
  wire [1:0] sg136;
  wire [1:0] sg137;
  wire [1:0] sg138;
  wire [1:0] sg139;
  wire [1:0] sg140;
  wire [1:0] sg141;
  wire [1:0] sg142;
  wire [1:0] sg143;
  wire [1:0] sg144;
  wire [1:0] sg145;
  wire [1:0] sg146;
  wire [1:0] sg147;
  wire [1:0] sg148;
  wire [1:0] sg149;
  wire [1:0] sg150;
  wire [1:0] sg151;
  wire [1:0] sg152;
  wire [1:0] sg153;
  wire [1:0] sg154;
  wire [1:0] sg155;
  wire [1:0] sg156;
  wire [1:0] sg157;
  wire [9:0] sg158;
  wire [1:0] sg161;
  wire [1:0] sg162;
  wire [1:0] sg163;
  wire [1:0] sg164;
  wire [1:0] sg165;
  wire [1:0] sg166;
  wire [1:0] sg167;
  wire [1:0] sg168;
  wire [1:0] sg169;
  wire [1:0] sg170;
  wire [1:0] sg171;
  wire [1:0] sg172;
  wire [1:0] sg173;
  wire [1:0] sg174;
  wire [1:0] sg175;
  wire [1:0] sg176;
  wire [1:0] sg177;
  wire [1:0] sg178;
  wire [1:0] sg179;
  wire [1:0] sg180;
  wire [1:0] sg181;
  wire [1:0] sg182;
  wire [1:0] sg183;
  wire [1:0] sg184;
  wire [1:0] sg185;
  wire [1:0] sg186;
  wire [1:0] sg187;
  wire [1:0] sg188;
  wire [1:0] sg189;
  wire [9:0] sg190;
  wire [1:0] sg193;
  wire [1:0] sg194;
  wire [1:0] sg195;
  wire [1:0] sg196;
  wire [1:0] sg197;
  wire [1:0] sg198;
  wire [1:0] sg199;
  wire [1:0] sg200;
  wire [1:0] sg201;
  wire [1:0] sg202;
  wire [1:0] sg203;
  wire [1:0] sg204;
  wire [1:0] sg205;
  wire [1:0] sg206;
  wire [1:0] sg207;
  wire [1:0] sg208;
  wire [1:0] sg209;
  wire [1:0] sg210;
  wire [1:0] sg211;
  wire [1:0] sg212;
  wire [1:0] sg213;
  wire [1:0] sg214;
  wire [1:0] sg215;
  wire [1:0] sg216;
  wire [1:0] sg217;
  wire [1:0] sg218;
  wire [1:0] sg219;
  wire [1:0] sg220;
  wire [1:0] sg221;
  wire [9:0] sg222;
  wire [1:0] sg225;
  wire [1:0] sg226;
  wire [1:0] sg227;
  wire [1:0] sg228;
  wire [1:0] sg229;
  wire [1:0] sg230;
  wire [1:0] sg231;
  wire [1:0] sg232;
  wire [1:0] sg233;
  wire [1:0] sg234;
  wire [1:0] sg235;
  wire [1:0] sg236;
  wire [1:0] sg237;
  wire [1:0] sg238;
  wire [1:0] sg239;
  wire [1:0] sg240;
  wire [1:0] sg241;
  wire [1:0] sg242;
  wire [1:0] sg243;
  wire [1:0] sg244;
  wire [1:0] sg245;
  wire [1:0] sg246;
  wire [1:0] sg247;
  wire [1:0] sg248;
  wire [1:0] sg249;
  wire [1:0] sg250;
  wire [1:0] sg251;
  wire [1:0] sg252;
  wire [1:0] sg253;
  wire [9:0] sg254;
  wire [1:0] sg257;
  wire [1:0] sg258;
  wire [1:0] sg259;
  wire [1:0] sg260;
  wire [1:0] sg261;
  wire [1:0] sg262;
  wire [1:0] sg263;
  wire [1:0] sg264;
  wire [1:0] sg265;
  wire [1:0] sg266;
  wire [1:0] sg267;
  wire [1:0] sg268;
  wire [1:0] sg269;
  wire [1:0] sg270;
  wire [1:0] sg271;
  wire [1:0] sg272;
  wire [1:0] sg273;
  wire [1:0] sg274;
  wire [1:0] sg275;
  wire [1:0] sg276;
  wire [1:0] sg277;
  wire [1:0] sg278;
  wire [1:0] sg279;
  wire [1:0] sg280;
  wire [1:0] sg281;
  wire [1:0] sg282;
  wire [1:0] sg283;
  wire [1:0] sg284;
  wire [1:0] sg285;
  wire [9:0] sg286;
  wire [1:0] sg289;
  wire [1:0] sg290;
  wire [1:0] sg291;
  wire [1:0] sg292;
  wire [1:0] sg293;
  wire [1:0] sg294;
  wire [1:0] sg295;
  wire [1:0] sg296;
  wire [1:0] sg297;
  wire [1:0] sg298;
  wire [1:0] sg299;
  wire [1:0] sg300;
  wire [1:0] sg301;
  wire [1:0] sg302;
  wire [1:0] sg303;
  wire [1:0] sg304;
  wire [1:0] sg305;
  wire [1:0] sg306;
  wire [1:0] sg307;
  wire [1:0] sg308;
  wire [1:0] sg309;
  wire [1:0] sg310;
  wire [1:0] sg311;
  wire [1:0] sg312;
  wire [1:0] sg313;
  wire [1:0] sg314;
  wire [1:0] sg315;
  wire [1:0] sg316;
  wire [1:0] sg317;
  wire [9:0] sg318;
  wire [1:0] sg321;
  wire [1:0] sg322;
  wire [1:0] sg323;
  wire [1:0] sg324;
  wire [1:0] sg325;
  wire [1:0] sg326;
  wire [1:0] sg327;
  wire [1:0] sg328;
  wire [1:0] sg329;
  wire [1:0] sg330;
  wire [1:0] sg331;
  wire [1:0] sg332;
  wire [1:0] sg333;
  wire [1:0] sg334;
  wire [1:0] sg335;
  wire [1:0] sg336;
  wire [1:0] sg337;
  wire [1:0] sg338;
  wire [1:0] sg339;
  wire [1:0] sg340;
  wire [1:0] sg341;
  wire [1:0] sg342;
  wire [1:0] sg343;
  wire [1:0] sg344;
  wire [1:0] sg345;
  wire [1:0] sg346;
  wire [1:0] sg347;
  wire [1:0] sg348;
  wire [1:0] sg349;
  wire [9:0] sg350;
  wire [1:0] sg353;
  wire [1:0] sg354;
  wire [1:0] sg355;
  wire [1:0] sg356;
  wire [1:0] sg357;
  wire [1:0] sg358;
  wire [1:0] sg359;
  wire [1:0] sg360;
  wire [1:0] sg361;
  wire [1:0] sg362;
  wire [1:0] sg363;
  wire [1:0] sg364;
  wire [1:0] sg365;
  wire [1:0] sg366;
  wire [1:0] sg367;
  wire [1:0] sg368;
  wire [1:0] sg369;
  wire [1:0] sg370;
  wire [1:0] sg371;
  wire [1:0] sg372;
  wire [1:0] sg373;
  wire [1:0] sg374;
  wire [1:0] sg375;
  wire [1:0] sg376;
  wire [1:0] sg377;
  wire [1:0] sg378;
  wire [1:0] sg379;
  wire [1:0] sg380;
  wire [1:0] sg381;
  wire [9:0] sg382;
  wire [1:0] sg385;
  wire [1:0] sg386;
  wire [1:0] sg387;
  wire [1:0] sg388;
  wire [1:0] sg389;
  wire [1:0] sg390;
  wire [1:0] sg391;
  wire [1:0] sg392;
  wire [1:0] sg393;
  wire [1:0] sg394;
  wire [1:0] sg395;
  wire [1:0] sg396;
  wire [1:0] sg397;
  wire [1:0] sg398;
  wire [1:0] sg399;
  wire [1:0] sg400;
  wire [1:0] sg401;
  wire [1:0] sg402;
  wire [1:0] sg403;
  wire [1:0] sg404;
  wire [1:0] sg405;
  wire [1:0] sg406;
  wire [1:0] sg407;
  wire [1:0] sg408;
  wire [1:0] sg409;
  wire [1:0] sg410;
  wire [1:0] sg411;
  wire [1:0] sg412;
  wire [1:0] sg413;
  wire [9:0] sg414;
  wire [1:0] sg417;
  wire [1:0] sg418;
  wire [1:0] sg419;
  wire [1:0] sg420;
  wire [1:0] sg421;
  wire [1:0] sg422;
  wire [1:0] sg423;
  wire [1:0] sg424;
  wire [1:0] sg425;
  wire [1:0] sg426;
  wire [1:0] sg427;
  wire [1:0] sg428;
  wire [1:0] sg429;
  wire [1:0] sg430;
  wire [1:0] sg431;
  wire [1:0] sg432;
  wire [1:0] sg433;
  wire [1:0] sg434;
  wire [1:0] sg435;
  wire [1:0] sg436;
  wire [1:0] sg437;
  wire [1:0] sg438;
  wire [1:0] sg439;
  wire [1:0] sg440;
  wire [1:0] sg441;
  wire [1:0] sg442;
  wire [1:0] sg443;
  wire [1:0] sg444;
  wire [1:0] sg445;
  wire [9:0] sg446;
  wire [1:0] sg449;
  wire [1:0] sg450;
  wire [1:0] sg451;
  wire [1:0] sg452;
  wire [1:0] sg453;
  wire [1:0] sg454;
  wire [1:0] sg455;
  wire [1:0] sg456;
  wire [1:0] sg457;
  wire [1:0] sg458;
  wire [1:0] sg459;
  wire [1:0] sg460;
  wire [1:0] sg461;
  wire [1:0] sg462;
  wire [1:0] sg463;
  wire [1:0] sg464;
  wire [1:0] sg465;
  wire [1:0] sg466;
  wire [1:0] sg467;
  wire [1:0] sg468;
  wire [1:0] sg469;
  wire [1:0] sg470;
  wire [1:0] sg471;
  wire [1:0] sg472;
  wire [1:0] sg473;
  wire [1:0] sg474;
  wire [1:0] sg475;
  wire [1:0] sg476;
  wire [1:0] sg477;
  wire [1:0] sg478;
  wire kanwa_s;
  wire _add_all_x_sig;
  wire [9:0] _add_all_x_start;
  wire [9:0] _add_all_x_goal;
  wire _add_all_x_dig_w;
  wire [9:0] _add_all_x_data_in33;
  wire [9:0] _add_all_x_data_in34;
  wire [9:0] _add_all_x_data_in35;
  wire [9:0] _add_all_x_data_in36;
  wire [9:0] _add_all_x_data_in37;
  wire [9:0] _add_all_x_data_in38;
  wire [9:0] _add_all_x_data_in39;
  wire [9:0] _add_all_x_data_in40;
  wire [9:0] _add_all_x_data_in41;
  wire [9:0] _add_all_x_data_in42;
  wire [9:0] _add_all_x_data_in43;
  wire [9:0] _add_all_x_data_in44;
  wire [9:0] _add_all_x_data_in45;
  wire [9:0] _add_all_x_data_in46;
  wire [9:0] _add_all_x_data_in47;
  wire [9:0] _add_all_x_data_in48;
  wire [9:0] _add_all_x_data_in49;
  wire [9:0] _add_all_x_data_in50;
  wire [9:0] _add_all_x_data_in51;
  wire [9:0] _add_all_x_data_in52;
  wire [9:0] _add_all_x_data_in53;
  wire [9:0] _add_all_x_data_in54;
  wire [9:0] _add_all_x_data_in55;
  wire [9:0] _add_all_x_data_in56;
  wire [9:0] _add_all_x_data_in57;
  wire [9:0] _add_all_x_data_in58;
  wire [9:0] _add_all_x_data_in59;
  wire [9:0] _add_all_x_data_in60;
  wire [9:0] _add_all_x_data_in61;
  wire [9:0] _add_all_x_data_in62;
  wire [9:0] _add_all_x_data_in65;
  wire [9:0] _add_all_x_data_in66;
  wire [9:0] _add_all_x_data_in67;
  wire [9:0] _add_all_x_data_in68;
  wire [9:0] _add_all_x_data_in69;
  wire [9:0] _add_all_x_data_in70;
  wire [9:0] _add_all_x_data_in71;
  wire [9:0] _add_all_x_data_in72;
  wire [9:0] _add_all_x_data_in73;
  wire [9:0] _add_all_x_data_in74;
  wire [9:0] _add_all_x_data_in75;
  wire [9:0] _add_all_x_data_in76;
  wire [9:0] _add_all_x_data_in77;
  wire [9:0] _add_all_x_data_in78;
  wire [9:0] _add_all_x_data_in79;
  wire [9:0] _add_all_x_data_in80;
  wire [9:0] _add_all_x_data_in81;
  wire [9:0] _add_all_x_data_in82;
  wire [9:0] _add_all_x_data_in83;
  wire [9:0] _add_all_x_data_in84;
  wire [9:0] _add_all_x_data_in85;
  wire [9:0] _add_all_x_data_in86;
  wire [9:0] _add_all_x_data_in87;
  wire [9:0] _add_all_x_data_in88;
  wire [9:0] _add_all_x_data_in89;
  wire [9:0] _add_all_x_data_in90;
  wire [9:0] _add_all_x_data_in91;
  wire [9:0] _add_all_x_data_in92;
  wire [9:0] _add_all_x_data_in93;
  wire [9:0] _add_all_x_data_in94;
  wire [9:0] _add_all_x_data_in97;
  wire [9:0] _add_all_x_data_in98;
  wire [9:0] _add_all_x_data_in99;
  wire [9:0] _add_all_x_data_in100;
  wire [9:0] _add_all_x_data_in101;
  wire [9:0] _add_all_x_data_in102;
  wire [9:0] _add_all_x_data_in103;
  wire [9:0] _add_all_x_data_in104;
  wire [9:0] _add_all_x_data_in105;
  wire [9:0] _add_all_x_data_in106;
  wire [9:0] _add_all_x_data_in107;
  wire [9:0] _add_all_x_data_in108;
  wire [9:0] _add_all_x_data_in109;
  wire [9:0] _add_all_x_data_in110;
  wire [9:0] _add_all_x_data_in111;
  wire [9:0] _add_all_x_data_in112;
  wire [9:0] _add_all_x_data_in113;
  wire [9:0] _add_all_x_data_in114;
  wire [9:0] _add_all_x_data_in115;
  wire [9:0] _add_all_x_data_in116;
  wire [9:0] _add_all_x_data_in117;
  wire [9:0] _add_all_x_data_in118;
  wire [9:0] _add_all_x_data_in119;
  wire [9:0] _add_all_x_data_in120;
  wire [9:0] _add_all_x_data_in121;
  wire [9:0] _add_all_x_data_in122;
  wire [9:0] _add_all_x_data_in123;
  wire [9:0] _add_all_x_data_in124;
  wire [9:0] _add_all_x_data_in125;
  wire [9:0] _add_all_x_data_in126;
  wire [9:0] _add_all_x_data_in129;
  wire [9:0] _add_all_x_data_in130;
  wire [9:0] _add_all_x_data_in131;
  wire [9:0] _add_all_x_data_in132;
  wire [9:0] _add_all_x_data_in133;
  wire [9:0] _add_all_x_data_in134;
  wire [9:0] _add_all_x_data_in135;
  wire [9:0] _add_all_x_data_in136;
  wire [9:0] _add_all_x_data_in137;
  wire [9:0] _add_all_x_data_in138;
  wire [9:0] _add_all_x_data_in139;
  wire [9:0] _add_all_x_data_in140;
  wire [9:0] _add_all_x_data_in141;
  wire [9:0] _add_all_x_data_in142;
  wire [9:0] _add_all_x_data_in143;
  wire [9:0] _add_all_x_data_in144;
  wire [9:0] _add_all_x_data_in145;
  wire [9:0] _add_all_x_data_in146;
  wire [9:0] _add_all_x_data_in147;
  wire [9:0] _add_all_x_data_in148;
  wire [9:0] _add_all_x_data_in149;
  wire [9:0] _add_all_x_data_in150;
  wire [9:0] _add_all_x_data_in151;
  wire [9:0] _add_all_x_data_in152;
  wire [9:0] _add_all_x_data_in153;
  wire [9:0] _add_all_x_data_in154;
  wire [9:0] _add_all_x_data_in155;
  wire [9:0] _add_all_x_data_in156;
  wire [9:0] _add_all_x_data_in157;
  wire [9:0] _add_all_x_data_in158;
  wire [9:0] _add_all_x_data_in161;
  wire [9:0] _add_all_x_data_in162;
  wire [9:0] _add_all_x_data_in163;
  wire [9:0] _add_all_x_data_in164;
  wire [9:0] _add_all_x_data_in165;
  wire [9:0] _add_all_x_data_in166;
  wire [9:0] _add_all_x_data_in167;
  wire [9:0] _add_all_x_data_in168;
  wire [9:0] _add_all_x_data_in169;
  wire [9:0] _add_all_x_data_in170;
  wire [9:0] _add_all_x_data_in171;
  wire [9:0] _add_all_x_data_in172;
  wire [9:0] _add_all_x_data_in173;
  wire [9:0] _add_all_x_data_in174;
  wire [9:0] _add_all_x_data_in175;
  wire [9:0] _add_all_x_data_in176;
  wire [9:0] _add_all_x_data_in177;
  wire [9:0] _add_all_x_data_in178;
  wire [9:0] _add_all_x_data_in179;
  wire [9:0] _add_all_x_data_in180;
  wire [9:0] _add_all_x_data_in181;
  wire [9:0] _add_all_x_data_in182;
  wire [9:0] _add_all_x_data_in183;
  wire [9:0] _add_all_x_data_in184;
  wire [9:0] _add_all_x_data_in185;
  wire [9:0] _add_all_x_data_in186;
  wire [9:0] _add_all_x_data_in187;
  wire [9:0] _add_all_x_data_in188;
  wire [9:0] _add_all_x_data_in189;
  wire [9:0] _add_all_x_data_in190;
  wire [9:0] _add_all_x_data_in193;
  wire [9:0] _add_all_x_data_in194;
  wire [9:0] _add_all_x_data_in195;
  wire [9:0] _add_all_x_data_in196;
  wire [9:0] _add_all_x_data_in197;
  wire [9:0] _add_all_x_data_in198;
  wire [9:0] _add_all_x_data_in199;
  wire [9:0] _add_all_x_data_in200;
  wire [9:0] _add_all_x_data_in201;
  wire [9:0] _add_all_x_data_in202;
  wire [9:0] _add_all_x_data_in203;
  wire [9:0] _add_all_x_data_in204;
  wire [9:0] _add_all_x_data_in205;
  wire [9:0] _add_all_x_data_in206;
  wire [9:0] _add_all_x_data_in207;
  wire [9:0] _add_all_x_data_in208;
  wire [9:0] _add_all_x_data_in209;
  wire [9:0] _add_all_x_data_in210;
  wire [9:0] _add_all_x_data_in211;
  wire [9:0] _add_all_x_data_in212;
  wire [9:0] _add_all_x_data_in213;
  wire [9:0] _add_all_x_data_in214;
  wire [9:0] _add_all_x_data_in215;
  wire [9:0] _add_all_x_data_in216;
  wire [9:0] _add_all_x_data_in217;
  wire [9:0] _add_all_x_data_in218;
  wire [9:0] _add_all_x_data_in219;
  wire [9:0] _add_all_x_data_in220;
  wire [9:0] _add_all_x_data_in221;
  wire [9:0] _add_all_x_data_in222;
  wire [9:0] _add_all_x_data_in225;
  wire [9:0] _add_all_x_data_in226;
  wire [9:0] _add_all_x_data_in227;
  wire [9:0] _add_all_x_data_in228;
  wire [9:0] _add_all_x_data_in229;
  wire [9:0] _add_all_x_data_in230;
  wire [9:0] _add_all_x_data_in231;
  wire [9:0] _add_all_x_data_in232;
  wire [9:0] _add_all_x_data_in233;
  wire [9:0] _add_all_x_data_in234;
  wire [9:0] _add_all_x_data_in235;
  wire [9:0] _add_all_x_data_in236;
  wire [9:0] _add_all_x_data_in237;
  wire [9:0] _add_all_x_data_in238;
  wire [9:0] _add_all_x_data_in239;
  wire [9:0] _add_all_x_data_in240;
  wire [9:0] _add_all_x_data_in241;
  wire [9:0] _add_all_x_data_in242;
  wire [9:0] _add_all_x_data_in243;
  wire [9:0] _add_all_x_data_in244;
  wire [9:0] _add_all_x_data_in245;
  wire [9:0] _add_all_x_data_in246;
  wire [9:0] _add_all_x_data_in247;
  wire [9:0] _add_all_x_data_in248;
  wire [9:0] _add_all_x_data_in249;
  wire [9:0] _add_all_x_data_in250;
  wire [9:0] _add_all_x_data_in251;
  wire [9:0] _add_all_x_data_in252;
  wire [9:0] _add_all_x_data_in253;
  wire [9:0] _add_all_x_data_in254;
  wire [9:0] _add_all_x_data_in257;
  wire [9:0] _add_all_x_data_in258;
  wire [9:0] _add_all_x_data_in259;
  wire [9:0] _add_all_x_data_in260;
  wire [9:0] _add_all_x_data_in261;
  wire [9:0] _add_all_x_data_in262;
  wire [9:0] _add_all_x_data_in263;
  wire [9:0] _add_all_x_data_in264;
  wire [9:0] _add_all_x_data_in265;
  wire [9:0] _add_all_x_data_in266;
  wire [9:0] _add_all_x_data_in267;
  wire [9:0] _add_all_x_data_in268;
  wire [9:0] _add_all_x_data_in269;
  wire [9:0] _add_all_x_data_in270;
  wire [9:0] _add_all_x_data_in271;
  wire [9:0] _add_all_x_data_in272;
  wire [9:0] _add_all_x_data_in273;
  wire [9:0] _add_all_x_data_in274;
  wire [9:0] _add_all_x_data_in275;
  wire [9:0] _add_all_x_data_in276;
  wire [9:0] _add_all_x_data_in277;
  wire [9:0] _add_all_x_data_in278;
  wire [9:0] _add_all_x_data_in279;
  wire [9:0] _add_all_x_data_in280;
  wire [9:0] _add_all_x_data_in281;
  wire [9:0] _add_all_x_data_in282;
  wire [9:0] _add_all_x_data_in283;
  wire [9:0] _add_all_x_data_in284;
  wire [9:0] _add_all_x_data_in285;
  wire [9:0] _add_all_x_data_in286;
  wire [9:0] _add_all_x_data_in289;
  wire [9:0] _add_all_x_data_in290;
  wire [9:0] _add_all_x_data_in291;
  wire [9:0] _add_all_x_data_in292;
  wire [9:0] _add_all_x_data_in293;
  wire [9:0] _add_all_x_data_in294;
  wire [9:0] _add_all_x_data_in295;
  wire [9:0] _add_all_x_data_in296;
  wire [9:0] _add_all_x_data_in297;
  wire [9:0] _add_all_x_data_in298;
  wire [9:0] _add_all_x_data_in299;
  wire [9:0] _add_all_x_data_in300;
  wire [9:0] _add_all_x_data_in301;
  wire [9:0] _add_all_x_data_in302;
  wire [9:0] _add_all_x_data_in303;
  wire [9:0] _add_all_x_data_in304;
  wire [9:0] _add_all_x_data_in305;
  wire [9:0] _add_all_x_data_in306;
  wire [9:0] _add_all_x_data_in307;
  wire [9:0] _add_all_x_data_in308;
  wire [9:0] _add_all_x_data_in309;
  wire [9:0] _add_all_x_data_in310;
  wire [9:0] _add_all_x_data_in311;
  wire [9:0] _add_all_x_data_in312;
  wire [9:0] _add_all_x_data_in313;
  wire [9:0] _add_all_x_data_in314;
  wire [9:0] _add_all_x_data_in315;
  wire [9:0] _add_all_x_data_in316;
  wire [9:0] _add_all_x_data_in317;
  wire [9:0] _add_all_x_data_in318;
  wire [9:0] _add_all_x_data_in321;
  wire [9:0] _add_all_x_data_in322;
  wire [9:0] _add_all_x_data_in323;
  wire [9:0] _add_all_x_data_in324;
  wire [9:0] _add_all_x_data_in325;
  wire [9:0] _add_all_x_data_in326;
  wire [9:0] _add_all_x_data_in327;
  wire [9:0] _add_all_x_data_in328;
  wire [9:0] _add_all_x_data_in329;
  wire [9:0] _add_all_x_data_in330;
  wire [9:0] _add_all_x_data_in331;
  wire [9:0] _add_all_x_data_in332;
  wire [9:0] _add_all_x_data_in333;
  wire [9:0] _add_all_x_data_in334;
  wire [9:0] _add_all_x_data_in335;
  wire [9:0] _add_all_x_data_in336;
  wire [9:0] _add_all_x_data_in337;
  wire [9:0] _add_all_x_data_in338;
  wire [9:0] _add_all_x_data_in339;
  wire [9:0] _add_all_x_data_in340;
  wire [9:0] _add_all_x_data_in341;
  wire [9:0] _add_all_x_data_in342;
  wire [9:0] _add_all_x_data_in343;
  wire [9:0] _add_all_x_data_in344;
  wire [9:0] _add_all_x_data_in345;
  wire [9:0] _add_all_x_data_in346;
  wire [9:0] _add_all_x_data_in347;
  wire [9:0] _add_all_x_data_in348;
  wire [9:0] _add_all_x_data_in349;
  wire [9:0] _add_all_x_data_in350;
  wire [9:0] _add_all_x_data_in353;
  wire [9:0] _add_all_x_data_in354;
  wire [9:0] _add_all_x_data_in355;
  wire [9:0] _add_all_x_data_in356;
  wire [9:0] _add_all_x_data_in357;
  wire [9:0] _add_all_x_data_in358;
  wire [9:0] _add_all_x_data_in359;
  wire [9:0] _add_all_x_data_in360;
  wire [9:0] _add_all_x_data_in361;
  wire [9:0] _add_all_x_data_in362;
  wire [9:0] _add_all_x_data_in363;
  wire [9:0] _add_all_x_data_in364;
  wire [9:0] _add_all_x_data_in365;
  wire [9:0] _add_all_x_data_in366;
  wire [9:0] _add_all_x_data_in367;
  wire [9:0] _add_all_x_data_in368;
  wire [9:0] _add_all_x_data_in369;
  wire [9:0] _add_all_x_data_in370;
  wire [9:0] _add_all_x_data_in371;
  wire [9:0] _add_all_x_data_in372;
  wire [9:0] _add_all_x_data_in373;
  wire [9:0] _add_all_x_data_in374;
  wire [9:0] _add_all_x_data_in375;
  wire [9:0] _add_all_x_data_in376;
  wire [9:0] _add_all_x_data_in377;
  wire [9:0] _add_all_x_data_in378;
  wire [9:0] _add_all_x_data_in379;
  wire [9:0] _add_all_x_data_in380;
  wire [9:0] _add_all_x_data_in381;
  wire [9:0] _add_all_x_data_in382;
  wire [9:0] _add_all_x_data_in385;
  wire [9:0] _add_all_x_data_in386;
  wire [9:0] _add_all_x_data_in387;
  wire [9:0] _add_all_x_data_in388;
  wire [9:0] _add_all_x_data_in389;
  wire [9:0] _add_all_x_data_in390;
  wire [9:0] _add_all_x_data_in391;
  wire [9:0] _add_all_x_data_in392;
  wire [9:0] _add_all_x_data_in393;
  wire [9:0] _add_all_x_data_in394;
  wire [9:0] _add_all_x_data_in395;
  wire [9:0] _add_all_x_data_in396;
  wire [9:0] _add_all_x_data_in397;
  wire [9:0] _add_all_x_data_in398;
  wire [9:0] _add_all_x_data_in399;
  wire [9:0] _add_all_x_data_in400;
  wire [9:0] _add_all_x_data_in401;
  wire [9:0] _add_all_x_data_in402;
  wire [9:0] _add_all_x_data_in403;
  wire [9:0] _add_all_x_data_in404;
  wire [9:0] _add_all_x_data_in405;
  wire [9:0] _add_all_x_data_in406;
  wire [9:0] _add_all_x_data_in407;
  wire [9:0] _add_all_x_data_in408;
  wire [9:0] _add_all_x_data_in409;
  wire [9:0] _add_all_x_data_in410;
  wire [9:0] _add_all_x_data_in411;
  wire [9:0] _add_all_x_data_in412;
  wire [9:0] _add_all_x_data_in413;
  wire [9:0] _add_all_x_data_in414;
  wire [9:0] _add_all_x_data_in417;
  wire [9:0] _add_all_x_data_in418;
  wire [9:0] _add_all_x_data_in419;
  wire [9:0] _add_all_x_data_in420;
  wire [9:0] _add_all_x_data_in421;
  wire [9:0] _add_all_x_data_in422;
  wire [9:0] _add_all_x_data_in423;
  wire [9:0] _add_all_x_data_in424;
  wire [9:0] _add_all_x_data_in425;
  wire [9:0] _add_all_x_data_in426;
  wire [9:0] _add_all_x_data_in427;
  wire [9:0] _add_all_x_data_in428;
  wire [9:0] _add_all_x_data_in429;
  wire [9:0] _add_all_x_data_in430;
  wire [9:0] _add_all_x_data_in431;
  wire [9:0] _add_all_x_data_in432;
  wire [9:0] _add_all_x_data_in433;
  wire [9:0] _add_all_x_data_in434;
  wire [9:0] _add_all_x_data_in435;
  wire [9:0] _add_all_x_data_in436;
  wire [9:0] _add_all_x_data_in437;
  wire [9:0] _add_all_x_data_in438;
  wire [9:0] _add_all_x_data_in439;
  wire [9:0] _add_all_x_data_in440;
  wire [9:0] _add_all_x_data_in441;
  wire [9:0] _add_all_x_data_in442;
  wire [9:0] _add_all_x_data_in443;
  wire [9:0] _add_all_x_data_in444;
  wire [9:0] _add_all_x_data_in445;
  wire [9:0] _add_all_x_data_in446;
  wire [9:0] _add_all_x_data_in449;
  wire [9:0] _add_all_x_data_in450;
  wire [9:0] _add_all_x_data_in451;
  wire [9:0] _add_all_x_data_in452;
  wire [9:0] _add_all_x_data_in453;
  wire [9:0] _add_all_x_data_in454;
  wire [9:0] _add_all_x_data_in455;
  wire [9:0] _add_all_x_data_in456;
  wire [9:0] _add_all_x_data_in457;
  wire [9:0] _add_all_x_data_in458;
  wire [9:0] _add_all_x_data_in459;
  wire [9:0] _add_all_x_data_in460;
  wire [9:0] _add_all_x_data_in461;
  wire [9:0] _add_all_x_data_in462;
  wire [9:0] _add_all_x_data_in463;
  wire [9:0] _add_all_x_data_in464;
  wire [9:0] _add_all_x_data_in465;
  wire [9:0] _add_all_x_data_in466;
  wire [9:0] _add_all_x_data_in467;
  wire [9:0] _add_all_x_data_in468;
  wire [9:0] _add_all_x_data_in469;
  wire [9:0] _add_all_x_data_in470;
  wire [9:0] _add_all_x_data_in471;
  wire [9:0] _add_all_x_data_in472;
  wire [9:0] _add_all_x_data_in473;
  wire [9:0] _add_all_x_data_in474;
  wire [9:0] _add_all_x_data_in475;
  wire [9:0] _add_all_x_data_in476;
  wire [9:0] _add_all_x_data_in477;
  wire [9:0] _add_all_x_data_in478;
  wire [9:0] _add_all_x_data_out_org33;
  wire [9:0] _add_all_x_data_out_org34;
  wire [9:0] _add_all_x_data_out_org35;
  wire [9:0] _add_all_x_data_out_org36;
  wire [9:0] _add_all_x_data_out_org37;
  wire [9:0] _add_all_x_data_out_org38;
  wire [9:0] _add_all_x_data_out_org39;
  wire [9:0] _add_all_x_data_out_org40;
  wire [9:0] _add_all_x_data_out_org41;
  wire [9:0] _add_all_x_data_out_org42;
  wire [9:0] _add_all_x_data_out_org43;
  wire [9:0] _add_all_x_data_out_org44;
  wire [9:0] _add_all_x_data_out_org45;
  wire [9:0] _add_all_x_data_out_org46;
  wire [9:0] _add_all_x_data_out_org47;
  wire [9:0] _add_all_x_data_out_org48;
  wire [9:0] _add_all_x_data_out_org49;
  wire [9:0] _add_all_x_data_out_org50;
  wire [9:0] _add_all_x_data_out_org51;
  wire [9:0] _add_all_x_data_out_org52;
  wire [9:0] _add_all_x_data_out_org53;
  wire [9:0] _add_all_x_data_out_org54;
  wire [9:0] _add_all_x_data_out_org55;
  wire [9:0] _add_all_x_data_out_org56;
  wire [9:0] _add_all_x_data_out_org57;
  wire [9:0] _add_all_x_data_out_org58;
  wire [9:0] _add_all_x_data_out_org59;
  wire [9:0] _add_all_x_data_out_org60;
  wire [9:0] _add_all_x_data_out_org61;
  wire [9:0] _add_all_x_data_out_org62;
  wire [9:0] _add_all_x_data_out_org65;
  wire [9:0] _add_all_x_data_out_org66;
  wire [9:0] _add_all_x_data_out_org67;
  wire [9:0] _add_all_x_data_out_org68;
  wire [9:0] _add_all_x_data_out_org69;
  wire [9:0] _add_all_x_data_out_org70;
  wire [9:0] _add_all_x_data_out_org71;
  wire [9:0] _add_all_x_data_out_org72;
  wire [9:0] _add_all_x_data_out_org73;
  wire [9:0] _add_all_x_data_out_org74;
  wire [9:0] _add_all_x_data_out_org75;
  wire [9:0] _add_all_x_data_out_org76;
  wire [9:0] _add_all_x_data_out_org77;
  wire [9:0] _add_all_x_data_out_org78;
  wire [9:0] _add_all_x_data_out_org79;
  wire [9:0] _add_all_x_data_out_org80;
  wire [9:0] _add_all_x_data_out_org81;
  wire [9:0] _add_all_x_data_out_org82;
  wire [9:0] _add_all_x_data_out_org83;
  wire [9:0] _add_all_x_data_out_org84;
  wire [9:0] _add_all_x_data_out_org85;
  wire [9:0] _add_all_x_data_out_org86;
  wire [9:0] _add_all_x_data_out_org87;
  wire [9:0] _add_all_x_data_out_org88;
  wire [9:0] _add_all_x_data_out_org89;
  wire [9:0] _add_all_x_data_out_org90;
  wire [9:0] _add_all_x_data_out_org91;
  wire [9:0] _add_all_x_data_out_org92;
  wire [9:0] _add_all_x_data_out_org93;
  wire [9:0] _add_all_x_data_out_org94;
  wire [9:0] _add_all_x_data_out_org97;
  wire [9:0] _add_all_x_data_out_org98;
  wire [9:0] _add_all_x_data_out_org99;
  wire [9:0] _add_all_x_data_out_org100;
  wire [9:0] _add_all_x_data_out_org101;
  wire [9:0] _add_all_x_data_out_org102;
  wire [9:0] _add_all_x_data_out_org103;
  wire [9:0] _add_all_x_data_out_org104;
  wire [9:0] _add_all_x_data_out_org105;
  wire [9:0] _add_all_x_data_out_org106;
  wire [9:0] _add_all_x_data_out_org107;
  wire [9:0] _add_all_x_data_out_org108;
  wire [9:0] _add_all_x_data_out_org109;
  wire [9:0] _add_all_x_data_out_org110;
  wire [9:0] _add_all_x_data_out_org111;
  wire [9:0] _add_all_x_data_out_org112;
  wire [9:0] _add_all_x_data_out_org113;
  wire [9:0] _add_all_x_data_out_org114;
  wire [9:0] _add_all_x_data_out_org115;
  wire [9:0] _add_all_x_data_out_org116;
  wire [9:0] _add_all_x_data_out_org117;
  wire [9:0] _add_all_x_data_out_org118;
  wire [9:0] _add_all_x_data_out_org119;
  wire [9:0] _add_all_x_data_out_org120;
  wire [9:0] _add_all_x_data_out_org121;
  wire [9:0] _add_all_x_data_out_org122;
  wire [9:0] _add_all_x_data_out_org123;
  wire [9:0] _add_all_x_data_out_org124;
  wire [9:0] _add_all_x_data_out_org125;
  wire [9:0] _add_all_x_data_out_org126;
  wire [9:0] _add_all_x_data_out_org129;
  wire [9:0] _add_all_x_data_out_org130;
  wire [9:0] _add_all_x_data_out_org131;
  wire [9:0] _add_all_x_data_out_org132;
  wire [9:0] _add_all_x_data_out_org133;
  wire [9:0] _add_all_x_data_out_org134;
  wire [9:0] _add_all_x_data_out_org135;
  wire [9:0] _add_all_x_data_out_org136;
  wire [9:0] _add_all_x_data_out_org137;
  wire [9:0] _add_all_x_data_out_org138;
  wire [9:0] _add_all_x_data_out_org139;
  wire [9:0] _add_all_x_data_out_org140;
  wire [9:0] _add_all_x_data_out_org141;
  wire [9:0] _add_all_x_data_out_org142;
  wire [9:0] _add_all_x_data_out_org143;
  wire [9:0] _add_all_x_data_out_org144;
  wire [9:0] _add_all_x_data_out_org145;
  wire [9:0] _add_all_x_data_out_org146;
  wire [9:0] _add_all_x_data_out_org147;
  wire [9:0] _add_all_x_data_out_org148;
  wire [9:0] _add_all_x_data_out_org149;
  wire [9:0] _add_all_x_data_out_org150;
  wire [9:0] _add_all_x_data_out_org151;
  wire [9:0] _add_all_x_data_out_org152;
  wire [9:0] _add_all_x_data_out_org153;
  wire [9:0] _add_all_x_data_out_org154;
  wire [9:0] _add_all_x_data_out_org155;
  wire [9:0] _add_all_x_data_out_org156;
  wire [9:0] _add_all_x_data_out_org157;
  wire [9:0] _add_all_x_data_out_org158;
  wire [9:0] _add_all_x_data_out_org161;
  wire [9:0] _add_all_x_data_out_org162;
  wire [9:0] _add_all_x_data_out_org163;
  wire [9:0] _add_all_x_data_out_org164;
  wire [9:0] _add_all_x_data_out_org165;
  wire [9:0] _add_all_x_data_out_org166;
  wire [9:0] _add_all_x_data_out_org167;
  wire [9:0] _add_all_x_data_out_org168;
  wire [9:0] _add_all_x_data_out_org169;
  wire [9:0] _add_all_x_data_out_org170;
  wire [9:0] _add_all_x_data_out_org171;
  wire [9:0] _add_all_x_data_out_org172;
  wire [9:0] _add_all_x_data_out_org173;
  wire [9:0] _add_all_x_data_out_org174;
  wire [9:0] _add_all_x_data_out_org175;
  wire [9:0] _add_all_x_data_out_org176;
  wire [9:0] _add_all_x_data_out_org177;
  wire [9:0] _add_all_x_data_out_org178;
  wire [9:0] _add_all_x_data_out_org179;
  wire [9:0] _add_all_x_data_out_org180;
  wire [9:0] _add_all_x_data_out_org181;
  wire [9:0] _add_all_x_data_out_org182;
  wire [9:0] _add_all_x_data_out_org183;
  wire [9:0] _add_all_x_data_out_org184;
  wire [9:0] _add_all_x_data_out_org185;
  wire [9:0] _add_all_x_data_out_org186;
  wire [9:0] _add_all_x_data_out_org187;
  wire [9:0] _add_all_x_data_out_org188;
  wire [9:0] _add_all_x_data_out_org189;
  wire [9:0] _add_all_x_data_out_org190;
  wire [9:0] _add_all_x_data_out_org193;
  wire [9:0] _add_all_x_data_out_org194;
  wire [9:0] _add_all_x_data_out_org195;
  wire [9:0] _add_all_x_data_out_org196;
  wire [9:0] _add_all_x_data_out_org197;
  wire [9:0] _add_all_x_data_out_org198;
  wire [9:0] _add_all_x_data_out_org199;
  wire [9:0] _add_all_x_data_out_org200;
  wire [9:0] _add_all_x_data_out_org201;
  wire [9:0] _add_all_x_data_out_org202;
  wire [9:0] _add_all_x_data_out_org203;
  wire [9:0] _add_all_x_data_out_org204;
  wire [9:0] _add_all_x_data_out_org205;
  wire [9:0] _add_all_x_data_out_org206;
  wire [9:0] _add_all_x_data_out_org207;
  wire [9:0] _add_all_x_data_out_org208;
  wire [9:0] _add_all_x_data_out_org209;
  wire [9:0] _add_all_x_data_out_org210;
  wire [9:0] _add_all_x_data_out_org211;
  wire [9:0] _add_all_x_data_out_org212;
  wire [9:0] _add_all_x_data_out_org213;
  wire [9:0] _add_all_x_data_out_org214;
  wire [9:0] _add_all_x_data_out_org215;
  wire [9:0] _add_all_x_data_out_org216;
  wire [9:0] _add_all_x_data_out_org217;
  wire [9:0] _add_all_x_data_out_org218;
  wire [9:0] _add_all_x_data_out_org219;
  wire [9:0] _add_all_x_data_out_org220;
  wire [9:0] _add_all_x_data_out_org221;
  wire [9:0] _add_all_x_data_out_org222;
  wire [9:0] _add_all_x_data_out_org225;
  wire [9:0] _add_all_x_data_out_org226;
  wire [9:0] _add_all_x_data_out_org227;
  wire [9:0] _add_all_x_data_out_org228;
  wire [9:0] _add_all_x_data_out_org229;
  wire [9:0] _add_all_x_data_out_org230;
  wire [9:0] _add_all_x_data_out_org231;
  wire [9:0] _add_all_x_data_out_org232;
  wire [9:0] _add_all_x_data_out_org233;
  wire [9:0] _add_all_x_data_out_org234;
  wire [9:0] _add_all_x_data_out_org235;
  wire [9:0] _add_all_x_data_out_org236;
  wire [9:0] _add_all_x_data_out_org237;
  wire [9:0] _add_all_x_data_out_org238;
  wire [9:0] _add_all_x_data_out_org239;
  wire [9:0] _add_all_x_data_out_org240;
  wire [9:0] _add_all_x_data_out_org241;
  wire [9:0] _add_all_x_data_out_org242;
  wire [9:0] _add_all_x_data_out_org243;
  wire [9:0] _add_all_x_data_out_org244;
  wire [9:0] _add_all_x_data_out_org245;
  wire [9:0] _add_all_x_data_out_org246;
  wire [9:0] _add_all_x_data_out_org247;
  wire [9:0] _add_all_x_data_out_org248;
  wire [9:0] _add_all_x_data_out_org249;
  wire [9:0] _add_all_x_data_out_org250;
  wire [9:0] _add_all_x_data_out_org251;
  wire [9:0] _add_all_x_data_out_org252;
  wire [9:0] _add_all_x_data_out_org253;
  wire [9:0] _add_all_x_data_out_org254;
  wire [9:0] _add_all_x_data_out_org257;
  wire [9:0] _add_all_x_data_out_org258;
  wire [9:0] _add_all_x_data_out_org259;
  wire [9:0] _add_all_x_data_out_org260;
  wire [9:0] _add_all_x_data_out_org261;
  wire [9:0] _add_all_x_data_out_org262;
  wire [9:0] _add_all_x_data_out_org263;
  wire [9:0] _add_all_x_data_out_org264;
  wire [9:0] _add_all_x_data_out_org265;
  wire [9:0] _add_all_x_data_out_org266;
  wire [9:0] _add_all_x_data_out_org267;
  wire [9:0] _add_all_x_data_out_org268;
  wire [9:0] _add_all_x_data_out_org269;
  wire [9:0] _add_all_x_data_out_org270;
  wire [9:0] _add_all_x_data_out_org271;
  wire [9:0] _add_all_x_data_out_org272;
  wire [9:0] _add_all_x_data_out_org273;
  wire [9:0] _add_all_x_data_out_org274;
  wire [9:0] _add_all_x_data_out_org275;
  wire [9:0] _add_all_x_data_out_org276;
  wire [9:0] _add_all_x_data_out_org277;
  wire [9:0] _add_all_x_data_out_org278;
  wire [9:0] _add_all_x_data_out_org279;
  wire [9:0] _add_all_x_data_out_org280;
  wire [9:0] _add_all_x_data_out_org281;
  wire [9:0] _add_all_x_data_out_org282;
  wire [9:0] _add_all_x_data_out_org283;
  wire [9:0] _add_all_x_data_out_org284;
  wire [9:0] _add_all_x_data_out_org285;
  wire [9:0] _add_all_x_data_out_org286;
  wire [9:0] _add_all_x_data_out_org289;
  wire [9:0] _add_all_x_data_out_org290;
  wire [9:0] _add_all_x_data_out_org291;
  wire [9:0] _add_all_x_data_out_org292;
  wire [9:0] _add_all_x_data_out_org293;
  wire [9:0] _add_all_x_data_out_org294;
  wire [9:0] _add_all_x_data_out_org295;
  wire [9:0] _add_all_x_data_out_org296;
  wire [9:0] _add_all_x_data_out_org297;
  wire [9:0] _add_all_x_data_out_org298;
  wire [9:0] _add_all_x_data_out_org299;
  wire [9:0] _add_all_x_data_out_org300;
  wire [9:0] _add_all_x_data_out_org301;
  wire [9:0] _add_all_x_data_out_org302;
  wire [9:0] _add_all_x_data_out_org303;
  wire [9:0] _add_all_x_data_out_org304;
  wire [9:0] _add_all_x_data_out_org305;
  wire [9:0] _add_all_x_data_out_org306;
  wire [9:0] _add_all_x_data_out_org307;
  wire [9:0] _add_all_x_data_out_org308;
  wire [9:0] _add_all_x_data_out_org309;
  wire [9:0] _add_all_x_data_out_org310;
  wire [9:0] _add_all_x_data_out_org311;
  wire [9:0] _add_all_x_data_out_org312;
  wire [9:0] _add_all_x_data_out_org313;
  wire [9:0] _add_all_x_data_out_org314;
  wire [9:0] _add_all_x_data_out_org315;
  wire [9:0] _add_all_x_data_out_org316;
  wire [9:0] _add_all_x_data_out_org317;
  wire [9:0] _add_all_x_data_out_org318;
  wire [9:0] _add_all_x_data_out_org321;
  wire [9:0] _add_all_x_data_out_org322;
  wire [9:0] _add_all_x_data_out_org323;
  wire [9:0] _add_all_x_data_out_org324;
  wire [9:0] _add_all_x_data_out_org325;
  wire [9:0] _add_all_x_data_out_org326;
  wire [9:0] _add_all_x_data_out_org327;
  wire [9:0] _add_all_x_data_out_org328;
  wire [9:0] _add_all_x_data_out_org329;
  wire [9:0] _add_all_x_data_out_org330;
  wire [9:0] _add_all_x_data_out_org331;
  wire [9:0] _add_all_x_data_out_org332;
  wire [9:0] _add_all_x_data_out_org333;
  wire [9:0] _add_all_x_data_out_org334;
  wire [9:0] _add_all_x_data_out_org335;
  wire [9:0] _add_all_x_data_out_org336;
  wire [9:0] _add_all_x_data_out_org337;
  wire [9:0] _add_all_x_data_out_org338;
  wire [9:0] _add_all_x_data_out_org339;
  wire [9:0] _add_all_x_data_out_org340;
  wire [9:0] _add_all_x_data_out_org341;
  wire [9:0] _add_all_x_data_out_org342;
  wire [9:0] _add_all_x_data_out_org343;
  wire [9:0] _add_all_x_data_out_org344;
  wire [9:0] _add_all_x_data_out_org345;
  wire [9:0] _add_all_x_data_out_org346;
  wire [9:0] _add_all_x_data_out_org347;
  wire [9:0] _add_all_x_data_out_org348;
  wire [9:0] _add_all_x_data_out_org349;
  wire [9:0] _add_all_x_data_out_org350;
  wire [9:0] _add_all_x_data_out_org353;
  wire [9:0] _add_all_x_data_out_org354;
  wire [9:0] _add_all_x_data_out_org355;
  wire [9:0] _add_all_x_data_out_org356;
  wire [9:0] _add_all_x_data_out_org357;
  wire [9:0] _add_all_x_data_out_org358;
  wire [9:0] _add_all_x_data_out_org359;
  wire [9:0] _add_all_x_data_out_org360;
  wire [9:0] _add_all_x_data_out_org361;
  wire [9:0] _add_all_x_data_out_org362;
  wire [9:0] _add_all_x_data_out_org363;
  wire [9:0] _add_all_x_data_out_org364;
  wire [9:0] _add_all_x_data_out_org365;
  wire [9:0] _add_all_x_data_out_org366;
  wire [9:0] _add_all_x_data_out_org367;
  wire [9:0] _add_all_x_data_out_org368;
  wire [9:0] _add_all_x_data_out_org369;
  wire [9:0] _add_all_x_data_out_org370;
  wire [9:0] _add_all_x_data_out_org371;
  wire [9:0] _add_all_x_data_out_org372;
  wire [9:0] _add_all_x_data_out_org373;
  wire [9:0] _add_all_x_data_out_org374;
  wire [9:0] _add_all_x_data_out_org375;
  wire [9:0] _add_all_x_data_out_org376;
  wire [9:0] _add_all_x_data_out_org377;
  wire [9:0] _add_all_x_data_out_org378;
  wire [9:0] _add_all_x_data_out_org379;
  wire [9:0] _add_all_x_data_out_org380;
  wire [9:0] _add_all_x_data_out_org381;
  wire [9:0] _add_all_x_data_out_org382;
  wire [9:0] _add_all_x_data_out_org385;
  wire [9:0] _add_all_x_data_out_org386;
  wire [9:0] _add_all_x_data_out_org387;
  wire [9:0] _add_all_x_data_out_org388;
  wire [9:0] _add_all_x_data_out_org389;
  wire [9:0] _add_all_x_data_out_org390;
  wire [9:0] _add_all_x_data_out_org391;
  wire [9:0] _add_all_x_data_out_org392;
  wire [9:0] _add_all_x_data_out_org393;
  wire [9:0] _add_all_x_data_out_org394;
  wire [9:0] _add_all_x_data_out_org395;
  wire [9:0] _add_all_x_data_out_org396;
  wire [9:0] _add_all_x_data_out_org397;
  wire [9:0] _add_all_x_data_out_org398;
  wire [9:0] _add_all_x_data_out_org399;
  wire [9:0] _add_all_x_data_out_org400;
  wire [9:0] _add_all_x_data_out_org401;
  wire [9:0] _add_all_x_data_out_org402;
  wire [9:0] _add_all_x_data_out_org403;
  wire [9:0] _add_all_x_data_out_org404;
  wire [9:0] _add_all_x_data_out_org405;
  wire [9:0] _add_all_x_data_out_org406;
  wire [9:0] _add_all_x_data_out_org407;
  wire [9:0] _add_all_x_data_out_org408;
  wire [9:0] _add_all_x_data_out_org409;
  wire [9:0] _add_all_x_data_out_org410;
  wire [9:0] _add_all_x_data_out_org411;
  wire [9:0] _add_all_x_data_out_org412;
  wire [9:0] _add_all_x_data_out_org413;
  wire [9:0] _add_all_x_data_out_org414;
  wire [9:0] _add_all_x_data_out_org417;
  wire [9:0] _add_all_x_data_out_org418;
  wire [9:0] _add_all_x_data_out_org419;
  wire [9:0] _add_all_x_data_out_org420;
  wire [9:0] _add_all_x_data_out_org421;
  wire [9:0] _add_all_x_data_out_org422;
  wire [9:0] _add_all_x_data_out_org423;
  wire [9:0] _add_all_x_data_out_org424;
  wire [9:0] _add_all_x_data_out_org425;
  wire [9:0] _add_all_x_data_out_org426;
  wire [9:0] _add_all_x_data_out_org427;
  wire [9:0] _add_all_x_data_out_org428;
  wire [9:0] _add_all_x_data_out_org429;
  wire [9:0] _add_all_x_data_out_org430;
  wire [9:0] _add_all_x_data_out_org431;
  wire [9:0] _add_all_x_data_out_org432;
  wire [9:0] _add_all_x_data_out_org433;
  wire [9:0] _add_all_x_data_out_org434;
  wire [9:0] _add_all_x_data_out_org435;
  wire [9:0] _add_all_x_data_out_org436;
  wire [9:0] _add_all_x_data_out_org437;
  wire [9:0] _add_all_x_data_out_org438;
  wire [9:0] _add_all_x_data_out_org439;
  wire [9:0] _add_all_x_data_out_org440;
  wire [9:0] _add_all_x_data_out_org441;
  wire [9:0] _add_all_x_data_out_org442;
  wire [9:0] _add_all_x_data_out_org443;
  wire [9:0] _add_all_x_data_out_org444;
  wire [9:0] _add_all_x_data_out_org445;
  wire [9:0] _add_all_x_data_out_org446;
  wire [9:0] _add_all_x_data_out_org449;
  wire [9:0] _add_all_x_data_out_org450;
  wire [9:0] _add_all_x_data_out_org451;
  wire [9:0] _add_all_x_data_out_org452;
  wire [9:0] _add_all_x_data_out_org453;
  wire [9:0] _add_all_x_data_out_org454;
  wire [9:0] _add_all_x_data_out_org455;
  wire [9:0] _add_all_x_data_out_org456;
  wire [9:0] _add_all_x_data_out_org457;
  wire [9:0] _add_all_x_data_out_org458;
  wire [9:0] _add_all_x_data_out_org459;
  wire [9:0] _add_all_x_data_out_org460;
  wire [9:0] _add_all_x_data_out_org461;
  wire [9:0] _add_all_x_data_out_org462;
  wire [9:0] _add_all_x_data_out_org463;
  wire [9:0] _add_all_x_data_out_org464;
  wire [9:0] _add_all_x_data_out_org465;
  wire [9:0] _add_all_x_data_out_org466;
  wire [9:0] _add_all_x_data_out_org467;
  wire [9:0] _add_all_x_data_out_org468;
  wire [9:0] _add_all_x_data_out_org469;
  wire [9:0] _add_all_x_data_out_org470;
  wire [9:0] _add_all_x_data_out_org471;
  wire [9:0] _add_all_x_data_out_org472;
  wire [9:0] _add_all_x_data_out_org473;
  wire [9:0] _add_all_x_data_out_org474;
  wire [9:0] _add_all_x_data_out_org475;
  wire [9:0] _add_all_x_data_out_org476;
  wire [9:0] _add_all_x_data_out_org477;
  wire [9:0] _add_all_x_data_out_org478;
  wire [9:0] _add_all_x_data_in_org33;
  wire [9:0] _add_all_x_data_in_org34;
  wire [9:0] _add_all_x_data_in_org35;
  wire [9:0] _add_all_x_data_in_org36;
  wire [9:0] _add_all_x_data_in_org37;
  wire [9:0] _add_all_x_data_in_org38;
  wire [9:0] _add_all_x_data_in_org39;
  wire [9:0] _add_all_x_data_in_org40;
  wire [9:0] _add_all_x_data_in_org41;
  wire [9:0] _add_all_x_data_in_org42;
  wire [9:0] _add_all_x_data_in_org43;
  wire [9:0] _add_all_x_data_in_org44;
  wire [9:0] _add_all_x_data_in_org45;
  wire [9:0] _add_all_x_data_in_org46;
  wire [9:0] _add_all_x_data_in_org47;
  wire [9:0] _add_all_x_data_in_org48;
  wire [9:0] _add_all_x_data_in_org49;
  wire [9:0] _add_all_x_data_in_org50;
  wire [9:0] _add_all_x_data_in_org51;
  wire [9:0] _add_all_x_data_in_org52;
  wire [9:0] _add_all_x_data_in_org53;
  wire [9:0] _add_all_x_data_in_org54;
  wire [9:0] _add_all_x_data_in_org55;
  wire [9:0] _add_all_x_data_in_org56;
  wire [9:0] _add_all_x_data_in_org57;
  wire [9:0] _add_all_x_data_in_org58;
  wire [9:0] _add_all_x_data_in_org59;
  wire [9:0] _add_all_x_data_in_org60;
  wire [9:0] _add_all_x_data_in_org61;
  wire [9:0] _add_all_x_data_in_org62;
  wire [9:0] _add_all_x_data_in_org65;
  wire [9:0] _add_all_x_data_in_org66;
  wire [9:0] _add_all_x_data_in_org67;
  wire [9:0] _add_all_x_data_in_org68;
  wire [9:0] _add_all_x_data_in_org69;
  wire [9:0] _add_all_x_data_in_org70;
  wire [9:0] _add_all_x_data_in_org71;
  wire [9:0] _add_all_x_data_in_org72;
  wire [9:0] _add_all_x_data_in_org73;
  wire [9:0] _add_all_x_data_in_org74;
  wire [9:0] _add_all_x_data_in_org75;
  wire [9:0] _add_all_x_data_in_org76;
  wire [9:0] _add_all_x_data_in_org77;
  wire [9:0] _add_all_x_data_in_org78;
  wire [9:0] _add_all_x_data_in_org79;
  wire [9:0] _add_all_x_data_in_org80;
  wire [9:0] _add_all_x_data_in_org81;
  wire [9:0] _add_all_x_data_in_org82;
  wire [9:0] _add_all_x_data_in_org83;
  wire [9:0] _add_all_x_data_in_org84;
  wire [9:0] _add_all_x_data_in_org85;
  wire [9:0] _add_all_x_data_in_org86;
  wire [9:0] _add_all_x_data_in_org87;
  wire [9:0] _add_all_x_data_in_org88;
  wire [9:0] _add_all_x_data_in_org89;
  wire [9:0] _add_all_x_data_in_org90;
  wire [9:0] _add_all_x_data_in_org91;
  wire [9:0] _add_all_x_data_in_org92;
  wire [9:0] _add_all_x_data_in_org93;
  wire [9:0] _add_all_x_data_in_org94;
  wire [9:0] _add_all_x_data_in_org97;
  wire [9:0] _add_all_x_data_in_org98;
  wire [9:0] _add_all_x_data_in_org99;
  wire [9:0] _add_all_x_data_in_org100;
  wire [9:0] _add_all_x_data_in_org101;
  wire [9:0] _add_all_x_data_in_org102;
  wire [9:0] _add_all_x_data_in_org103;
  wire [9:0] _add_all_x_data_in_org104;
  wire [9:0] _add_all_x_data_in_org105;
  wire [9:0] _add_all_x_data_in_org106;
  wire [9:0] _add_all_x_data_in_org107;
  wire [9:0] _add_all_x_data_in_org108;
  wire [9:0] _add_all_x_data_in_org109;
  wire [9:0] _add_all_x_data_in_org110;
  wire [9:0] _add_all_x_data_in_org111;
  wire [9:0] _add_all_x_data_in_org112;
  wire [9:0] _add_all_x_data_in_org113;
  wire [9:0] _add_all_x_data_in_org114;
  wire [9:0] _add_all_x_data_in_org115;
  wire [9:0] _add_all_x_data_in_org116;
  wire [9:0] _add_all_x_data_in_org117;
  wire [9:0] _add_all_x_data_in_org118;
  wire [9:0] _add_all_x_data_in_org119;
  wire [9:0] _add_all_x_data_in_org120;
  wire [9:0] _add_all_x_data_in_org121;
  wire [9:0] _add_all_x_data_in_org122;
  wire [9:0] _add_all_x_data_in_org123;
  wire [9:0] _add_all_x_data_in_org124;
  wire [9:0] _add_all_x_data_in_org125;
  wire [9:0] _add_all_x_data_in_org126;
  wire [9:0] _add_all_x_data_in_org129;
  wire [9:0] _add_all_x_data_in_org130;
  wire [9:0] _add_all_x_data_in_org131;
  wire [9:0] _add_all_x_data_in_org132;
  wire [9:0] _add_all_x_data_in_org133;
  wire [9:0] _add_all_x_data_in_org134;
  wire [9:0] _add_all_x_data_in_org135;
  wire [9:0] _add_all_x_data_in_org136;
  wire [9:0] _add_all_x_data_in_org137;
  wire [9:0] _add_all_x_data_in_org138;
  wire [9:0] _add_all_x_data_in_org139;
  wire [9:0] _add_all_x_data_in_org140;
  wire [9:0] _add_all_x_data_in_org141;
  wire [9:0] _add_all_x_data_in_org142;
  wire [9:0] _add_all_x_data_in_org143;
  wire [9:0] _add_all_x_data_in_org144;
  wire [9:0] _add_all_x_data_in_org145;
  wire [9:0] _add_all_x_data_in_org146;
  wire [9:0] _add_all_x_data_in_org147;
  wire [9:0] _add_all_x_data_in_org148;
  wire [9:0] _add_all_x_data_in_org149;
  wire [9:0] _add_all_x_data_in_org150;
  wire [9:0] _add_all_x_data_in_org151;
  wire [9:0] _add_all_x_data_in_org152;
  wire [9:0] _add_all_x_data_in_org153;
  wire [9:0] _add_all_x_data_in_org154;
  wire [9:0] _add_all_x_data_in_org155;
  wire [9:0] _add_all_x_data_in_org156;
  wire [9:0] _add_all_x_data_in_org157;
  wire [9:0] _add_all_x_data_in_org158;
  wire [9:0] _add_all_x_data_in_org161;
  wire [9:0] _add_all_x_data_in_org162;
  wire [9:0] _add_all_x_data_in_org163;
  wire [9:0] _add_all_x_data_in_org164;
  wire [9:0] _add_all_x_data_in_org165;
  wire [9:0] _add_all_x_data_in_org166;
  wire [9:0] _add_all_x_data_in_org167;
  wire [9:0] _add_all_x_data_in_org168;
  wire [9:0] _add_all_x_data_in_org169;
  wire [9:0] _add_all_x_data_in_org170;
  wire [9:0] _add_all_x_data_in_org171;
  wire [9:0] _add_all_x_data_in_org172;
  wire [9:0] _add_all_x_data_in_org173;
  wire [9:0] _add_all_x_data_in_org174;
  wire [9:0] _add_all_x_data_in_org175;
  wire [9:0] _add_all_x_data_in_org176;
  wire [9:0] _add_all_x_data_in_org177;
  wire [9:0] _add_all_x_data_in_org178;
  wire [9:0] _add_all_x_data_in_org179;
  wire [9:0] _add_all_x_data_in_org180;
  wire [9:0] _add_all_x_data_in_org181;
  wire [9:0] _add_all_x_data_in_org182;
  wire [9:0] _add_all_x_data_in_org183;
  wire [9:0] _add_all_x_data_in_org184;
  wire [9:0] _add_all_x_data_in_org185;
  wire [9:0] _add_all_x_data_in_org186;
  wire [9:0] _add_all_x_data_in_org187;
  wire [9:0] _add_all_x_data_in_org188;
  wire [9:0] _add_all_x_data_in_org189;
  wire [9:0] _add_all_x_data_in_org190;
  wire [9:0] _add_all_x_data_in_org193;
  wire [9:0] _add_all_x_data_in_org194;
  wire [9:0] _add_all_x_data_in_org195;
  wire [9:0] _add_all_x_data_in_org196;
  wire [9:0] _add_all_x_data_in_org197;
  wire [9:0] _add_all_x_data_in_org198;
  wire [9:0] _add_all_x_data_in_org199;
  wire [9:0] _add_all_x_data_in_org200;
  wire [9:0] _add_all_x_data_in_org201;
  wire [9:0] _add_all_x_data_in_org202;
  wire [9:0] _add_all_x_data_in_org203;
  wire [9:0] _add_all_x_data_in_org204;
  wire [9:0] _add_all_x_data_in_org205;
  wire [9:0] _add_all_x_data_in_org206;
  wire [9:0] _add_all_x_data_in_org207;
  wire [9:0] _add_all_x_data_in_org208;
  wire [9:0] _add_all_x_data_in_org209;
  wire [9:0] _add_all_x_data_in_org210;
  wire [9:0] _add_all_x_data_in_org211;
  wire [9:0] _add_all_x_data_in_org212;
  wire [9:0] _add_all_x_data_in_org213;
  wire [9:0] _add_all_x_data_in_org214;
  wire [9:0] _add_all_x_data_in_org215;
  wire [9:0] _add_all_x_data_in_org216;
  wire [9:0] _add_all_x_data_in_org217;
  wire [9:0] _add_all_x_data_in_org218;
  wire [9:0] _add_all_x_data_in_org219;
  wire [9:0] _add_all_x_data_in_org220;
  wire [9:0] _add_all_x_data_in_org221;
  wire [9:0] _add_all_x_data_in_org222;
  wire [9:0] _add_all_x_data_in_org225;
  wire [9:0] _add_all_x_data_in_org226;
  wire [9:0] _add_all_x_data_in_org227;
  wire [9:0] _add_all_x_data_in_org228;
  wire [9:0] _add_all_x_data_in_org229;
  wire [9:0] _add_all_x_data_in_org230;
  wire [9:0] _add_all_x_data_in_org231;
  wire [9:0] _add_all_x_data_in_org232;
  wire [9:0] _add_all_x_data_in_org233;
  wire [9:0] _add_all_x_data_in_org234;
  wire [9:0] _add_all_x_data_in_org235;
  wire [9:0] _add_all_x_data_in_org236;
  wire [9:0] _add_all_x_data_in_org237;
  wire [9:0] _add_all_x_data_in_org238;
  wire [9:0] _add_all_x_data_in_org239;
  wire [9:0] _add_all_x_data_in_org240;
  wire [9:0] _add_all_x_data_in_org241;
  wire [9:0] _add_all_x_data_in_org242;
  wire [9:0] _add_all_x_data_in_org243;
  wire [9:0] _add_all_x_data_in_org244;
  wire [9:0] _add_all_x_data_in_org245;
  wire [9:0] _add_all_x_data_in_org246;
  wire [9:0] _add_all_x_data_in_org247;
  wire [9:0] _add_all_x_data_in_org248;
  wire [9:0] _add_all_x_data_in_org249;
  wire [9:0] _add_all_x_data_in_org250;
  wire [9:0] _add_all_x_data_in_org251;
  wire [9:0] _add_all_x_data_in_org252;
  wire [9:0] _add_all_x_data_in_org253;
  wire [9:0] _add_all_x_data_in_org254;
  wire [9:0] _add_all_x_data_in_org257;
  wire [9:0] _add_all_x_data_in_org258;
  wire [9:0] _add_all_x_data_in_org259;
  wire [9:0] _add_all_x_data_in_org260;
  wire [9:0] _add_all_x_data_in_org261;
  wire [9:0] _add_all_x_data_in_org262;
  wire [9:0] _add_all_x_data_in_org263;
  wire [9:0] _add_all_x_data_in_org264;
  wire [9:0] _add_all_x_data_in_org265;
  wire [9:0] _add_all_x_data_in_org266;
  wire [9:0] _add_all_x_data_in_org267;
  wire [9:0] _add_all_x_data_in_org268;
  wire [9:0] _add_all_x_data_in_org269;
  wire [9:0] _add_all_x_data_in_org270;
  wire [9:0] _add_all_x_data_in_org271;
  wire [9:0] _add_all_x_data_in_org272;
  wire [9:0] _add_all_x_data_in_org273;
  wire [9:0] _add_all_x_data_in_org274;
  wire [9:0] _add_all_x_data_in_org275;
  wire [9:0] _add_all_x_data_in_org276;
  wire [9:0] _add_all_x_data_in_org277;
  wire [9:0] _add_all_x_data_in_org278;
  wire [9:0] _add_all_x_data_in_org279;
  wire [9:0] _add_all_x_data_in_org280;
  wire [9:0] _add_all_x_data_in_org281;
  wire [9:0] _add_all_x_data_in_org282;
  wire [9:0] _add_all_x_data_in_org283;
  wire [9:0] _add_all_x_data_in_org284;
  wire [9:0] _add_all_x_data_in_org285;
  wire [9:0] _add_all_x_data_in_org286;
  wire [9:0] _add_all_x_data_in_org289;
  wire [9:0] _add_all_x_data_in_org290;
  wire [9:0] _add_all_x_data_in_org291;
  wire [9:0] _add_all_x_data_in_org292;
  wire [9:0] _add_all_x_data_in_org293;
  wire [9:0] _add_all_x_data_in_org294;
  wire [9:0] _add_all_x_data_in_org295;
  wire [9:0] _add_all_x_data_in_org296;
  wire [9:0] _add_all_x_data_in_org297;
  wire [9:0] _add_all_x_data_in_org298;
  wire [9:0] _add_all_x_data_in_org299;
  wire [9:0] _add_all_x_data_in_org300;
  wire [9:0] _add_all_x_data_in_org301;
  wire [9:0] _add_all_x_data_in_org302;
  wire [9:0] _add_all_x_data_in_org303;
  wire [9:0] _add_all_x_data_in_org304;
  wire [9:0] _add_all_x_data_in_org305;
  wire [9:0] _add_all_x_data_in_org306;
  wire [9:0] _add_all_x_data_in_org307;
  wire [9:0] _add_all_x_data_in_org308;
  wire [9:0] _add_all_x_data_in_org309;
  wire [9:0] _add_all_x_data_in_org310;
  wire [9:0] _add_all_x_data_in_org311;
  wire [9:0] _add_all_x_data_in_org312;
  wire [9:0] _add_all_x_data_in_org313;
  wire [9:0] _add_all_x_data_in_org314;
  wire [9:0] _add_all_x_data_in_org315;
  wire [9:0] _add_all_x_data_in_org316;
  wire [9:0] _add_all_x_data_in_org317;
  wire [9:0] _add_all_x_data_in_org318;
  wire [9:0] _add_all_x_data_in_org321;
  wire [9:0] _add_all_x_data_in_org322;
  wire [9:0] _add_all_x_data_in_org323;
  wire [9:0] _add_all_x_data_in_org324;
  wire [9:0] _add_all_x_data_in_org325;
  wire [9:0] _add_all_x_data_in_org326;
  wire [9:0] _add_all_x_data_in_org327;
  wire [9:0] _add_all_x_data_in_org328;
  wire [9:0] _add_all_x_data_in_org329;
  wire [9:0] _add_all_x_data_in_org330;
  wire [9:0] _add_all_x_data_in_org331;
  wire [9:0] _add_all_x_data_in_org332;
  wire [9:0] _add_all_x_data_in_org333;
  wire [9:0] _add_all_x_data_in_org334;
  wire [9:0] _add_all_x_data_in_org335;
  wire [9:0] _add_all_x_data_in_org336;
  wire [9:0] _add_all_x_data_in_org337;
  wire [9:0] _add_all_x_data_in_org338;
  wire [9:0] _add_all_x_data_in_org339;
  wire [9:0] _add_all_x_data_in_org340;
  wire [9:0] _add_all_x_data_in_org341;
  wire [9:0] _add_all_x_data_in_org342;
  wire [9:0] _add_all_x_data_in_org343;
  wire [9:0] _add_all_x_data_in_org344;
  wire [9:0] _add_all_x_data_in_org345;
  wire [9:0] _add_all_x_data_in_org346;
  wire [9:0] _add_all_x_data_in_org347;
  wire [9:0] _add_all_x_data_in_org348;
  wire [9:0] _add_all_x_data_in_org349;
  wire [9:0] _add_all_x_data_in_org350;
  wire [9:0] _add_all_x_data_in_org353;
  wire [9:0] _add_all_x_data_in_org354;
  wire [9:0] _add_all_x_data_in_org355;
  wire [9:0] _add_all_x_data_in_org356;
  wire [9:0] _add_all_x_data_in_org357;
  wire [9:0] _add_all_x_data_in_org358;
  wire [9:0] _add_all_x_data_in_org359;
  wire [9:0] _add_all_x_data_in_org360;
  wire [9:0] _add_all_x_data_in_org361;
  wire [9:0] _add_all_x_data_in_org362;
  wire [9:0] _add_all_x_data_in_org363;
  wire [9:0] _add_all_x_data_in_org364;
  wire [9:0] _add_all_x_data_in_org365;
  wire [9:0] _add_all_x_data_in_org366;
  wire [9:0] _add_all_x_data_in_org367;
  wire [9:0] _add_all_x_data_in_org368;
  wire [9:0] _add_all_x_data_in_org369;
  wire [9:0] _add_all_x_data_in_org370;
  wire [9:0] _add_all_x_data_in_org371;
  wire [9:0] _add_all_x_data_in_org372;
  wire [9:0] _add_all_x_data_in_org373;
  wire [9:0] _add_all_x_data_in_org374;
  wire [9:0] _add_all_x_data_in_org375;
  wire [9:0] _add_all_x_data_in_org376;
  wire [9:0] _add_all_x_data_in_org377;
  wire [9:0] _add_all_x_data_in_org378;
  wire [9:0] _add_all_x_data_in_org379;
  wire [9:0] _add_all_x_data_in_org380;
  wire [9:0] _add_all_x_data_in_org381;
  wire [9:0] _add_all_x_data_in_org382;
  wire [9:0] _add_all_x_data_in_org385;
  wire [9:0] _add_all_x_data_in_org386;
  wire [9:0] _add_all_x_data_in_org387;
  wire [9:0] _add_all_x_data_in_org388;
  wire [9:0] _add_all_x_data_in_org389;
  wire [9:0] _add_all_x_data_in_org390;
  wire [9:0] _add_all_x_data_in_org391;
  wire [9:0] _add_all_x_data_in_org392;
  wire [9:0] _add_all_x_data_in_org393;
  wire [9:0] _add_all_x_data_in_org394;
  wire [9:0] _add_all_x_data_in_org395;
  wire [9:0] _add_all_x_data_in_org396;
  wire [9:0] _add_all_x_data_in_org397;
  wire [9:0] _add_all_x_data_in_org398;
  wire [9:0] _add_all_x_data_in_org399;
  wire [9:0] _add_all_x_data_in_org400;
  wire [9:0] _add_all_x_data_in_org401;
  wire [9:0] _add_all_x_data_in_org402;
  wire [9:0] _add_all_x_data_in_org403;
  wire [9:0] _add_all_x_data_in_org404;
  wire [9:0] _add_all_x_data_in_org405;
  wire [9:0] _add_all_x_data_in_org406;
  wire [9:0] _add_all_x_data_in_org407;
  wire [9:0] _add_all_x_data_in_org408;
  wire [9:0] _add_all_x_data_in_org409;
  wire [9:0] _add_all_x_data_in_org410;
  wire [9:0] _add_all_x_data_in_org411;
  wire [9:0] _add_all_x_data_in_org412;
  wire [9:0] _add_all_x_data_in_org413;
  wire [9:0] _add_all_x_data_in_org414;
  wire [9:0] _add_all_x_data_in_org417;
  wire [9:0] _add_all_x_data_in_org418;
  wire [9:0] _add_all_x_data_in_org419;
  wire [9:0] _add_all_x_data_in_org420;
  wire [9:0] _add_all_x_data_in_org421;
  wire [9:0] _add_all_x_data_in_org422;
  wire [9:0] _add_all_x_data_in_org423;
  wire [9:0] _add_all_x_data_in_org424;
  wire [9:0] _add_all_x_data_in_org425;
  wire [9:0] _add_all_x_data_in_org426;
  wire [9:0] _add_all_x_data_in_org427;
  wire [9:0] _add_all_x_data_in_org428;
  wire [9:0] _add_all_x_data_in_org429;
  wire [9:0] _add_all_x_data_in_org430;
  wire [9:0] _add_all_x_data_in_org431;
  wire [9:0] _add_all_x_data_in_org432;
  wire [9:0] _add_all_x_data_in_org433;
  wire [9:0] _add_all_x_data_in_org434;
  wire [9:0] _add_all_x_data_in_org435;
  wire [9:0] _add_all_x_data_in_org436;
  wire [9:0] _add_all_x_data_in_org437;
  wire [9:0] _add_all_x_data_in_org438;
  wire [9:0] _add_all_x_data_in_org439;
  wire [9:0] _add_all_x_data_in_org440;
  wire [9:0] _add_all_x_data_in_org441;
  wire [9:0] _add_all_x_data_in_org442;
  wire [9:0] _add_all_x_data_in_org443;
  wire [9:0] _add_all_x_data_in_org444;
  wire [9:0] _add_all_x_data_in_org445;
  wire [9:0] _add_all_x_data_in_org446;
  wire [9:0] _add_all_x_data_in_org449;
  wire [9:0] _add_all_x_data_in_org450;
  wire [9:0] _add_all_x_data_in_org451;
  wire [9:0] _add_all_x_data_in_org452;
  wire [9:0] _add_all_x_data_in_org453;
  wire [9:0] _add_all_x_data_in_org454;
  wire [9:0] _add_all_x_data_in_org455;
  wire [9:0] _add_all_x_data_in_org456;
  wire [9:0] _add_all_x_data_in_org457;
  wire [9:0] _add_all_x_data_in_org458;
  wire [9:0] _add_all_x_data_in_org459;
  wire [9:0] _add_all_x_data_in_org460;
  wire [9:0] _add_all_x_data_in_org461;
  wire [9:0] _add_all_x_data_in_org462;
  wire [9:0] _add_all_x_data_in_org463;
  wire [9:0] _add_all_x_data_in_org464;
  wire [9:0] _add_all_x_data_in_org465;
  wire [9:0] _add_all_x_data_in_org466;
  wire [9:0] _add_all_x_data_in_org467;
  wire [9:0] _add_all_x_data_in_org468;
  wire [9:0] _add_all_x_data_in_org469;
  wire [9:0] _add_all_x_data_in_org470;
  wire [9:0] _add_all_x_data_in_org471;
  wire [9:0] _add_all_x_data_in_org472;
  wire [9:0] _add_all_x_data_in_org473;
  wire [9:0] _add_all_x_data_in_org474;
  wire [9:0] _add_all_x_data_in_org475;
  wire [9:0] _add_all_x_data_in_org476;
  wire [9:0] _add_all_x_data_in_org477;
  wire [9:0] _add_all_x_data_in_org478;
  wire [9:0] _add_all_x_data_out33;
  wire [9:0] _add_all_x_data_out34;
  wire [9:0] _add_all_x_data_out35;
  wire [9:0] _add_all_x_data_out36;
  wire [9:0] _add_all_x_data_out37;
  wire [9:0] _add_all_x_data_out38;
  wire [9:0] _add_all_x_data_out39;
  wire [9:0] _add_all_x_data_out40;
  wire [9:0] _add_all_x_data_out41;
  wire [9:0] _add_all_x_data_out42;
  wire [9:0] _add_all_x_data_out43;
  wire [9:0] _add_all_x_data_out44;
  wire [9:0] _add_all_x_data_out45;
  wire [9:0] _add_all_x_data_out46;
  wire [9:0] _add_all_x_data_out47;
  wire [9:0] _add_all_x_data_out48;
  wire [9:0] _add_all_x_data_out49;
  wire [9:0] _add_all_x_data_out50;
  wire [9:0] _add_all_x_data_out51;
  wire [9:0] _add_all_x_data_out52;
  wire [9:0] _add_all_x_data_out53;
  wire [9:0] _add_all_x_data_out54;
  wire [9:0] _add_all_x_data_out55;
  wire [9:0] _add_all_x_data_out56;
  wire [9:0] _add_all_x_data_out57;
  wire [9:0] _add_all_x_data_out58;
  wire [9:0] _add_all_x_data_out59;
  wire [9:0] _add_all_x_data_out60;
  wire [9:0] _add_all_x_data_out61;
  wire [9:0] _add_all_x_data_out62;
  wire [9:0] _add_all_x_data_out65;
  wire [9:0] _add_all_x_data_out66;
  wire [9:0] _add_all_x_data_out67;
  wire [9:0] _add_all_x_data_out68;
  wire [9:0] _add_all_x_data_out69;
  wire [9:0] _add_all_x_data_out70;
  wire [9:0] _add_all_x_data_out71;
  wire [9:0] _add_all_x_data_out72;
  wire [9:0] _add_all_x_data_out73;
  wire [9:0] _add_all_x_data_out74;
  wire [9:0] _add_all_x_data_out75;
  wire [9:0] _add_all_x_data_out76;
  wire [9:0] _add_all_x_data_out77;
  wire [9:0] _add_all_x_data_out78;
  wire [9:0] _add_all_x_data_out79;
  wire [9:0] _add_all_x_data_out80;
  wire [9:0] _add_all_x_data_out81;
  wire [9:0] _add_all_x_data_out82;
  wire [9:0] _add_all_x_data_out83;
  wire [9:0] _add_all_x_data_out84;
  wire [9:0] _add_all_x_data_out85;
  wire [9:0] _add_all_x_data_out86;
  wire [9:0] _add_all_x_data_out87;
  wire [9:0] _add_all_x_data_out88;
  wire [9:0] _add_all_x_data_out89;
  wire [9:0] _add_all_x_data_out90;
  wire [9:0] _add_all_x_data_out91;
  wire [9:0] _add_all_x_data_out92;
  wire [9:0] _add_all_x_data_out93;
  wire [9:0] _add_all_x_data_out94;
  wire [9:0] _add_all_x_data_out97;
  wire [9:0] _add_all_x_data_out98;
  wire [9:0] _add_all_x_data_out99;
  wire [9:0] _add_all_x_data_out100;
  wire [9:0] _add_all_x_data_out101;
  wire [9:0] _add_all_x_data_out102;
  wire [9:0] _add_all_x_data_out103;
  wire [9:0] _add_all_x_data_out104;
  wire [9:0] _add_all_x_data_out105;
  wire [9:0] _add_all_x_data_out106;
  wire [9:0] _add_all_x_data_out107;
  wire [9:0] _add_all_x_data_out108;
  wire [9:0] _add_all_x_data_out109;
  wire [9:0] _add_all_x_data_out110;
  wire [9:0] _add_all_x_data_out111;
  wire [9:0] _add_all_x_data_out112;
  wire [9:0] _add_all_x_data_out113;
  wire [9:0] _add_all_x_data_out114;
  wire [9:0] _add_all_x_data_out115;
  wire [9:0] _add_all_x_data_out116;
  wire [9:0] _add_all_x_data_out117;
  wire [9:0] _add_all_x_data_out118;
  wire [9:0] _add_all_x_data_out119;
  wire [9:0] _add_all_x_data_out120;
  wire [9:0] _add_all_x_data_out121;
  wire [9:0] _add_all_x_data_out122;
  wire [9:0] _add_all_x_data_out123;
  wire [9:0] _add_all_x_data_out124;
  wire [9:0] _add_all_x_data_out125;
  wire [9:0] _add_all_x_data_out126;
  wire [9:0] _add_all_x_data_out129;
  wire [9:0] _add_all_x_data_out130;
  wire [9:0] _add_all_x_data_out131;
  wire [9:0] _add_all_x_data_out132;
  wire [9:0] _add_all_x_data_out133;
  wire [9:0] _add_all_x_data_out134;
  wire [9:0] _add_all_x_data_out135;
  wire [9:0] _add_all_x_data_out136;
  wire [9:0] _add_all_x_data_out137;
  wire [9:0] _add_all_x_data_out138;
  wire [9:0] _add_all_x_data_out139;
  wire [9:0] _add_all_x_data_out140;
  wire [9:0] _add_all_x_data_out141;
  wire [9:0] _add_all_x_data_out142;
  wire [9:0] _add_all_x_data_out143;
  wire [9:0] _add_all_x_data_out144;
  wire [9:0] _add_all_x_data_out145;
  wire [9:0] _add_all_x_data_out146;
  wire [9:0] _add_all_x_data_out147;
  wire [9:0] _add_all_x_data_out148;
  wire [9:0] _add_all_x_data_out149;
  wire [9:0] _add_all_x_data_out150;
  wire [9:0] _add_all_x_data_out151;
  wire [9:0] _add_all_x_data_out152;
  wire [9:0] _add_all_x_data_out153;
  wire [9:0] _add_all_x_data_out154;
  wire [9:0] _add_all_x_data_out155;
  wire [9:0] _add_all_x_data_out156;
  wire [9:0] _add_all_x_data_out157;
  wire [9:0] _add_all_x_data_out158;
  wire [9:0] _add_all_x_data_out161;
  wire [9:0] _add_all_x_data_out162;
  wire [9:0] _add_all_x_data_out163;
  wire [9:0] _add_all_x_data_out164;
  wire [9:0] _add_all_x_data_out165;
  wire [9:0] _add_all_x_data_out166;
  wire [9:0] _add_all_x_data_out167;
  wire [9:0] _add_all_x_data_out168;
  wire [9:0] _add_all_x_data_out169;
  wire [9:0] _add_all_x_data_out170;
  wire [9:0] _add_all_x_data_out171;
  wire [9:0] _add_all_x_data_out172;
  wire [9:0] _add_all_x_data_out173;
  wire [9:0] _add_all_x_data_out174;
  wire [9:0] _add_all_x_data_out175;
  wire [9:0] _add_all_x_data_out176;
  wire [9:0] _add_all_x_data_out177;
  wire [9:0] _add_all_x_data_out178;
  wire [9:0] _add_all_x_data_out179;
  wire [9:0] _add_all_x_data_out180;
  wire [9:0] _add_all_x_data_out181;
  wire [9:0] _add_all_x_data_out182;
  wire [9:0] _add_all_x_data_out183;
  wire [9:0] _add_all_x_data_out184;
  wire [9:0] _add_all_x_data_out185;
  wire [9:0] _add_all_x_data_out186;
  wire [9:0] _add_all_x_data_out187;
  wire [9:0] _add_all_x_data_out188;
  wire [9:0] _add_all_x_data_out189;
  wire [9:0] _add_all_x_data_out190;
  wire [9:0] _add_all_x_data_out193;
  wire [9:0] _add_all_x_data_out194;
  wire [9:0] _add_all_x_data_out195;
  wire [9:0] _add_all_x_data_out196;
  wire [9:0] _add_all_x_data_out197;
  wire [9:0] _add_all_x_data_out198;
  wire [9:0] _add_all_x_data_out199;
  wire [9:0] _add_all_x_data_out200;
  wire [9:0] _add_all_x_data_out201;
  wire [9:0] _add_all_x_data_out202;
  wire [9:0] _add_all_x_data_out203;
  wire [9:0] _add_all_x_data_out204;
  wire [9:0] _add_all_x_data_out205;
  wire [9:0] _add_all_x_data_out206;
  wire [9:0] _add_all_x_data_out207;
  wire [9:0] _add_all_x_data_out208;
  wire [9:0] _add_all_x_data_out209;
  wire [9:0] _add_all_x_data_out210;
  wire [9:0] _add_all_x_data_out211;
  wire [9:0] _add_all_x_data_out212;
  wire [9:0] _add_all_x_data_out213;
  wire [9:0] _add_all_x_data_out214;
  wire [9:0] _add_all_x_data_out215;
  wire [9:0] _add_all_x_data_out216;
  wire [9:0] _add_all_x_data_out217;
  wire [9:0] _add_all_x_data_out218;
  wire [9:0] _add_all_x_data_out219;
  wire [9:0] _add_all_x_data_out220;
  wire [9:0] _add_all_x_data_out221;
  wire [9:0] _add_all_x_data_out222;
  wire [9:0] _add_all_x_data_out225;
  wire [9:0] _add_all_x_data_out226;
  wire [9:0] _add_all_x_data_out227;
  wire [9:0] _add_all_x_data_out228;
  wire [9:0] _add_all_x_data_out229;
  wire [9:0] _add_all_x_data_out230;
  wire [9:0] _add_all_x_data_out231;
  wire [9:0] _add_all_x_data_out232;
  wire [9:0] _add_all_x_data_out233;
  wire [9:0] _add_all_x_data_out234;
  wire [9:0] _add_all_x_data_out235;
  wire [9:0] _add_all_x_data_out236;
  wire [9:0] _add_all_x_data_out237;
  wire [9:0] _add_all_x_data_out238;
  wire [9:0] _add_all_x_data_out239;
  wire [9:0] _add_all_x_data_out240;
  wire [9:0] _add_all_x_data_out241;
  wire [9:0] _add_all_x_data_out242;
  wire [9:0] _add_all_x_data_out243;
  wire [9:0] _add_all_x_data_out244;
  wire [9:0] _add_all_x_data_out245;
  wire [9:0] _add_all_x_data_out246;
  wire [9:0] _add_all_x_data_out247;
  wire [9:0] _add_all_x_data_out248;
  wire [9:0] _add_all_x_data_out249;
  wire [9:0] _add_all_x_data_out250;
  wire [9:0] _add_all_x_data_out251;
  wire [9:0] _add_all_x_data_out252;
  wire [9:0] _add_all_x_data_out253;
  wire [9:0] _add_all_x_data_out254;
  wire [9:0] _add_all_x_data_out257;
  wire [9:0] _add_all_x_data_out258;
  wire [9:0] _add_all_x_data_out259;
  wire [9:0] _add_all_x_data_out260;
  wire [9:0] _add_all_x_data_out261;
  wire [9:0] _add_all_x_data_out262;
  wire [9:0] _add_all_x_data_out263;
  wire [9:0] _add_all_x_data_out264;
  wire [9:0] _add_all_x_data_out265;
  wire [9:0] _add_all_x_data_out266;
  wire [9:0] _add_all_x_data_out267;
  wire [9:0] _add_all_x_data_out268;
  wire [9:0] _add_all_x_data_out269;
  wire [9:0] _add_all_x_data_out270;
  wire [9:0] _add_all_x_data_out271;
  wire [9:0] _add_all_x_data_out272;
  wire [9:0] _add_all_x_data_out273;
  wire [9:0] _add_all_x_data_out274;
  wire [9:0] _add_all_x_data_out275;
  wire [9:0] _add_all_x_data_out276;
  wire [9:0] _add_all_x_data_out277;
  wire [9:0] _add_all_x_data_out278;
  wire [9:0] _add_all_x_data_out279;
  wire [9:0] _add_all_x_data_out280;
  wire [9:0] _add_all_x_data_out281;
  wire [9:0] _add_all_x_data_out282;
  wire [9:0] _add_all_x_data_out283;
  wire [9:0] _add_all_x_data_out284;
  wire [9:0] _add_all_x_data_out285;
  wire [9:0] _add_all_x_data_out286;
  wire [9:0] _add_all_x_data_out289;
  wire [9:0] _add_all_x_data_out290;
  wire [9:0] _add_all_x_data_out291;
  wire [9:0] _add_all_x_data_out292;
  wire [9:0] _add_all_x_data_out293;
  wire [9:0] _add_all_x_data_out294;
  wire [9:0] _add_all_x_data_out295;
  wire [9:0] _add_all_x_data_out296;
  wire [9:0] _add_all_x_data_out297;
  wire [9:0] _add_all_x_data_out298;
  wire [9:0] _add_all_x_data_out299;
  wire [9:0] _add_all_x_data_out300;
  wire [9:0] _add_all_x_data_out301;
  wire [9:0] _add_all_x_data_out302;
  wire [9:0] _add_all_x_data_out303;
  wire [9:0] _add_all_x_data_out304;
  wire [9:0] _add_all_x_data_out305;
  wire [9:0] _add_all_x_data_out306;
  wire [9:0] _add_all_x_data_out307;
  wire [9:0] _add_all_x_data_out308;
  wire [9:0] _add_all_x_data_out309;
  wire [9:0] _add_all_x_data_out310;
  wire [9:0] _add_all_x_data_out311;
  wire [9:0] _add_all_x_data_out312;
  wire [9:0] _add_all_x_data_out313;
  wire [9:0] _add_all_x_data_out314;
  wire [9:0] _add_all_x_data_out315;
  wire [9:0] _add_all_x_data_out316;
  wire [9:0] _add_all_x_data_out317;
  wire [9:0] _add_all_x_data_out318;
  wire [9:0] _add_all_x_data_out321;
  wire [9:0] _add_all_x_data_out322;
  wire [9:0] _add_all_x_data_out323;
  wire [9:0] _add_all_x_data_out324;
  wire [9:0] _add_all_x_data_out325;
  wire [9:0] _add_all_x_data_out326;
  wire [9:0] _add_all_x_data_out327;
  wire [9:0] _add_all_x_data_out328;
  wire [9:0] _add_all_x_data_out329;
  wire [9:0] _add_all_x_data_out330;
  wire [9:0] _add_all_x_data_out331;
  wire [9:0] _add_all_x_data_out332;
  wire [9:0] _add_all_x_data_out333;
  wire [9:0] _add_all_x_data_out334;
  wire [9:0] _add_all_x_data_out335;
  wire [9:0] _add_all_x_data_out336;
  wire [9:0] _add_all_x_data_out337;
  wire [9:0] _add_all_x_data_out338;
  wire [9:0] _add_all_x_data_out339;
  wire [9:0] _add_all_x_data_out340;
  wire [9:0] _add_all_x_data_out341;
  wire [9:0] _add_all_x_data_out342;
  wire [9:0] _add_all_x_data_out343;
  wire [9:0] _add_all_x_data_out344;
  wire [9:0] _add_all_x_data_out345;
  wire [9:0] _add_all_x_data_out346;
  wire [9:0] _add_all_x_data_out347;
  wire [9:0] _add_all_x_data_out348;
  wire [9:0] _add_all_x_data_out349;
  wire [9:0] _add_all_x_data_out350;
  wire [9:0] _add_all_x_data_out353;
  wire [9:0] _add_all_x_data_out354;
  wire [9:0] _add_all_x_data_out355;
  wire [9:0] _add_all_x_data_out356;
  wire [9:0] _add_all_x_data_out357;
  wire [9:0] _add_all_x_data_out358;
  wire [9:0] _add_all_x_data_out359;
  wire [9:0] _add_all_x_data_out360;
  wire [9:0] _add_all_x_data_out361;
  wire [9:0] _add_all_x_data_out362;
  wire [9:0] _add_all_x_data_out363;
  wire [9:0] _add_all_x_data_out364;
  wire [9:0] _add_all_x_data_out365;
  wire [9:0] _add_all_x_data_out366;
  wire [9:0] _add_all_x_data_out367;
  wire [9:0] _add_all_x_data_out368;
  wire [9:0] _add_all_x_data_out369;
  wire [9:0] _add_all_x_data_out370;
  wire [9:0] _add_all_x_data_out371;
  wire [9:0] _add_all_x_data_out372;
  wire [9:0] _add_all_x_data_out373;
  wire [9:0] _add_all_x_data_out374;
  wire [9:0] _add_all_x_data_out375;
  wire [9:0] _add_all_x_data_out376;
  wire [9:0] _add_all_x_data_out377;
  wire [9:0] _add_all_x_data_out378;
  wire [9:0] _add_all_x_data_out379;
  wire [9:0] _add_all_x_data_out380;
  wire [9:0] _add_all_x_data_out381;
  wire [9:0] _add_all_x_data_out382;
  wire [9:0] _add_all_x_data_out385;
  wire [9:0] _add_all_x_data_out386;
  wire [9:0] _add_all_x_data_out387;
  wire [9:0] _add_all_x_data_out388;
  wire [9:0] _add_all_x_data_out389;
  wire [9:0] _add_all_x_data_out390;
  wire [9:0] _add_all_x_data_out391;
  wire [9:0] _add_all_x_data_out392;
  wire [9:0] _add_all_x_data_out393;
  wire [9:0] _add_all_x_data_out394;
  wire [9:0] _add_all_x_data_out395;
  wire [9:0] _add_all_x_data_out396;
  wire [9:0] _add_all_x_data_out397;
  wire [9:0] _add_all_x_data_out398;
  wire [9:0] _add_all_x_data_out399;
  wire [9:0] _add_all_x_data_out400;
  wire [9:0] _add_all_x_data_out401;
  wire [9:0] _add_all_x_data_out402;
  wire [9:0] _add_all_x_data_out403;
  wire [9:0] _add_all_x_data_out404;
  wire [9:0] _add_all_x_data_out405;
  wire [9:0] _add_all_x_data_out406;
  wire [9:0] _add_all_x_data_out407;
  wire [9:0] _add_all_x_data_out408;
  wire [9:0] _add_all_x_data_out409;
  wire [9:0] _add_all_x_data_out410;
  wire [9:0] _add_all_x_data_out411;
  wire [9:0] _add_all_x_data_out412;
  wire [9:0] _add_all_x_data_out413;
  wire [9:0] _add_all_x_data_out414;
  wire [9:0] _add_all_x_data_out417;
  wire [9:0] _add_all_x_data_out418;
  wire [9:0] _add_all_x_data_out419;
  wire [9:0] _add_all_x_data_out420;
  wire [9:0] _add_all_x_data_out421;
  wire [9:0] _add_all_x_data_out422;
  wire [9:0] _add_all_x_data_out423;
  wire [9:0] _add_all_x_data_out424;
  wire [9:0] _add_all_x_data_out425;
  wire [9:0] _add_all_x_data_out426;
  wire [9:0] _add_all_x_data_out427;
  wire [9:0] _add_all_x_data_out428;
  wire [9:0] _add_all_x_data_out429;
  wire [9:0] _add_all_x_data_out430;
  wire [9:0] _add_all_x_data_out431;
  wire [9:0] _add_all_x_data_out432;
  wire [9:0] _add_all_x_data_out433;
  wire [9:0] _add_all_x_data_out434;
  wire [9:0] _add_all_x_data_out435;
  wire [9:0] _add_all_x_data_out436;
  wire [9:0] _add_all_x_data_out437;
  wire [9:0] _add_all_x_data_out438;
  wire [9:0] _add_all_x_data_out439;
  wire [9:0] _add_all_x_data_out440;
  wire [9:0] _add_all_x_data_out441;
  wire [9:0] _add_all_x_data_out442;
  wire [9:0] _add_all_x_data_out443;
  wire [9:0] _add_all_x_data_out444;
  wire [9:0] _add_all_x_data_out445;
  wire [9:0] _add_all_x_data_out446;
  wire [9:0] _add_all_x_data_out449;
  wire [9:0] _add_all_x_data_out450;
  wire [9:0] _add_all_x_data_out451;
  wire [9:0] _add_all_x_data_out452;
  wire [9:0] _add_all_x_data_out453;
  wire [9:0] _add_all_x_data_out454;
  wire [9:0] _add_all_x_data_out455;
  wire [9:0] _add_all_x_data_out456;
  wire [9:0] _add_all_x_data_out457;
  wire [9:0] _add_all_x_data_out458;
  wire [9:0] _add_all_x_data_out459;
  wire [9:0] _add_all_x_data_out460;
  wire [9:0] _add_all_x_data_out461;
  wire [9:0] _add_all_x_data_out462;
  wire [9:0] _add_all_x_data_out463;
  wire [9:0] _add_all_x_data_out464;
  wire [9:0] _add_all_x_data_out465;
  wire [9:0] _add_all_x_data_out466;
  wire [9:0] _add_all_x_data_out467;
  wire [9:0] _add_all_x_data_out468;
  wire [9:0] _add_all_x_data_out469;
  wire [9:0] _add_all_x_data_out470;
  wire [9:0] _add_all_x_data_out471;
  wire [9:0] _add_all_x_data_out472;
  wire [9:0] _add_all_x_data_out473;
  wire [9:0] _add_all_x_data_out474;
  wire [9:0] _add_all_x_data_out475;
  wire [9:0] _add_all_x_data_out476;
  wire [9:0] _add_all_x_data_out477;
  wire [9:0] _add_all_x_data_out478;
  wire [9:0] _add_all_x_data_out_index33;
  wire [9:0] _add_all_x_data_out_index34;
  wire [9:0] _add_all_x_data_out_index35;
  wire [9:0] _add_all_x_data_out_index36;
  wire [9:0] _add_all_x_data_out_index37;
  wire [9:0] _add_all_x_data_out_index38;
  wire [9:0] _add_all_x_data_out_index39;
  wire [9:0] _add_all_x_data_out_index40;
  wire [9:0] _add_all_x_data_out_index41;
  wire [9:0] _add_all_x_data_out_index42;
  wire [9:0] _add_all_x_data_out_index43;
  wire [9:0] _add_all_x_data_out_index44;
  wire [9:0] _add_all_x_data_out_index45;
  wire [9:0] _add_all_x_data_out_index46;
  wire [9:0] _add_all_x_data_out_index47;
  wire [9:0] _add_all_x_data_out_index48;
  wire [9:0] _add_all_x_data_out_index49;
  wire [9:0] _add_all_x_data_out_index50;
  wire [9:0] _add_all_x_data_out_index51;
  wire [9:0] _add_all_x_data_out_index52;
  wire [9:0] _add_all_x_data_out_index53;
  wire [9:0] _add_all_x_data_out_index54;
  wire [9:0] _add_all_x_data_out_index55;
  wire [9:0] _add_all_x_data_out_index56;
  wire [9:0] _add_all_x_data_out_index57;
  wire [9:0] _add_all_x_data_out_index58;
  wire [9:0] _add_all_x_data_out_index59;
  wire [9:0] _add_all_x_data_out_index60;
  wire [9:0] _add_all_x_data_out_index61;
  wire [9:0] _add_all_x_data_out_index62;
  wire [9:0] _add_all_x_data_out_index65;
  wire [9:0] _add_all_x_data_out_index66;
  wire [9:0] _add_all_x_data_out_index67;
  wire [9:0] _add_all_x_data_out_index68;
  wire [9:0] _add_all_x_data_out_index69;
  wire [9:0] _add_all_x_data_out_index70;
  wire [9:0] _add_all_x_data_out_index71;
  wire [9:0] _add_all_x_data_out_index72;
  wire [9:0] _add_all_x_data_out_index73;
  wire [9:0] _add_all_x_data_out_index74;
  wire [9:0] _add_all_x_data_out_index75;
  wire [9:0] _add_all_x_data_out_index76;
  wire [9:0] _add_all_x_data_out_index77;
  wire [9:0] _add_all_x_data_out_index78;
  wire [9:0] _add_all_x_data_out_index79;
  wire [9:0] _add_all_x_data_out_index80;
  wire [9:0] _add_all_x_data_out_index81;
  wire [9:0] _add_all_x_data_out_index82;
  wire [9:0] _add_all_x_data_out_index83;
  wire [9:0] _add_all_x_data_out_index84;
  wire [9:0] _add_all_x_data_out_index85;
  wire [9:0] _add_all_x_data_out_index86;
  wire [9:0] _add_all_x_data_out_index87;
  wire [9:0] _add_all_x_data_out_index88;
  wire [9:0] _add_all_x_data_out_index89;
  wire [9:0] _add_all_x_data_out_index90;
  wire [9:0] _add_all_x_data_out_index91;
  wire [9:0] _add_all_x_data_out_index92;
  wire [9:0] _add_all_x_data_out_index93;
  wire [9:0] _add_all_x_data_out_index94;
  wire [9:0] _add_all_x_data_out_index97;
  wire [9:0] _add_all_x_data_out_index98;
  wire [9:0] _add_all_x_data_out_index99;
  wire [9:0] _add_all_x_data_out_index100;
  wire [9:0] _add_all_x_data_out_index101;
  wire [9:0] _add_all_x_data_out_index102;
  wire [9:0] _add_all_x_data_out_index103;
  wire [9:0] _add_all_x_data_out_index104;
  wire [9:0] _add_all_x_data_out_index105;
  wire [9:0] _add_all_x_data_out_index106;
  wire [9:0] _add_all_x_data_out_index107;
  wire [9:0] _add_all_x_data_out_index108;
  wire [9:0] _add_all_x_data_out_index109;
  wire [9:0] _add_all_x_data_out_index110;
  wire [9:0] _add_all_x_data_out_index111;
  wire [9:0] _add_all_x_data_out_index112;
  wire [9:0] _add_all_x_data_out_index113;
  wire [9:0] _add_all_x_data_out_index114;
  wire [9:0] _add_all_x_data_out_index115;
  wire [9:0] _add_all_x_data_out_index116;
  wire [9:0] _add_all_x_data_out_index117;
  wire [9:0] _add_all_x_data_out_index118;
  wire [9:0] _add_all_x_data_out_index119;
  wire [9:0] _add_all_x_data_out_index120;
  wire [9:0] _add_all_x_data_out_index121;
  wire [9:0] _add_all_x_data_out_index122;
  wire [9:0] _add_all_x_data_out_index123;
  wire [9:0] _add_all_x_data_out_index124;
  wire [9:0] _add_all_x_data_out_index125;
  wire [9:0] _add_all_x_data_out_index126;
  wire [9:0] _add_all_x_data_out_index129;
  wire [9:0] _add_all_x_data_out_index130;
  wire [9:0] _add_all_x_data_out_index131;
  wire [9:0] _add_all_x_data_out_index132;
  wire [9:0] _add_all_x_data_out_index133;
  wire [9:0] _add_all_x_data_out_index134;
  wire [9:0] _add_all_x_data_out_index135;
  wire [9:0] _add_all_x_data_out_index136;
  wire [9:0] _add_all_x_data_out_index137;
  wire [9:0] _add_all_x_data_out_index138;
  wire [9:0] _add_all_x_data_out_index139;
  wire [9:0] _add_all_x_data_out_index140;
  wire [9:0] _add_all_x_data_out_index141;
  wire [9:0] _add_all_x_data_out_index142;
  wire [9:0] _add_all_x_data_out_index143;
  wire [9:0] _add_all_x_data_out_index144;
  wire [9:0] _add_all_x_data_out_index145;
  wire [9:0] _add_all_x_data_out_index146;
  wire [9:0] _add_all_x_data_out_index147;
  wire [9:0] _add_all_x_data_out_index148;
  wire [9:0] _add_all_x_data_out_index149;
  wire [9:0] _add_all_x_data_out_index150;
  wire [9:0] _add_all_x_data_out_index151;
  wire [9:0] _add_all_x_data_out_index152;
  wire [9:0] _add_all_x_data_out_index153;
  wire [9:0] _add_all_x_data_out_index154;
  wire [9:0] _add_all_x_data_out_index155;
  wire [9:0] _add_all_x_data_out_index156;
  wire [9:0] _add_all_x_data_out_index157;
  wire [9:0] _add_all_x_data_out_index158;
  wire [9:0] _add_all_x_data_out_index161;
  wire [9:0] _add_all_x_data_out_index162;
  wire [9:0] _add_all_x_data_out_index163;
  wire [9:0] _add_all_x_data_out_index164;
  wire [9:0] _add_all_x_data_out_index165;
  wire [9:0] _add_all_x_data_out_index166;
  wire [9:0] _add_all_x_data_out_index167;
  wire [9:0] _add_all_x_data_out_index168;
  wire [9:0] _add_all_x_data_out_index169;
  wire [9:0] _add_all_x_data_out_index170;
  wire [9:0] _add_all_x_data_out_index171;
  wire [9:0] _add_all_x_data_out_index172;
  wire [9:0] _add_all_x_data_out_index173;
  wire [9:0] _add_all_x_data_out_index174;
  wire [9:0] _add_all_x_data_out_index175;
  wire [9:0] _add_all_x_data_out_index176;
  wire [9:0] _add_all_x_data_out_index177;
  wire [9:0] _add_all_x_data_out_index178;
  wire [9:0] _add_all_x_data_out_index179;
  wire [9:0] _add_all_x_data_out_index180;
  wire [9:0] _add_all_x_data_out_index181;
  wire [9:0] _add_all_x_data_out_index182;
  wire [9:0] _add_all_x_data_out_index183;
  wire [9:0] _add_all_x_data_out_index184;
  wire [9:0] _add_all_x_data_out_index185;
  wire [9:0] _add_all_x_data_out_index186;
  wire [9:0] _add_all_x_data_out_index187;
  wire [9:0] _add_all_x_data_out_index188;
  wire [9:0] _add_all_x_data_out_index189;
  wire [9:0] _add_all_x_data_out_index190;
  wire [9:0] _add_all_x_data_out_index193;
  wire [9:0] _add_all_x_data_out_index194;
  wire [9:0] _add_all_x_data_out_index195;
  wire [9:0] _add_all_x_data_out_index196;
  wire [9:0] _add_all_x_data_out_index197;
  wire [9:0] _add_all_x_data_out_index198;
  wire [9:0] _add_all_x_data_out_index199;
  wire [9:0] _add_all_x_data_out_index200;
  wire [9:0] _add_all_x_data_out_index201;
  wire [9:0] _add_all_x_data_out_index202;
  wire [9:0] _add_all_x_data_out_index203;
  wire [9:0] _add_all_x_data_out_index204;
  wire [9:0] _add_all_x_data_out_index205;
  wire [9:0] _add_all_x_data_out_index206;
  wire [9:0] _add_all_x_data_out_index207;
  wire [9:0] _add_all_x_data_out_index208;
  wire [9:0] _add_all_x_data_out_index209;
  wire [9:0] _add_all_x_data_out_index210;
  wire [9:0] _add_all_x_data_out_index211;
  wire [9:0] _add_all_x_data_out_index212;
  wire [9:0] _add_all_x_data_out_index213;
  wire [9:0] _add_all_x_data_out_index214;
  wire [9:0] _add_all_x_data_out_index215;
  wire [9:0] _add_all_x_data_out_index216;
  wire [9:0] _add_all_x_data_out_index217;
  wire [9:0] _add_all_x_data_out_index218;
  wire [9:0] _add_all_x_data_out_index219;
  wire [9:0] _add_all_x_data_out_index220;
  wire [9:0] _add_all_x_data_out_index221;
  wire [9:0] _add_all_x_data_out_index222;
  wire [9:0] _add_all_x_data_out_index225;
  wire [9:0] _add_all_x_data_out_index226;
  wire [9:0] _add_all_x_data_out_index227;
  wire [9:0] _add_all_x_data_out_index228;
  wire [9:0] _add_all_x_data_out_index229;
  wire [9:0] _add_all_x_data_out_index230;
  wire [9:0] _add_all_x_data_out_index231;
  wire [9:0] _add_all_x_data_out_index232;
  wire [9:0] _add_all_x_data_out_index233;
  wire [9:0] _add_all_x_data_out_index234;
  wire [9:0] _add_all_x_data_out_index235;
  wire [9:0] _add_all_x_data_out_index236;
  wire [9:0] _add_all_x_data_out_index237;
  wire [9:0] _add_all_x_data_out_index238;
  wire [9:0] _add_all_x_data_out_index239;
  wire [9:0] _add_all_x_data_out_index240;
  wire [9:0] _add_all_x_data_out_index241;
  wire [9:0] _add_all_x_data_out_index242;
  wire [9:0] _add_all_x_data_out_index243;
  wire [9:0] _add_all_x_data_out_index244;
  wire [9:0] _add_all_x_data_out_index245;
  wire [9:0] _add_all_x_data_out_index246;
  wire [9:0] _add_all_x_data_out_index247;
  wire [9:0] _add_all_x_data_out_index248;
  wire [9:0] _add_all_x_data_out_index249;
  wire [9:0] _add_all_x_data_out_index250;
  wire [9:0] _add_all_x_data_out_index251;
  wire [9:0] _add_all_x_data_out_index252;
  wire [9:0] _add_all_x_data_out_index253;
  wire [9:0] _add_all_x_data_out_index254;
  wire [9:0] _add_all_x_data_out_index257;
  wire [9:0] _add_all_x_data_out_index258;
  wire [9:0] _add_all_x_data_out_index259;
  wire [9:0] _add_all_x_data_out_index260;
  wire [9:0] _add_all_x_data_out_index261;
  wire [9:0] _add_all_x_data_out_index262;
  wire [9:0] _add_all_x_data_out_index263;
  wire [9:0] _add_all_x_data_out_index264;
  wire [9:0] _add_all_x_data_out_index265;
  wire [9:0] _add_all_x_data_out_index266;
  wire [9:0] _add_all_x_data_out_index267;
  wire [9:0] _add_all_x_data_out_index268;
  wire [9:0] _add_all_x_data_out_index269;
  wire [9:0] _add_all_x_data_out_index270;
  wire [9:0] _add_all_x_data_out_index271;
  wire [9:0] _add_all_x_data_out_index272;
  wire [9:0] _add_all_x_data_out_index273;
  wire [9:0] _add_all_x_data_out_index274;
  wire [9:0] _add_all_x_data_out_index275;
  wire [9:0] _add_all_x_data_out_index276;
  wire [9:0] _add_all_x_data_out_index277;
  wire [9:0] _add_all_x_data_out_index278;
  wire [9:0] _add_all_x_data_out_index279;
  wire [9:0] _add_all_x_data_out_index280;
  wire [9:0] _add_all_x_data_out_index281;
  wire [9:0] _add_all_x_data_out_index282;
  wire [9:0] _add_all_x_data_out_index283;
  wire [9:0] _add_all_x_data_out_index284;
  wire [9:0] _add_all_x_data_out_index285;
  wire [9:0] _add_all_x_data_out_index286;
  wire [9:0] _add_all_x_data_out_index289;
  wire [9:0] _add_all_x_data_out_index290;
  wire [9:0] _add_all_x_data_out_index291;
  wire [9:0] _add_all_x_data_out_index292;
  wire [9:0] _add_all_x_data_out_index293;
  wire [9:0] _add_all_x_data_out_index294;
  wire [9:0] _add_all_x_data_out_index295;
  wire [9:0] _add_all_x_data_out_index296;
  wire [9:0] _add_all_x_data_out_index297;
  wire [9:0] _add_all_x_data_out_index298;
  wire [9:0] _add_all_x_data_out_index299;
  wire [9:0] _add_all_x_data_out_index300;
  wire [9:0] _add_all_x_data_out_index301;
  wire [9:0] _add_all_x_data_out_index302;
  wire [9:0] _add_all_x_data_out_index303;
  wire [9:0] _add_all_x_data_out_index304;
  wire [9:0] _add_all_x_data_out_index305;
  wire [9:0] _add_all_x_data_out_index306;
  wire [9:0] _add_all_x_data_out_index307;
  wire [9:0] _add_all_x_data_out_index308;
  wire [9:0] _add_all_x_data_out_index309;
  wire [9:0] _add_all_x_data_out_index310;
  wire [9:0] _add_all_x_data_out_index311;
  wire [9:0] _add_all_x_data_out_index312;
  wire [9:0] _add_all_x_data_out_index313;
  wire [9:0] _add_all_x_data_out_index314;
  wire [9:0] _add_all_x_data_out_index315;
  wire [9:0] _add_all_x_data_out_index316;
  wire [9:0] _add_all_x_data_out_index317;
  wire [9:0] _add_all_x_data_out_index318;
  wire [9:0] _add_all_x_data_out_index321;
  wire [9:0] _add_all_x_data_out_index322;
  wire [9:0] _add_all_x_data_out_index323;
  wire [9:0] _add_all_x_data_out_index324;
  wire [9:0] _add_all_x_data_out_index325;
  wire [9:0] _add_all_x_data_out_index326;
  wire [9:0] _add_all_x_data_out_index327;
  wire [9:0] _add_all_x_data_out_index328;
  wire [9:0] _add_all_x_data_out_index329;
  wire [9:0] _add_all_x_data_out_index330;
  wire [9:0] _add_all_x_data_out_index331;
  wire [9:0] _add_all_x_data_out_index332;
  wire [9:0] _add_all_x_data_out_index333;
  wire [9:0] _add_all_x_data_out_index334;
  wire [9:0] _add_all_x_data_out_index335;
  wire [9:0] _add_all_x_data_out_index336;
  wire [9:0] _add_all_x_data_out_index337;
  wire [9:0] _add_all_x_data_out_index338;
  wire [9:0] _add_all_x_data_out_index339;
  wire [9:0] _add_all_x_data_out_index340;
  wire [9:0] _add_all_x_data_out_index341;
  wire [9:0] _add_all_x_data_out_index342;
  wire [9:0] _add_all_x_data_out_index343;
  wire [9:0] _add_all_x_data_out_index344;
  wire [9:0] _add_all_x_data_out_index345;
  wire [9:0] _add_all_x_data_out_index346;
  wire [9:0] _add_all_x_data_out_index347;
  wire [9:0] _add_all_x_data_out_index348;
  wire [9:0] _add_all_x_data_out_index349;
  wire [9:0] _add_all_x_data_out_index350;
  wire [9:0] _add_all_x_data_out_index353;
  wire [9:0] _add_all_x_data_out_index354;
  wire [9:0] _add_all_x_data_out_index355;
  wire [9:0] _add_all_x_data_out_index356;
  wire [9:0] _add_all_x_data_out_index357;
  wire [9:0] _add_all_x_data_out_index358;
  wire [9:0] _add_all_x_data_out_index359;
  wire [9:0] _add_all_x_data_out_index360;
  wire [9:0] _add_all_x_data_out_index361;
  wire [9:0] _add_all_x_data_out_index362;
  wire [9:0] _add_all_x_data_out_index363;
  wire [9:0] _add_all_x_data_out_index364;
  wire [9:0] _add_all_x_data_out_index365;
  wire [9:0] _add_all_x_data_out_index366;
  wire [9:0] _add_all_x_data_out_index367;
  wire [9:0] _add_all_x_data_out_index368;
  wire [9:0] _add_all_x_data_out_index369;
  wire [9:0] _add_all_x_data_out_index370;
  wire [9:0] _add_all_x_data_out_index371;
  wire [9:0] _add_all_x_data_out_index372;
  wire [9:0] _add_all_x_data_out_index373;
  wire [9:0] _add_all_x_data_out_index374;
  wire [9:0] _add_all_x_data_out_index375;
  wire [9:0] _add_all_x_data_out_index376;
  wire [9:0] _add_all_x_data_out_index377;
  wire [9:0] _add_all_x_data_out_index378;
  wire [9:0] _add_all_x_data_out_index379;
  wire [9:0] _add_all_x_data_out_index380;
  wire [9:0] _add_all_x_data_out_index381;
  wire [9:0] _add_all_x_data_out_index382;
  wire [9:0] _add_all_x_data_out_index385;
  wire [9:0] _add_all_x_data_out_index386;
  wire [9:0] _add_all_x_data_out_index387;
  wire [9:0] _add_all_x_data_out_index388;
  wire [9:0] _add_all_x_data_out_index389;
  wire [9:0] _add_all_x_data_out_index390;
  wire [9:0] _add_all_x_data_out_index391;
  wire [9:0] _add_all_x_data_out_index392;
  wire [9:0] _add_all_x_data_out_index393;
  wire [9:0] _add_all_x_data_out_index394;
  wire [9:0] _add_all_x_data_out_index395;
  wire [9:0] _add_all_x_data_out_index396;
  wire [9:0] _add_all_x_data_out_index397;
  wire [9:0] _add_all_x_data_out_index398;
  wire [9:0] _add_all_x_data_out_index399;
  wire [9:0] _add_all_x_data_out_index400;
  wire [9:0] _add_all_x_data_out_index401;
  wire [9:0] _add_all_x_data_out_index402;
  wire [9:0] _add_all_x_data_out_index403;
  wire [9:0] _add_all_x_data_out_index404;
  wire [9:0] _add_all_x_data_out_index405;
  wire [9:0] _add_all_x_data_out_index406;
  wire [9:0] _add_all_x_data_out_index407;
  wire [9:0] _add_all_x_data_out_index408;
  wire [9:0] _add_all_x_data_out_index409;
  wire [9:0] _add_all_x_data_out_index410;
  wire [9:0] _add_all_x_data_out_index411;
  wire [9:0] _add_all_x_data_out_index412;
  wire [9:0] _add_all_x_data_out_index413;
  wire [9:0] _add_all_x_data_out_index414;
  wire [9:0] _add_all_x_data_out_index417;
  wire [9:0] _add_all_x_data_out_index418;
  wire [9:0] _add_all_x_data_out_index419;
  wire [9:0] _add_all_x_data_out_index420;
  wire [9:0] _add_all_x_data_out_index421;
  wire [9:0] _add_all_x_data_out_index422;
  wire [9:0] _add_all_x_data_out_index423;
  wire [9:0] _add_all_x_data_out_index424;
  wire [9:0] _add_all_x_data_out_index425;
  wire [9:0] _add_all_x_data_out_index426;
  wire [9:0] _add_all_x_data_out_index427;
  wire [9:0] _add_all_x_data_out_index428;
  wire [9:0] _add_all_x_data_out_index429;
  wire [9:0] _add_all_x_data_out_index430;
  wire [9:0] _add_all_x_data_out_index431;
  wire [9:0] _add_all_x_data_out_index432;
  wire [9:0] _add_all_x_data_out_index433;
  wire [9:0] _add_all_x_data_out_index434;
  wire [9:0] _add_all_x_data_out_index435;
  wire [9:0] _add_all_x_data_out_index436;
  wire [9:0] _add_all_x_data_out_index437;
  wire [9:0] _add_all_x_data_out_index438;
  wire [9:0] _add_all_x_data_out_index439;
  wire [9:0] _add_all_x_data_out_index440;
  wire [9:0] _add_all_x_data_out_index441;
  wire [9:0] _add_all_x_data_out_index442;
  wire [9:0] _add_all_x_data_out_index443;
  wire [9:0] _add_all_x_data_out_index444;
  wire [9:0] _add_all_x_data_out_index445;
  wire [9:0] _add_all_x_data_out_index446;
  wire [9:0] _add_all_x_data_out_index449;
  wire [9:0] _add_all_x_data_out_index450;
  wire [9:0] _add_all_x_data_out_index451;
  wire [9:0] _add_all_x_data_out_index452;
  wire [9:0] _add_all_x_data_out_index453;
  wire [9:0] _add_all_x_data_out_index454;
  wire [9:0] _add_all_x_data_out_index455;
  wire [9:0] _add_all_x_data_out_index456;
  wire [9:0] _add_all_x_data_out_index457;
  wire [9:0] _add_all_x_data_out_index458;
  wire [9:0] _add_all_x_data_out_index459;
  wire [9:0] _add_all_x_data_out_index460;
  wire [9:0] _add_all_x_data_out_index461;
  wire [9:0] _add_all_x_data_out_index462;
  wire [9:0] _add_all_x_data_out_index463;
  wire [9:0] _add_all_x_data_out_index464;
  wire [9:0] _add_all_x_data_out_index465;
  wire [9:0] _add_all_x_data_out_index466;
  wire [9:0] _add_all_x_data_out_index467;
  wire [9:0] _add_all_x_data_out_index468;
  wire [9:0] _add_all_x_data_out_index469;
  wire [9:0] _add_all_x_data_out_index470;
  wire [9:0] _add_all_x_data_out_index471;
  wire [9:0] _add_all_x_data_out_index472;
  wire [9:0] _add_all_x_data_out_index473;
  wire [9:0] _add_all_x_data_out_index474;
  wire [9:0] _add_all_x_data_out_index475;
  wire [9:0] _add_all_x_data_out_index476;
  wire [9:0] _add_all_x_data_out_index477;
  wire [9:0] _add_all_x_data_out_index478;
  wire [1:0] _add_all_x_sg_in33;
  wire [1:0] _add_all_x_sg_in34;
  wire [1:0] _add_all_x_sg_in35;
  wire [1:0] _add_all_x_sg_in36;
  wire [1:0] _add_all_x_sg_in37;
  wire [1:0] _add_all_x_sg_in38;
  wire [1:0] _add_all_x_sg_in39;
  wire [1:0] _add_all_x_sg_in40;
  wire [1:0] _add_all_x_sg_in41;
  wire [1:0] _add_all_x_sg_in42;
  wire [1:0] _add_all_x_sg_in43;
  wire [1:0] _add_all_x_sg_in44;
  wire [1:0] _add_all_x_sg_in45;
  wire [1:0] _add_all_x_sg_in46;
  wire [1:0] _add_all_x_sg_in47;
  wire [1:0] _add_all_x_sg_in48;
  wire [1:0] _add_all_x_sg_in49;
  wire [1:0] _add_all_x_sg_in50;
  wire [1:0] _add_all_x_sg_in51;
  wire [1:0] _add_all_x_sg_in52;
  wire [1:0] _add_all_x_sg_in53;
  wire [1:0] _add_all_x_sg_in54;
  wire [1:0] _add_all_x_sg_in55;
  wire [1:0] _add_all_x_sg_in56;
  wire [1:0] _add_all_x_sg_in57;
  wire [1:0] _add_all_x_sg_in58;
  wire [1:0] _add_all_x_sg_in59;
  wire [1:0] _add_all_x_sg_in60;
  wire [1:0] _add_all_x_sg_in61;
  wire [1:0] _add_all_x_sg_in62;
  wire [1:0] _add_all_x_sg_in65;
  wire [1:0] _add_all_x_sg_in66;
  wire [1:0] _add_all_x_sg_in67;
  wire [1:0] _add_all_x_sg_in68;
  wire [1:0] _add_all_x_sg_in69;
  wire [1:0] _add_all_x_sg_in70;
  wire [1:0] _add_all_x_sg_in71;
  wire [1:0] _add_all_x_sg_in72;
  wire [1:0] _add_all_x_sg_in73;
  wire [1:0] _add_all_x_sg_in74;
  wire [1:0] _add_all_x_sg_in75;
  wire [1:0] _add_all_x_sg_in76;
  wire [1:0] _add_all_x_sg_in77;
  wire [1:0] _add_all_x_sg_in78;
  wire [1:0] _add_all_x_sg_in79;
  wire [1:0] _add_all_x_sg_in80;
  wire [1:0] _add_all_x_sg_in81;
  wire [1:0] _add_all_x_sg_in82;
  wire [1:0] _add_all_x_sg_in83;
  wire [1:0] _add_all_x_sg_in84;
  wire [1:0] _add_all_x_sg_in85;
  wire [1:0] _add_all_x_sg_in86;
  wire [1:0] _add_all_x_sg_in87;
  wire [1:0] _add_all_x_sg_in88;
  wire [1:0] _add_all_x_sg_in89;
  wire [1:0] _add_all_x_sg_in90;
  wire [1:0] _add_all_x_sg_in91;
  wire [1:0] _add_all_x_sg_in92;
  wire [1:0] _add_all_x_sg_in93;
  wire [1:0] _add_all_x_sg_in94;
  wire [1:0] _add_all_x_sg_in97;
  wire [1:0] _add_all_x_sg_in98;
  wire [1:0] _add_all_x_sg_in99;
  wire [1:0] _add_all_x_sg_in100;
  wire [1:0] _add_all_x_sg_in101;
  wire [1:0] _add_all_x_sg_in102;
  wire [1:0] _add_all_x_sg_in103;
  wire [1:0] _add_all_x_sg_in104;
  wire [1:0] _add_all_x_sg_in105;
  wire [1:0] _add_all_x_sg_in106;
  wire [1:0] _add_all_x_sg_in107;
  wire [1:0] _add_all_x_sg_in108;
  wire [1:0] _add_all_x_sg_in109;
  wire [1:0] _add_all_x_sg_in110;
  wire [1:0] _add_all_x_sg_in111;
  wire [1:0] _add_all_x_sg_in112;
  wire [1:0] _add_all_x_sg_in113;
  wire [1:0] _add_all_x_sg_in114;
  wire [1:0] _add_all_x_sg_in115;
  wire [1:0] _add_all_x_sg_in116;
  wire [1:0] _add_all_x_sg_in117;
  wire [1:0] _add_all_x_sg_in118;
  wire [1:0] _add_all_x_sg_in119;
  wire [1:0] _add_all_x_sg_in120;
  wire [1:0] _add_all_x_sg_in121;
  wire [1:0] _add_all_x_sg_in122;
  wire [1:0] _add_all_x_sg_in123;
  wire [1:0] _add_all_x_sg_in124;
  wire [1:0] _add_all_x_sg_in125;
  wire [1:0] _add_all_x_sg_in126;
  wire [1:0] _add_all_x_sg_in129;
  wire [1:0] _add_all_x_sg_in130;
  wire [1:0] _add_all_x_sg_in131;
  wire [1:0] _add_all_x_sg_in132;
  wire [1:0] _add_all_x_sg_in133;
  wire [1:0] _add_all_x_sg_in134;
  wire [1:0] _add_all_x_sg_in135;
  wire [1:0] _add_all_x_sg_in136;
  wire [1:0] _add_all_x_sg_in137;
  wire [1:0] _add_all_x_sg_in138;
  wire [1:0] _add_all_x_sg_in139;
  wire [1:0] _add_all_x_sg_in140;
  wire [1:0] _add_all_x_sg_in141;
  wire [1:0] _add_all_x_sg_in142;
  wire [1:0] _add_all_x_sg_in143;
  wire [1:0] _add_all_x_sg_in144;
  wire [1:0] _add_all_x_sg_in145;
  wire [1:0] _add_all_x_sg_in146;
  wire [1:0] _add_all_x_sg_in147;
  wire [1:0] _add_all_x_sg_in148;
  wire [1:0] _add_all_x_sg_in149;
  wire [1:0] _add_all_x_sg_in150;
  wire [1:0] _add_all_x_sg_in151;
  wire [1:0] _add_all_x_sg_in152;
  wire [1:0] _add_all_x_sg_in153;
  wire [1:0] _add_all_x_sg_in154;
  wire [1:0] _add_all_x_sg_in155;
  wire [1:0] _add_all_x_sg_in156;
  wire [1:0] _add_all_x_sg_in157;
  wire [1:0] _add_all_x_sg_in158;
  wire [1:0] _add_all_x_sg_in161;
  wire [1:0] _add_all_x_sg_in162;
  wire [1:0] _add_all_x_sg_in163;
  wire [1:0] _add_all_x_sg_in164;
  wire [1:0] _add_all_x_sg_in165;
  wire [1:0] _add_all_x_sg_in166;
  wire [1:0] _add_all_x_sg_in167;
  wire [1:0] _add_all_x_sg_in168;
  wire [1:0] _add_all_x_sg_in169;
  wire [1:0] _add_all_x_sg_in170;
  wire [1:0] _add_all_x_sg_in171;
  wire [1:0] _add_all_x_sg_in172;
  wire [1:0] _add_all_x_sg_in173;
  wire [1:0] _add_all_x_sg_in174;
  wire [1:0] _add_all_x_sg_in175;
  wire [1:0] _add_all_x_sg_in176;
  wire [1:0] _add_all_x_sg_in177;
  wire [1:0] _add_all_x_sg_in178;
  wire [1:0] _add_all_x_sg_in179;
  wire [1:0] _add_all_x_sg_in180;
  wire [1:0] _add_all_x_sg_in181;
  wire [1:0] _add_all_x_sg_in182;
  wire [1:0] _add_all_x_sg_in183;
  wire [1:0] _add_all_x_sg_in184;
  wire [1:0] _add_all_x_sg_in185;
  wire [1:0] _add_all_x_sg_in186;
  wire [1:0] _add_all_x_sg_in187;
  wire [1:0] _add_all_x_sg_in188;
  wire [1:0] _add_all_x_sg_in189;
  wire [1:0] _add_all_x_sg_in190;
  wire [1:0] _add_all_x_sg_in193;
  wire [1:0] _add_all_x_sg_in194;
  wire [1:0] _add_all_x_sg_in195;
  wire [1:0] _add_all_x_sg_in196;
  wire [1:0] _add_all_x_sg_in197;
  wire [1:0] _add_all_x_sg_in198;
  wire [1:0] _add_all_x_sg_in199;
  wire [1:0] _add_all_x_sg_in200;
  wire [1:0] _add_all_x_sg_in201;
  wire [1:0] _add_all_x_sg_in202;
  wire [1:0] _add_all_x_sg_in203;
  wire [1:0] _add_all_x_sg_in204;
  wire [1:0] _add_all_x_sg_in205;
  wire [1:0] _add_all_x_sg_in206;
  wire [1:0] _add_all_x_sg_in207;
  wire [1:0] _add_all_x_sg_in208;
  wire [1:0] _add_all_x_sg_in209;
  wire [1:0] _add_all_x_sg_in210;
  wire [1:0] _add_all_x_sg_in211;
  wire [1:0] _add_all_x_sg_in212;
  wire [1:0] _add_all_x_sg_in213;
  wire [1:0] _add_all_x_sg_in214;
  wire [1:0] _add_all_x_sg_in215;
  wire [1:0] _add_all_x_sg_in216;
  wire [1:0] _add_all_x_sg_in217;
  wire [1:0] _add_all_x_sg_in218;
  wire [1:0] _add_all_x_sg_in219;
  wire [1:0] _add_all_x_sg_in220;
  wire [1:0] _add_all_x_sg_in221;
  wire [1:0] _add_all_x_sg_in222;
  wire [1:0] _add_all_x_sg_in225;
  wire [1:0] _add_all_x_sg_in226;
  wire [1:0] _add_all_x_sg_in227;
  wire [1:0] _add_all_x_sg_in228;
  wire [1:0] _add_all_x_sg_in229;
  wire [1:0] _add_all_x_sg_in230;
  wire [1:0] _add_all_x_sg_in231;
  wire [1:0] _add_all_x_sg_in232;
  wire [1:0] _add_all_x_sg_in233;
  wire [1:0] _add_all_x_sg_in234;
  wire [1:0] _add_all_x_sg_in235;
  wire [1:0] _add_all_x_sg_in236;
  wire [1:0] _add_all_x_sg_in237;
  wire [1:0] _add_all_x_sg_in238;
  wire [1:0] _add_all_x_sg_in239;
  wire [1:0] _add_all_x_sg_in240;
  wire [1:0] _add_all_x_sg_in241;
  wire [1:0] _add_all_x_sg_in242;
  wire [1:0] _add_all_x_sg_in243;
  wire [1:0] _add_all_x_sg_in244;
  wire [1:0] _add_all_x_sg_in245;
  wire [1:0] _add_all_x_sg_in246;
  wire [1:0] _add_all_x_sg_in247;
  wire [1:0] _add_all_x_sg_in248;
  wire [1:0] _add_all_x_sg_in249;
  wire [1:0] _add_all_x_sg_in250;
  wire [1:0] _add_all_x_sg_in251;
  wire [1:0] _add_all_x_sg_in252;
  wire [1:0] _add_all_x_sg_in253;
  wire [1:0] _add_all_x_sg_in254;
  wire [1:0] _add_all_x_sg_in257;
  wire [1:0] _add_all_x_sg_in258;
  wire [1:0] _add_all_x_sg_in259;
  wire [1:0] _add_all_x_sg_in260;
  wire [1:0] _add_all_x_sg_in261;
  wire [1:0] _add_all_x_sg_in262;
  wire [1:0] _add_all_x_sg_in263;
  wire [1:0] _add_all_x_sg_in264;
  wire [1:0] _add_all_x_sg_in265;
  wire [1:0] _add_all_x_sg_in266;
  wire [1:0] _add_all_x_sg_in267;
  wire [1:0] _add_all_x_sg_in268;
  wire [1:0] _add_all_x_sg_in269;
  wire [1:0] _add_all_x_sg_in270;
  wire [1:0] _add_all_x_sg_in271;
  wire [1:0] _add_all_x_sg_in272;
  wire [1:0] _add_all_x_sg_in273;
  wire [1:0] _add_all_x_sg_in274;
  wire [1:0] _add_all_x_sg_in275;
  wire [1:0] _add_all_x_sg_in276;
  wire [1:0] _add_all_x_sg_in277;
  wire [1:0] _add_all_x_sg_in278;
  wire [1:0] _add_all_x_sg_in279;
  wire [1:0] _add_all_x_sg_in280;
  wire [1:0] _add_all_x_sg_in281;
  wire [1:0] _add_all_x_sg_in282;
  wire [1:0] _add_all_x_sg_in283;
  wire [1:0] _add_all_x_sg_in284;
  wire [1:0] _add_all_x_sg_in285;
  wire [1:0] _add_all_x_sg_in286;
  wire [1:0] _add_all_x_sg_in289;
  wire [1:0] _add_all_x_sg_in290;
  wire [1:0] _add_all_x_sg_in291;
  wire [1:0] _add_all_x_sg_in292;
  wire [1:0] _add_all_x_sg_in293;
  wire [1:0] _add_all_x_sg_in294;
  wire [1:0] _add_all_x_sg_in295;
  wire [1:0] _add_all_x_sg_in296;
  wire [1:0] _add_all_x_sg_in297;
  wire [1:0] _add_all_x_sg_in298;
  wire [1:0] _add_all_x_sg_in299;
  wire [1:0] _add_all_x_sg_in300;
  wire [1:0] _add_all_x_sg_in301;
  wire [1:0] _add_all_x_sg_in302;
  wire [1:0] _add_all_x_sg_in303;
  wire [1:0] _add_all_x_sg_in304;
  wire [1:0] _add_all_x_sg_in305;
  wire [1:0] _add_all_x_sg_in306;
  wire [1:0] _add_all_x_sg_in307;
  wire [1:0] _add_all_x_sg_in308;
  wire [1:0] _add_all_x_sg_in309;
  wire [1:0] _add_all_x_sg_in310;
  wire [1:0] _add_all_x_sg_in311;
  wire [1:0] _add_all_x_sg_in312;
  wire [1:0] _add_all_x_sg_in313;
  wire [1:0] _add_all_x_sg_in314;
  wire [1:0] _add_all_x_sg_in315;
  wire [1:0] _add_all_x_sg_in316;
  wire [1:0] _add_all_x_sg_in317;
  wire [1:0] _add_all_x_sg_in318;
  wire [1:0] _add_all_x_sg_in321;
  wire [1:0] _add_all_x_sg_in322;
  wire [1:0] _add_all_x_sg_in323;
  wire [1:0] _add_all_x_sg_in324;
  wire [1:0] _add_all_x_sg_in325;
  wire [1:0] _add_all_x_sg_in326;
  wire [1:0] _add_all_x_sg_in327;
  wire [1:0] _add_all_x_sg_in328;
  wire [1:0] _add_all_x_sg_in329;
  wire [1:0] _add_all_x_sg_in330;
  wire [1:0] _add_all_x_sg_in331;
  wire [1:0] _add_all_x_sg_in332;
  wire [1:0] _add_all_x_sg_in333;
  wire [1:0] _add_all_x_sg_in334;
  wire [1:0] _add_all_x_sg_in335;
  wire [1:0] _add_all_x_sg_in336;
  wire [1:0] _add_all_x_sg_in337;
  wire [1:0] _add_all_x_sg_in338;
  wire [1:0] _add_all_x_sg_in339;
  wire [1:0] _add_all_x_sg_in340;
  wire [1:0] _add_all_x_sg_in341;
  wire [1:0] _add_all_x_sg_in342;
  wire [1:0] _add_all_x_sg_in343;
  wire [1:0] _add_all_x_sg_in344;
  wire [1:0] _add_all_x_sg_in345;
  wire [1:0] _add_all_x_sg_in346;
  wire [1:0] _add_all_x_sg_in347;
  wire [1:0] _add_all_x_sg_in348;
  wire [1:0] _add_all_x_sg_in349;
  wire [1:0] _add_all_x_sg_in350;
  wire [1:0] _add_all_x_sg_in353;
  wire [1:0] _add_all_x_sg_in354;
  wire [1:0] _add_all_x_sg_in355;
  wire [1:0] _add_all_x_sg_in356;
  wire [1:0] _add_all_x_sg_in357;
  wire [1:0] _add_all_x_sg_in358;
  wire [1:0] _add_all_x_sg_in359;
  wire [1:0] _add_all_x_sg_in360;
  wire [1:0] _add_all_x_sg_in361;
  wire [1:0] _add_all_x_sg_in362;
  wire [1:0] _add_all_x_sg_in363;
  wire [1:0] _add_all_x_sg_in364;
  wire [1:0] _add_all_x_sg_in365;
  wire [1:0] _add_all_x_sg_in366;
  wire [1:0] _add_all_x_sg_in367;
  wire [1:0] _add_all_x_sg_in368;
  wire [1:0] _add_all_x_sg_in369;
  wire [1:0] _add_all_x_sg_in370;
  wire [1:0] _add_all_x_sg_in371;
  wire [1:0] _add_all_x_sg_in372;
  wire [1:0] _add_all_x_sg_in373;
  wire [1:0] _add_all_x_sg_in374;
  wire [1:0] _add_all_x_sg_in375;
  wire [1:0] _add_all_x_sg_in376;
  wire [1:0] _add_all_x_sg_in377;
  wire [1:0] _add_all_x_sg_in378;
  wire [1:0] _add_all_x_sg_in379;
  wire [1:0] _add_all_x_sg_in380;
  wire [1:0] _add_all_x_sg_in381;
  wire [1:0] _add_all_x_sg_in382;
  wire [1:0] _add_all_x_sg_in385;
  wire [1:0] _add_all_x_sg_in386;
  wire [1:0] _add_all_x_sg_in387;
  wire [1:0] _add_all_x_sg_in388;
  wire [1:0] _add_all_x_sg_in389;
  wire [1:0] _add_all_x_sg_in390;
  wire [1:0] _add_all_x_sg_in391;
  wire [1:0] _add_all_x_sg_in392;
  wire [1:0] _add_all_x_sg_in393;
  wire [1:0] _add_all_x_sg_in394;
  wire [1:0] _add_all_x_sg_in395;
  wire [1:0] _add_all_x_sg_in396;
  wire [1:0] _add_all_x_sg_in397;
  wire [1:0] _add_all_x_sg_in398;
  wire [1:0] _add_all_x_sg_in399;
  wire [1:0] _add_all_x_sg_in400;
  wire [1:0] _add_all_x_sg_in401;
  wire [1:0] _add_all_x_sg_in402;
  wire [1:0] _add_all_x_sg_in403;
  wire [1:0] _add_all_x_sg_in404;
  wire [1:0] _add_all_x_sg_in405;
  wire [1:0] _add_all_x_sg_in406;
  wire [1:0] _add_all_x_sg_in407;
  wire [1:0] _add_all_x_sg_in408;
  wire [1:0] _add_all_x_sg_in409;
  wire [1:0] _add_all_x_sg_in410;
  wire [1:0] _add_all_x_sg_in411;
  wire [1:0] _add_all_x_sg_in412;
  wire [1:0] _add_all_x_sg_in413;
  wire [1:0] _add_all_x_sg_in414;
  wire [1:0] _add_all_x_sg_in417;
  wire [1:0] _add_all_x_sg_in418;
  wire [1:0] _add_all_x_sg_in419;
  wire [1:0] _add_all_x_sg_in420;
  wire [1:0] _add_all_x_sg_in421;
  wire [1:0] _add_all_x_sg_in422;
  wire [1:0] _add_all_x_sg_in423;
  wire [1:0] _add_all_x_sg_in424;
  wire [1:0] _add_all_x_sg_in425;
  wire [1:0] _add_all_x_sg_in426;
  wire [1:0] _add_all_x_sg_in427;
  wire [1:0] _add_all_x_sg_in428;
  wire [1:0] _add_all_x_sg_in429;
  wire [1:0] _add_all_x_sg_in430;
  wire [1:0] _add_all_x_sg_in431;
  wire [1:0] _add_all_x_sg_in432;
  wire [1:0] _add_all_x_sg_in433;
  wire [1:0] _add_all_x_sg_in434;
  wire [1:0] _add_all_x_sg_in435;
  wire [1:0] _add_all_x_sg_in436;
  wire [1:0] _add_all_x_sg_in437;
  wire [1:0] _add_all_x_sg_in438;
  wire [1:0] _add_all_x_sg_in439;
  wire [1:0] _add_all_x_sg_in440;
  wire [1:0] _add_all_x_sg_in441;
  wire [1:0] _add_all_x_sg_in442;
  wire [1:0] _add_all_x_sg_in443;
  wire [1:0] _add_all_x_sg_in444;
  wire [1:0] _add_all_x_sg_in445;
  wire [1:0] _add_all_x_sg_in446;
  wire [1:0] _add_all_x_sg_in449;
  wire [1:0] _add_all_x_sg_in450;
  wire [1:0] _add_all_x_sg_in451;
  wire [1:0] _add_all_x_sg_in452;
  wire [1:0] _add_all_x_sg_in453;
  wire [1:0] _add_all_x_sg_in454;
  wire [1:0] _add_all_x_sg_in455;
  wire [1:0] _add_all_x_sg_in456;
  wire [1:0] _add_all_x_sg_in457;
  wire [1:0] _add_all_x_sg_in458;
  wire [1:0] _add_all_x_sg_in459;
  wire [1:0] _add_all_x_sg_in460;
  wire [1:0] _add_all_x_sg_in461;
  wire [1:0] _add_all_x_sg_in462;
  wire [1:0] _add_all_x_sg_in463;
  wire [1:0] _add_all_x_sg_in464;
  wire [1:0] _add_all_x_sg_in465;
  wire [1:0] _add_all_x_sg_in466;
  wire [1:0] _add_all_x_sg_in467;
  wire [1:0] _add_all_x_sg_in468;
  wire [1:0] _add_all_x_sg_in469;
  wire [1:0] _add_all_x_sg_in470;
  wire [1:0] _add_all_x_sg_in471;
  wire [1:0] _add_all_x_sg_in472;
  wire [1:0] _add_all_x_sg_in473;
  wire [1:0] _add_all_x_sg_in474;
  wire [1:0] _add_all_x_sg_in475;
  wire [1:0] _add_all_x_sg_in476;
  wire [1:0] _add_all_x_sg_in477;
  wire [1:0] _add_all_x_sg_in478;
  wire [1:0] _add_all_x_sg_out33;
  wire [1:0] _add_all_x_sg_out34;
  wire [1:0] _add_all_x_sg_out35;
  wire [1:0] _add_all_x_sg_out36;
  wire [1:0] _add_all_x_sg_out37;
  wire [1:0] _add_all_x_sg_out38;
  wire [1:0] _add_all_x_sg_out39;
  wire [1:0] _add_all_x_sg_out40;
  wire [1:0] _add_all_x_sg_out41;
  wire [1:0] _add_all_x_sg_out42;
  wire [1:0] _add_all_x_sg_out43;
  wire [1:0] _add_all_x_sg_out44;
  wire [1:0] _add_all_x_sg_out45;
  wire [1:0] _add_all_x_sg_out46;
  wire [1:0] _add_all_x_sg_out47;
  wire [1:0] _add_all_x_sg_out48;
  wire [1:0] _add_all_x_sg_out49;
  wire [1:0] _add_all_x_sg_out50;
  wire [1:0] _add_all_x_sg_out51;
  wire [1:0] _add_all_x_sg_out52;
  wire [1:0] _add_all_x_sg_out53;
  wire [1:0] _add_all_x_sg_out54;
  wire [1:0] _add_all_x_sg_out55;
  wire [1:0] _add_all_x_sg_out56;
  wire [1:0] _add_all_x_sg_out57;
  wire [1:0] _add_all_x_sg_out58;
  wire [1:0] _add_all_x_sg_out59;
  wire [1:0] _add_all_x_sg_out60;
  wire [1:0] _add_all_x_sg_out61;
  wire [9:0] _add_all_x_sg_out62;
  wire [1:0] _add_all_x_sg_out65;
  wire [1:0] _add_all_x_sg_out66;
  wire [1:0] _add_all_x_sg_out67;
  wire [1:0] _add_all_x_sg_out68;
  wire [1:0] _add_all_x_sg_out69;
  wire [1:0] _add_all_x_sg_out70;
  wire [1:0] _add_all_x_sg_out71;
  wire [1:0] _add_all_x_sg_out72;
  wire [1:0] _add_all_x_sg_out73;
  wire [1:0] _add_all_x_sg_out74;
  wire [1:0] _add_all_x_sg_out75;
  wire [1:0] _add_all_x_sg_out76;
  wire [1:0] _add_all_x_sg_out77;
  wire [1:0] _add_all_x_sg_out78;
  wire [1:0] _add_all_x_sg_out79;
  wire [1:0] _add_all_x_sg_out80;
  wire [1:0] _add_all_x_sg_out81;
  wire [1:0] _add_all_x_sg_out82;
  wire [1:0] _add_all_x_sg_out83;
  wire [1:0] _add_all_x_sg_out84;
  wire [1:0] _add_all_x_sg_out85;
  wire [1:0] _add_all_x_sg_out86;
  wire [1:0] _add_all_x_sg_out87;
  wire [1:0] _add_all_x_sg_out88;
  wire [1:0] _add_all_x_sg_out89;
  wire [1:0] _add_all_x_sg_out90;
  wire [1:0] _add_all_x_sg_out91;
  wire [1:0] _add_all_x_sg_out92;
  wire [1:0] _add_all_x_sg_out93;
  wire [1:0] _add_all_x_sg_out94;
  wire [1:0] _add_all_x_sg_out97;
  wire [1:0] _add_all_x_sg_out98;
  wire [1:0] _add_all_x_sg_out99;
  wire [1:0] _add_all_x_sg_out100;
  wire [1:0] _add_all_x_sg_out101;
  wire [1:0] _add_all_x_sg_out102;
  wire [1:0] _add_all_x_sg_out103;
  wire [1:0] _add_all_x_sg_out104;
  wire [1:0] _add_all_x_sg_out105;
  wire [1:0] _add_all_x_sg_out106;
  wire [1:0] _add_all_x_sg_out107;
  wire [1:0] _add_all_x_sg_out108;
  wire [1:0] _add_all_x_sg_out109;
  wire [1:0] _add_all_x_sg_out110;
  wire [1:0] _add_all_x_sg_out111;
  wire [1:0] _add_all_x_sg_out112;
  wire [1:0] _add_all_x_sg_out113;
  wire [1:0] _add_all_x_sg_out114;
  wire [1:0] _add_all_x_sg_out115;
  wire [1:0] _add_all_x_sg_out116;
  wire [1:0] _add_all_x_sg_out117;
  wire [1:0] _add_all_x_sg_out118;
  wire [1:0] _add_all_x_sg_out119;
  wire [1:0] _add_all_x_sg_out120;
  wire [1:0] _add_all_x_sg_out121;
  wire [1:0] _add_all_x_sg_out122;
  wire [1:0] _add_all_x_sg_out123;
  wire [1:0] _add_all_x_sg_out124;
  wire [1:0] _add_all_x_sg_out125;
  wire [1:0] _add_all_x_sg_out126;
  wire [1:0] _add_all_x_sg_out129;
  wire [1:0] _add_all_x_sg_out130;
  wire [1:0] _add_all_x_sg_out131;
  wire [1:0] _add_all_x_sg_out132;
  wire [1:0] _add_all_x_sg_out133;
  wire [1:0] _add_all_x_sg_out134;
  wire [1:0] _add_all_x_sg_out135;
  wire [1:0] _add_all_x_sg_out136;
  wire [1:0] _add_all_x_sg_out137;
  wire [1:0] _add_all_x_sg_out138;
  wire [1:0] _add_all_x_sg_out139;
  wire [1:0] _add_all_x_sg_out140;
  wire [1:0] _add_all_x_sg_out141;
  wire [1:0] _add_all_x_sg_out142;
  wire [1:0] _add_all_x_sg_out143;
  wire [1:0] _add_all_x_sg_out144;
  wire [1:0] _add_all_x_sg_out145;
  wire [1:0] _add_all_x_sg_out146;
  wire [1:0] _add_all_x_sg_out147;
  wire [1:0] _add_all_x_sg_out148;
  wire [1:0] _add_all_x_sg_out149;
  wire [1:0] _add_all_x_sg_out150;
  wire [1:0] _add_all_x_sg_out151;
  wire [1:0] _add_all_x_sg_out152;
  wire [1:0] _add_all_x_sg_out153;
  wire [1:0] _add_all_x_sg_out154;
  wire [1:0] _add_all_x_sg_out155;
  wire [1:0] _add_all_x_sg_out156;
  wire [1:0] _add_all_x_sg_out157;
  wire [1:0] _add_all_x_sg_out158;
  wire [1:0] _add_all_x_sg_out161;
  wire [1:0] _add_all_x_sg_out162;
  wire [1:0] _add_all_x_sg_out163;
  wire [1:0] _add_all_x_sg_out164;
  wire [1:0] _add_all_x_sg_out165;
  wire [1:0] _add_all_x_sg_out166;
  wire [1:0] _add_all_x_sg_out167;
  wire [1:0] _add_all_x_sg_out168;
  wire [1:0] _add_all_x_sg_out169;
  wire [1:0] _add_all_x_sg_out170;
  wire [1:0] _add_all_x_sg_out171;
  wire [1:0] _add_all_x_sg_out172;
  wire [1:0] _add_all_x_sg_out173;
  wire [1:0] _add_all_x_sg_out174;
  wire [1:0] _add_all_x_sg_out175;
  wire [1:0] _add_all_x_sg_out176;
  wire [1:0] _add_all_x_sg_out177;
  wire [1:0] _add_all_x_sg_out178;
  wire [1:0] _add_all_x_sg_out179;
  wire [1:0] _add_all_x_sg_out180;
  wire [1:0] _add_all_x_sg_out181;
  wire [1:0] _add_all_x_sg_out182;
  wire [1:0] _add_all_x_sg_out183;
  wire [1:0] _add_all_x_sg_out184;
  wire [1:0] _add_all_x_sg_out185;
  wire [1:0] _add_all_x_sg_out186;
  wire [1:0] _add_all_x_sg_out187;
  wire [1:0] _add_all_x_sg_out188;
  wire [1:0] _add_all_x_sg_out189;
  wire [1:0] _add_all_x_sg_out190;
  wire [1:0] _add_all_x_sg_out193;
  wire [1:0] _add_all_x_sg_out194;
  wire [1:0] _add_all_x_sg_out195;
  wire [1:0] _add_all_x_sg_out196;
  wire [1:0] _add_all_x_sg_out197;
  wire [1:0] _add_all_x_sg_out198;
  wire [1:0] _add_all_x_sg_out199;
  wire [1:0] _add_all_x_sg_out200;
  wire [1:0] _add_all_x_sg_out201;
  wire [1:0] _add_all_x_sg_out202;
  wire [1:0] _add_all_x_sg_out203;
  wire [1:0] _add_all_x_sg_out204;
  wire [1:0] _add_all_x_sg_out205;
  wire [1:0] _add_all_x_sg_out206;
  wire [1:0] _add_all_x_sg_out207;
  wire [1:0] _add_all_x_sg_out208;
  wire [1:0] _add_all_x_sg_out209;
  wire [1:0] _add_all_x_sg_out210;
  wire [1:0] _add_all_x_sg_out211;
  wire [1:0] _add_all_x_sg_out212;
  wire [1:0] _add_all_x_sg_out213;
  wire [1:0] _add_all_x_sg_out214;
  wire [1:0] _add_all_x_sg_out215;
  wire [1:0] _add_all_x_sg_out216;
  wire [1:0] _add_all_x_sg_out217;
  wire [1:0] _add_all_x_sg_out218;
  wire [1:0] _add_all_x_sg_out219;
  wire [1:0] _add_all_x_sg_out220;
  wire [1:0] _add_all_x_sg_out221;
  wire [1:0] _add_all_x_sg_out222;
  wire [1:0] _add_all_x_sg_out225;
  wire [1:0] _add_all_x_sg_out226;
  wire [1:0] _add_all_x_sg_out227;
  wire [1:0] _add_all_x_sg_out228;
  wire [1:0] _add_all_x_sg_out229;
  wire [1:0] _add_all_x_sg_out230;
  wire [1:0] _add_all_x_sg_out231;
  wire [1:0] _add_all_x_sg_out232;
  wire [1:0] _add_all_x_sg_out233;
  wire [1:0] _add_all_x_sg_out234;
  wire [1:0] _add_all_x_sg_out235;
  wire [1:0] _add_all_x_sg_out236;
  wire [1:0] _add_all_x_sg_out237;
  wire [1:0] _add_all_x_sg_out238;
  wire [1:0] _add_all_x_sg_out239;
  wire [1:0] _add_all_x_sg_out240;
  wire [1:0] _add_all_x_sg_out241;
  wire [1:0] _add_all_x_sg_out242;
  wire [1:0] _add_all_x_sg_out243;
  wire [1:0] _add_all_x_sg_out244;
  wire [1:0] _add_all_x_sg_out245;
  wire [1:0] _add_all_x_sg_out246;
  wire [1:0] _add_all_x_sg_out247;
  wire [1:0] _add_all_x_sg_out248;
  wire [1:0] _add_all_x_sg_out249;
  wire [1:0] _add_all_x_sg_out250;
  wire [1:0] _add_all_x_sg_out251;
  wire [1:0] _add_all_x_sg_out252;
  wire [1:0] _add_all_x_sg_out253;
  wire [1:0] _add_all_x_sg_out254;
  wire [1:0] _add_all_x_sg_out257;
  wire [1:0] _add_all_x_sg_out258;
  wire [1:0] _add_all_x_sg_out259;
  wire [1:0] _add_all_x_sg_out260;
  wire [1:0] _add_all_x_sg_out261;
  wire [1:0] _add_all_x_sg_out262;
  wire [1:0] _add_all_x_sg_out263;
  wire [1:0] _add_all_x_sg_out264;
  wire [1:0] _add_all_x_sg_out265;
  wire [1:0] _add_all_x_sg_out266;
  wire [1:0] _add_all_x_sg_out267;
  wire [1:0] _add_all_x_sg_out268;
  wire [1:0] _add_all_x_sg_out269;
  wire [1:0] _add_all_x_sg_out270;
  wire [1:0] _add_all_x_sg_out271;
  wire [1:0] _add_all_x_sg_out272;
  wire [1:0] _add_all_x_sg_out273;
  wire [1:0] _add_all_x_sg_out274;
  wire [1:0] _add_all_x_sg_out275;
  wire [1:0] _add_all_x_sg_out276;
  wire [1:0] _add_all_x_sg_out277;
  wire [1:0] _add_all_x_sg_out278;
  wire [1:0] _add_all_x_sg_out279;
  wire [1:0] _add_all_x_sg_out280;
  wire [1:0] _add_all_x_sg_out281;
  wire [1:0] _add_all_x_sg_out282;
  wire [1:0] _add_all_x_sg_out283;
  wire [1:0] _add_all_x_sg_out284;
  wire [1:0] _add_all_x_sg_out285;
  wire [1:0] _add_all_x_sg_out286;
  wire [1:0] _add_all_x_sg_out289;
  wire [1:0] _add_all_x_sg_out290;
  wire [1:0] _add_all_x_sg_out291;
  wire [1:0] _add_all_x_sg_out292;
  wire [1:0] _add_all_x_sg_out293;
  wire [1:0] _add_all_x_sg_out294;
  wire [1:0] _add_all_x_sg_out295;
  wire [1:0] _add_all_x_sg_out296;
  wire [1:0] _add_all_x_sg_out297;
  wire [1:0] _add_all_x_sg_out298;
  wire [1:0] _add_all_x_sg_out299;
  wire [1:0] _add_all_x_sg_out300;
  wire [1:0] _add_all_x_sg_out301;
  wire [1:0] _add_all_x_sg_out302;
  wire [1:0] _add_all_x_sg_out303;
  wire [1:0] _add_all_x_sg_out304;
  wire [1:0] _add_all_x_sg_out305;
  wire [1:0] _add_all_x_sg_out306;
  wire [1:0] _add_all_x_sg_out307;
  wire [1:0] _add_all_x_sg_out308;
  wire [1:0] _add_all_x_sg_out309;
  wire [1:0] _add_all_x_sg_out310;
  wire [1:0] _add_all_x_sg_out311;
  wire [1:0] _add_all_x_sg_out312;
  wire [1:0] _add_all_x_sg_out313;
  wire [1:0] _add_all_x_sg_out314;
  wire [1:0] _add_all_x_sg_out315;
  wire [1:0] _add_all_x_sg_out316;
  wire [1:0] _add_all_x_sg_out317;
  wire [1:0] _add_all_x_sg_out318;
  wire [1:0] _add_all_x_sg_out321;
  wire [1:0] _add_all_x_sg_out322;
  wire [1:0] _add_all_x_sg_out323;
  wire [1:0] _add_all_x_sg_out324;
  wire [1:0] _add_all_x_sg_out325;
  wire [1:0] _add_all_x_sg_out326;
  wire [1:0] _add_all_x_sg_out327;
  wire [1:0] _add_all_x_sg_out328;
  wire [1:0] _add_all_x_sg_out329;
  wire [1:0] _add_all_x_sg_out330;
  wire [1:0] _add_all_x_sg_out331;
  wire [1:0] _add_all_x_sg_out332;
  wire [1:0] _add_all_x_sg_out333;
  wire [1:0] _add_all_x_sg_out334;
  wire [1:0] _add_all_x_sg_out335;
  wire [1:0] _add_all_x_sg_out336;
  wire [1:0] _add_all_x_sg_out337;
  wire [1:0] _add_all_x_sg_out338;
  wire [1:0] _add_all_x_sg_out339;
  wire [1:0] _add_all_x_sg_out340;
  wire [1:0] _add_all_x_sg_out341;
  wire [1:0] _add_all_x_sg_out342;
  wire [1:0] _add_all_x_sg_out343;
  wire [1:0] _add_all_x_sg_out344;
  wire [1:0] _add_all_x_sg_out345;
  wire [1:0] _add_all_x_sg_out346;
  wire [1:0] _add_all_x_sg_out347;
  wire [1:0] _add_all_x_sg_out348;
  wire [1:0] _add_all_x_sg_out349;
  wire [1:0] _add_all_x_sg_out350;
  wire [1:0] _add_all_x_sg_out353;
  wire [1:0] _add_all_x_sg_out354;
  wire [1:0] _add_all_x_sg_out355;
  wire [1:0] _add_all_x_sg_out356;
  wire [1:0] _add_all_x_sg_out357;
  wire [1:0] _add_all_x_sg_out358;
  wire [1:0] _add_all_x_sg_out359;
  wire [1:0] _add_all_x_sg_out360;
  wire [1:0] _add_all_x_sg_out361;
  wire [1:0] _add_all_x_sg_out362;
  wire [1:0] _add_all_x_sg_out363;
  wire [1:0] _add_all_x_sg_out364;
  wire [1:0] _add_all_x_sg_out365;
  wire [1:0] _add_all_x_sg_out366;
  wire [1:0] _add_all_x_sg_out367;
  wire [1:0] _add_all_x_sg_out368;
  wire [1:0] _add_all_x_sg_out369;
  wire [1:0] _add_all_x_sg_out370;
  wire [1:0] _add_all_x_sg_out371;
  wire [1:0] _add_all_x_sg_out372;
  wire [1:0] _add_all_x_sg_out373;
  wire [1:0] _add_all_x_sg_out374;
  wire [1:0] _add_all_x_sg_out375;
  wire [1:0] _add_all_x_sg_out376;
  wire [1:0] _add_all_x_sg_out377;
  wire [1:0] _add_all_x_sg_out378;
  wire [1:0] _add_all_x_sg_out379;
  wire [1:0] _add_all_x_sg_out380;
  wire [1:0] _add_all_x_sg_out381;
  wire [1:0] _add_all_x_sg_out382;
  wire [1:0] _add_all_x_sg_out385;
  wire [1:0] _add_all_x_sg_out386;
  wire [1:0] _add_all_x_sg_out387;
  wire [1:0] _add_all_x_sg_out388;
  wire [1:0] _add_all_x_sg_out389;
  wire [1:0] _add_all_x_sg_out390;
  wire [1:0] _add_all_x_sg_out391;
  wire [1:0] _add_all_x_sg_out392;
  wire [1:0] _add_all_x_sg_out393;
  wire [1:0] _add_all_x_sg_out394;
  wire [1:0] _add_all_x_sg_out395;
  wire [1:0] _add_all_x_sg_out396;
  wire [1:0] _add_all_x_sg_out397;
  wire [1:0] _add_all_x_sg_out398;
  wire [1:0] _add_all_x_sg_out399;
  wire [1:0] _add_all_x_sg_out400;
  wire [1:0] _add_all_x_sg_out401;
  wire [1:0] _add_all_x_sg_out402;
  wire [1:0] _add_all_x_sg_out403;
  wire [1:0] _add_all_x_sg_out404;
  wire [1:0] _add_all_x_sg_out405;
  wire [1:0] _add_all_x_sg_out406;
  wire [1:0] _add_all_x_sg_out407;
  wire [1:0] _add_all_x_sg_out408;
  wire [1:0] _add_all_x_sg_out409;
  wire [1:0] _add_all_x_sg_out410;
  wire [1:0] _add_all_x_sg_out411;
  wire [1:0] _add_all_x_sg_out412;
  wire [1:0] _add_all_x_sg_out413;
  wire [1:0] _add_all_x_sg_out414;
  wire [1:0] _add_all_x_sg_out417;
  wire [1:0] _add_all_x_sg_out418;
  wire [1:0] _add_all_x_sg_out419;
  wire [1:0] _add_all_x_sg_out420;
  wire [1:0] _add_all_x_sg_out421;
  wire [1:0] _add_all_x_sg_out422;
  wire [1:0] _add_all_x_sg_out423;
  wire [1:0] _add_all_x_sg_out424;
  wire [1:0] _add_all_x_sg_out425;
  wire [1:0] _add_all_x_sg_out426;
  wire [1:0] _add_all_x_sg_out427;
  wire [1:0] _add_all_x_sg_out428;
  wire [1:0] _add_all_x_sg_out429;
  wire [1:0] _add_all_x_sg_out430;
  wire [1:0] _add_all_x_sg_out431;
  wire [1:0] _add_all_x_sg_out432;
  wire [1:0] _add_all_x_sg_out433;
  wire [1:0] _add_all_x_sg_out434;
  wire [1:0] _add_all_x_sg_out435;
  wire [1:0] _add_all_x_sg_out436;
  wire [1:0] _add_all_x_sg_out437;
  wire [1:0] _add_all_x_sg_out438;
  wire [1:0] _add_all_x_sg_out439;
  wire [1:0] _add_all_x_sg_out440;
  wire [1:0] _add_all_x_sg_out441;
  wire [1:0] _add_all_x_sg_out442;
  wire [1:0] _add_all_x_sg_out443;
  wire [1:0] _add_all_x_sg_out444;
  wire [1:0] _add_all_x_sg_out445;
  wire [1:0] _add_all_x_sg_out446;
  wire [1:0] _add_all_x_sg_out449;
  wire [1:0] _add_all_x_sg_out450;
  wire [1:0] _add_all_x_sg_out451;
  wire [1:0] _add_all_x_sg_out452;
  wire [1:0] _add_all_x_sg_out453;
  wire [1:0] _add_all_x_sg_out454;
  wire [1:0] _add_all_x_sg_out455;
  wire [1:0] _add_all_x_sg_out456;
  wire [1:0] _add_all_x_sg_out457;
  wire [1:0] _add_all_x_sg_out458;
  wire [1:0] _add_all_x_sg_out459;
  wire [1:0] _add_all_x_sg_out460;
  wire [1:0] _add_all_x_sg_out461;
  wire [1:0] _add_all_x_sg_out462;
  wire [1:0] _add_all_x_sg_out463;
  wire [1:0] _add_all_x_sg_out464;
  wire [1:0] _add_all_x_sg_out465;
  wire [1:0] _add_all_x_sg_out466;
  wire [1:0] _add_all_x_sg_out467;
  wire [1:0] _add_all_x_sg_out468;
  wire [1:0] _add_all_x_sg_out469;
  wire [1:0] _add_all_x_sg_out470;
  wire [1:0] _add_all_x_sg_out471;
  wire [1:0] _add_all_x_sg_out472;
  wire [1:0] _add_all_x_sg_out473;
  wire [1:0] _add_all_x_sg_out474;
  wire [1:0] _add_all_x_sg_out475;
  wire [1:0] _add_all_x_sg_out476;
  wire [1:0] _add_all_x_sg_out477;
  wire [1:0] _add_all_x_sg_out478;
  wire _add_all_x_dig_t0;
  wire _add_all_x_dig_t1;
  wire _add_all_x_dig_t2;
  wire _add_all_x_dig_t3;
  wire _add_all_x_dig_t4;
  wire _add_all_x_dig_t5;
  wire _add_all_x_dig_t6;
  wire _add_all_x_dig_t7;
  wire _add_all_x_dig_t8;
  wire _add_all_x_dig_t9;
  wire _add_all_x_dig_t10;
  wire _add_all_x_dig_t11;
  wire _add_all_x_dig_t12;
  wire _add_all_x_dig_t13;
  wire _add_all_x_dig_t14;
  wire _add_all_x_dig_t15;
  wire _add_all_x_dig_t16;
  wire _add_all_x_dig_t17;
  wire _add_all_x_dig_t18;
  wire _add_all_x_dig_t19;
  wire _add_all_x_dig_t20;
  wire _add_all_x_dig_t21;
  wire _add_all_x_dig_t22;
  wire _add_all_x_dig_t23;
  wire _add_all_x_dig_t24;
  wire _add_all_x_dig_t25;
  wire _add_all_x_dig_t26;
  wire _add_all_x_dig_t27;
  wire _add_all_x_dig_t28;
  wire _add_all_x_dig_t29;
  wire _add_all_x_dig_t30;
  wire _add_all_x_dig_t31;
  wire _add_all_x_dig_t32;
  wire _add_all_x_dig_t33;
  wire _add_all_x_dig_t34;
  wire _add_all_x_dig_t35;
  wire _add_all_x_dig_t36;
  wire _add_all_x_dig_t37;
  wire _add_all_x_dig_t38;
  wire _add_all_x_dig_t39;
  wire _add_all_x_dig_t40;
  wire _add_all_x_dig_t41;
  wire _add_all_x_dig_t42;
  wire _add_all_x_dig_t43;
  wire _add_all_x_dig_t44;
  wire _add_all_x_dig_t45;
  wire _add_all_x_dig_t46;
  wire _add_all_x_dig_t47;
  wire _add_all_x_dig_t48;
  wire _add_all_x_dig_t49;
  wire _add_all_x_dig_t50;
  wire _add_all_x_dig_t51;
  wire _add_all_x_dig_t52;
  wire _add_all_x_dig_t53;
  wire _add_all_x_dig_t54;
  wire _add_all_x_dig_t55;
  wire _add_all_x_dig_t56;
  wire _add_all_x_dig_t57;
  wire _add_all_x_dig_t58;
  wire _add_all_x_dig_t59;
  wire _add_all_x_dig_t60;
  wire _add_all_x_dig_t61;
  wire _add_all_x_dig_t62;
  wire _add_all_x_dig_t63;
  wire _add_all_x_dig_t64;
  wire _add_all_x_dig_t65;
  wire _add_all_x_dig_t66;
  wire _add_all_x_dig_t67;
  wire _add_all_x_dig_t68;
  wire _add_all_x_dig_t69;
  wire _add_all_x_dig_t70;
  wire _add_all_x_dig_t71;
  wire _add_all_x_dig_t72;
  wire _add_all_x_dig_t73;
  wire _add_all_x_dig_t74;
  wire _add_all_x_dig_t75;
  wire _add_all_x_dig_t76;
  wire _add_all_x_dig_t77;
  wire _add_all_x_dig_t78;
  wire _add_all_x_dig_t79;
  wire _add_all_x_dig_t80;
  wire _add_all_x_dig_t81;
  wire _add_all_x_dig_t82;
  wire _add_all_x_dig_t83;
  wire _add_all_x_dig_t84;
  wire _add_all_x_dig_t85;
  wire _add_all_x_dig_t86;
  wire _add_all_x_dig_t87;
  wire _add_all_x_dig_t88;
  wire _add_all_x_dig_t89;
  wire _add_all_x_dig_t90;
  wire _add_all_x_dig_t91;
  wire _add_all_x_dig_t92;
  wire _add_all_x_dig_t93;
  wire _add_all_x_dig_t94;
  wire _add_all_x_dig_t95;
  wire _add_all_x_dig_t96;
  wire _add_all_x_dig_t97;
  wire _add_all_x_dig_t98;
  wire _add_all_x_dig_t99;
  wire _add_all_x_dig_t100;
  wire _add_all_x_dig_t101;
  wire _add_all_x_dig_t102;
  wire _add_all_x_dig_t103;
  wire _add_all_x_dig_t104;
  wire _add_all_x_dig_t105;
  wire _add_all_x_dig_t106;
  wire _add_all_x_dig_t107;
  wire _add_all_x_dig_t108;
  wire _add_all_x_dig_t109;
  wire _add_all_x_dig_t110;
  wire _add_all_x_dig_t111;
  wire _add_all_x_dig_t112;
  wire _add_all_x_dig_t113;
  wire _add_all_x_dig_t114;
  wire _add_all_x_dig_t115;
  wire _add_all_x_dig_t116;
  wire _add_all_x_dig_t117;
  wire _add_all_x_dig_t118;
  wire _add_all_x_dig_t119;
  wire _add_all_x_dig_t120;
  wire _add_all_x_dig_t121;
  wire _add_all_x_dig_t122;
  wire _add_all_x_dig_t123;
  wire _add_all_x_dig_t124;
  wire _add_all_x_dig_t125;
  wire _add_all_x_dig_t126;
  wire _add_all_x_dig_t127;
  wire _add_all_x_dig_t128;
  wire _add_all_x_dig_t129;
  wire _add_all_x_dig_t130;
  wire _add_all_x_dig_t131;
  wire _add_all_x_dig_t132;
  wire _add_all_x_dig_t133;
  wire _add_all_x_dig_t134;
  wire _add_all_x_dig_t135;
  wire _add_all_x_dig_t136;
  wire _add_all_x_dig_t137;
  wire _add_all_x_dig_t138;
  wire _add_all_x_dig_t139;
  wire _add_all_x_dig_t140;
  wire _add_all_x_dig_t141;
  wire _add_all_x_dig_t142;
  wire _add_all_x_dig_t143;
  wire _add_all_x_dig_t144;
  wire _add_all_x_dig_t145;
  wire _add_all_x_dig_t146;
  wire _add_all_x_dig_t147;
  wire _add_all_x_dig_t148;
  wire _add_all_x_dig_t149;
  wire _add_all_x_dig_t150;
  wire _add_all_x_dig_t151;
  wire _add_all_x_dig_t152;
  wire _add_all_x_dig_t153;
  wire _add_all_x_dig_t154;
  wire _add_all_x_dig_t155;
  wire _add_all_x_dig_t156;
  wire _add_all_x_dig_t157;
  wire _add_all_x_dig_t158;
  wire _add_all_x_dig_t159;
  wire _add_all_x_dig_t160;
  wire _add_all_x_dig_t161;
  wire _add_all_x_dig_t162;
  wire _add_all_x_dig_t163;
  wire _add_all_x_dig_t164;
  wire _add_all_x_dig_t165;
  wire _add_all_x_dig_t166;
  wire _add_all_x_dig_t167;
  wire _add_all_x_dig_t168;
  wire _add_all_x_dig_t169;
  wire _add_all_x_dig_t170;
  wire _add_all_x_dig_t171;
  wire _add_all_x_dig_t172;
  wire _add_all_x_dig_t173;
  wire _add_all_x_dig_t174;
  wire _add_all_x_dig_t175;
  wire _add_all_x_dig_t176;
  wire _add_all_x_dig_t177;
  wire _add_all_x_dig_t178;
  wire _add_all_x_dig_t179;
  wire _add_all_x_dig_t180;
  wire _add_all_x_dig_t181;
  wire _add_all_x_dig_t182;
  wire _add_all_x_dig_t183;
  wire _add_all_x_dig_t184;
  wire _add_all_x_dig_t185;
  wire _add_all_x_dig_t186;
  wire _add_all_x_dig_t187;
  wire _add_all_x_dig_t188;
  wire _add_all_x_dig_t189;
  wire _add_all_x_dig_t190;
  wire _add_all_x_dig_t191;
  wire _add_all_x_dig_t192;
  wire _add_all_x_dig_t193;
  wire _add_all_x_dig_t194;
  wire _add_all_x_dig_t195;
  wire _add_all_x_dig_t196;
  wire _add_all_x_dig_t197;
  wire _add_all_x_dig_t198;
  wire _add_all_x_dig_t199;
  wire _add_all_x_dig_t200;
  wire _add_all_x_dig_t201;
  wire _add_all_x_dig_t202;
  wire _add_all_x_dig_t203;
  wire _add_all_x_dig_t204;
  wire _add_all_x_dig_t205;
  wire _add_all_x_dig_t206;
  wire _add_all_x_dig_t207;
  wire _add_all_x_dig_t208;
  wire _add_all_x_dig_t209;
  wire _add_all_x_in_do;
  wire _add_all_x_out_do;
  wire _add_all_x_out_data;
  wire _add_all_x_p_reset;
  wire _add_all_x_m_clock;
  wire [9:0] _sub_x_data_in33;
  wire [9:0] _sub_x_data_in35;
  wire [9:0] _sub_x_data_in37;
  wire [9:0] _sub_x_data_in39;
  wire [9:0] _sub_x_data_in41;
  wire [9:0] _sub_x_data_in43;
  wire [9:0] _sub_x_data_in45;
  wire [9:0] _sub_x_data_in47;
  wire [9:0] _sub_x_data_in49;
  wire [9:0] _sub_x_data_in51;
  wire [9:0] _sub_x_data_in53;
  wire [9:0] _sub_x_data_in55;
  wire [9:0] _sub_x_data_in57;
  wire [9:0] _sub_x_data_in59;
  wire [9:0] _sub_x_data_in61;
  wire [9:0] _sub_x_data_in65;
  wire [9:0] _sub_x_data_in67;
  wire [9:0] _sub_x_data_in69;
  wire [9:0] _sub_x_data_in71;
  wire [9:0] _sub_x_data_in73;
  wire [9:0] _sub_x_data_in75;
  wire [9:0] _sub_x_data_in77;
  wire [9:0] _sub_x_data_in79;
  wire [9:0] _sub_x_data_in81;
  wire [9:0] _sub_x_data_in83;
  wire [9:0] _sub_x_data_in85;
  wire [9:0] _sub_x_data_in87;
  wire [9:0] _sub_x_data_in89;
  wire [9:0] _sub_x_data_in91;
  wire [9:0] _sub_x_data_in93;
  wire [9:0] _sub_x_data_in97;
  wire [9:0] _sub_x_data_in99;
  wire [9:0] _sub_x_data_in101;
  wire [9:0] _sub_x_data_in103;
  wire [9:0] _sub_x_data_in105;
  wire [9:0] _sub_x_data_in107;
  wire [9:0] _sub_x_data_in109;
  wire [9:0] _sub_x_data_in111;
  wire [9:0] _sub_x_data_in113;
  wire [9:0] _sub_x_data_in115;
  wire [9:0] _sub_x_data_in117;
  wire [9:0] _sub_x_data_in119;
  wire [9:0] _sub_x_data_in121;
  wire [9:0] _sub_x_data_in123;
  wire [9:0] _sub_x_data_in125;
  wire [9:0] _sub_x_data_in129;
  wire [9:0] _sub_x_data_in131;
  wire [9:0] _sub_x_data_in133;
  wire [9:0] _sub_x_data_in135;
  wire [9:0] _sub_x_data_in137;
  wire [9:0] _sub_x_data_in139;
  wire [9:0] _sub_x_data_in141;
  wire [9:0] _sub_x_data_in143;
  wire [9:0] _sub_x_data_in145;
  wire [9:0] _sub_x_data_in147;
  wire [9:0] _sub_x_data_in149;
  wire [9:0] _sub_x_data_in151;
  wire [9:0] _sub_x_data_in153;
  wire [9:0] _sub_x_data_in155;
  wire [9:0] _sub_x_data_in157;
  wire [9:0] _sub_x_data_in161;
  wire [9:0] _sub_x_data_in163;
  wire [9:0] _sub_x_data_in165;
  wire [9:0] _sub_x_data_in167;
  wire [9:0] _sub_x_data_in169;
  wire [9:0] _sub_x_data_in171;
  wire [9:0] _sub_x_data_in173;
  wire [9:0] _sub_x_data_in175;
  wire [9:0] _sub_x_data_in177;
  wire [9:0] _sub_x_data_in179;
  wire [9:0] _sub_x_data_in181;
  wire [9:0] _sub_x_data_in183;
  wire [9:0] _sub_x_data_in185;
  wire [9:0] _sub_x_data_in187;
  wire [9:0] _sub_x_data_in189;
  wire [9:0] _sub_x_data_in193;
  wire [9:0] _sub_x_data_in195;
  wire [9:0] _sub_x_data_in197;
  wire [9:0] _sub_x_data_in199;
  wire [9:0] _sub_x_data_in201;
  wire [9:0] _sub_x_data_in203;
  wire [9:0] _sub_x_data_in205;
  wire [9:0] _sub_x_data_in207;
  wire [9:0] _sub_x_data_in209;
  wire [9:0] _sub_x_data_in211;
  wire [9:0] _sub_x_data_in213;
  wire [9:0] _sub_x_data_in215;
  wire [9:0] _sub_x_data_in217;
  wire [9:0] _sub_x_data_in219;
  wire [9:0] _sub_x_data_in221;
  wire [9:0] _sub_x_data_in225;
  wire [9:0] _sub_x_data_in227;
  wire [9:0] _sub_x_data_in229;
  wire [9:0] _sub_x_data_in231;
  wire [9:0] _sub_x_data_in233;
  wire [9:0] _sub_x_data_in235;
  wire [9:0] _sub_x_data_in237;
  wire [9:0] _sub_x_data_in239;
  wire [9:0] _sub_x_data_in241;
  wire [9:0] _sub_x_data_in243;
  wire [9:0] _sub_x_data_in245;
  wire [9:0] _sub_x_data_in247;
  wire [9:0] _sub_x_data_in249;
  wire [9:0] _sub_x_data_in251;
  wire [9:0] _sub_x_data_in253;
  wire [9:0] _sub_x_data_in257;
  wire [9:0] _sub_x_data_in259;
  wire [9:0] _sub_x_data_in261;
  wire [9:0] _sub_x_data_in263;
  wire [9:0] _sub_x_data_in265;
  wire [9:0] _sub_x_data_in267;
  wire [9:0] _sub_x_data_in269;
  wire [9:0] _sub_x_data_in271;
  wire [9:0] _sub_x_data_in273;
  wire [9:0] _sub_x_data_in275;
  wire [9:0] _sub_x_data_in277;
  wire [9:0] _sub_x_data_in279;
  wire [9:0] _sub_x_data_in281;
  wire [9:0] _sub_x_data_in283;
  wire [9:0] _sub_x_data_in285;
  wire [9:0] _sub_x_data_in289;
  wire [9:0] _sub_x_data_in291;
  wire [9:0] _sub_x_data_in293;
  wire [9:0] _sub_x_data_in295;
  wire [9:0] _sub_x_data_in297;
  wire [9:0] _sub_x_data_in299;
  wire [9:0] _sub_x_data_in301;
  wire [9:0] _sub_x_data_in303;
  wire [9:0] _sub_x_data_in305;
  wire [9:0] _sub_x_data_in307;
  wire [9:0] _sub_x_data_in309;
  wire [9:0] _sub_x_data_in311;
  wire [9:0] _sub_x_data_in313;
  wire [9:0] _sub_x_data_in315;
  wire [9:0] _sub_x_data_in317;
  wire [9:0] _sub_x_data_in321;
  wire [9:0] _sub_x_data_in323;
  wire [9:0] _sub_x_data_in325;
  wire [9:0] _sub_x_data_in327;
  wire [9:0] _sub_x_data_in329;
  wire [9:0] _sub_x_data_in331;
  wire [9:0] _sub_x_data_in333;
  wire [9:0] _sub_x_data_in335;
  wire [9:0] _sub_x_data_in337;
  wire [9:0] _sub_x_data_in339;
  wire [9:0] _sub_x_data_in341;
  wire [9:0] _sub_x_data_in343;
  wire [9:0] _sub_x_data_in345;
  wire [9:0] _sub_x_data_in347;
  wire [9:0] _sub_x_data_in349;
  wire [9:0] _sub_x_data_in353;
  wire [9:0] _sub_x_data_in355;
  wire [9:0] _sub_x_data_in357;
  wire [9:0] _sub_x_data_in359;
  wire [9:0] _sub_x_data_in361;
  wire [9:0] _sub_x_data_in363;
  wire [9:0] _sub_x_data_in365;
  wire [9:0] _sub_x_data_in367;
  wire [9:0] _sub_x_data_in369;
  wire [9:0] _sub_x_data_in371;
  wire [9:0] _sub_x_data_in373;
  wire [9:0] _sub_x_data_in375;
  wire [9:0] _sub_x_data_in377;
  wire [9:0] _sub_x_data_in379;
  wire [9:0] _sub_x_data_in381;
  wire [9:0] _sub_x_data_in385;
  wire [9:0] _sub_x_data_in387;
  wire [9:0] _sub_x_data_in389;
  wire [9:0] _sub_x_data_in391;
  wire [9:0] _sub_x_data_in393;
  wire [9:0] _sub_x_data_in395;
  wire [9:0] _sub_x_data_in397;
  wire [9:0] _sub_x_data_in399;
  wire [9:0] _sub_x_data_in401;
  wire [9:0] _sub_x_data_in403;
  wire [9:0] _sub_x_data_in405;
  wire [9:0] _sub_x_data_in407;
  wire [9:0] _sub_x_data_in409;
  wire [9:0] _sub_x_data_in411;
  wire [9:0] _sub_x_data_in413;
  wire [9:0] _sub_x_data_in417;
  wire [9:0] _sub_x_data_in419;
  wire [9:0] _sub_x_data_in421;
  wire [9:0] _sub_x_data_in423;
  wire [9:0] _sub_x_data_in425;
  wire [9:0] _sub_x_data_in427;
  wire [9:0] _sub_x_data_in429;
  wire [9:0] _sub_x_data_in431;
  wire [9:0] _sub_x_data_in433;
  wire [9:0] _sub_x_data_in435;
  wire [9:0] _sub_x_data_in437;
  wire [9:0] _sub_x_data_in439;
  wire [9:0] _sub_x_data_in441;
  wire [9:0] _sub_x_data_in443;
  wire [9:0] _sub_x_data_in445;
  wire [9:0] _sub_x_data_in449;
  wire [9:0] _sub_x_data_in451;
  wire [9:0] _sub_x_data_in453;
  wire [9:0] _sub_x_data_in455;
  wire [9:0] _sub_x_data_in457;
  wire [9:0] _sub_x_data_in459;
  wire [9:0] _sub_x_data_in461;
  wire [9:0] _sub_x_data_in463;
  wire [9:0] _sub_x_data_in465;
  wire [9:0] _sub_x_data_in467;
  wire [9:0] _sub_x_data_in469;
  wire [9:0] _sub_x_data_in471;
  wire [9:0] _sub_x_data_in473;
  wire [9:0] _sub_x_data_in475;
  wire [9:0] _sub_x_data_in477;
  wire [9:0] _sub_x_data_in_index33;
  wire [9:0] _sub_x_data_in_index35;
  wire [9:0] _sub_x_data_in_index37;
  wire [9:0] _sub_x_data_in_index39;
  wire [9:0] _sub_x_data_in_index41;
  wire [9:0] _sub_x_data_in_index43;
  wire [9:0] _sub_x_data_in_index45;
  wire [9:0] _sub_x_data_in_index47;
  wire [9:0] _sub_x_data_in_index49;
  wire [9:0] _sub_x_data_in_index51;
  wire [9:0] _sub_x_data_in_index53;
  wire [9:0] _sub_x_data_in_index55;
  wire [9:0] _sub_x_data_in_index57;
  wire [9:0] _sub_x_data_in_index59;
  wire [9:0] _sub_x_data_in_index61;
  wire [9:0] _sub_x_data_in_index65;
  wire [9:0] _sub_x_data_in_index67;
  wire [9:0] _sub_x_data_in_index69;
  wire [9:0] _sub_x_data_in_index71;
  wire [9:0] _sub_x_data_in_index73;
  wire [9:0] _sub_x_data_in_index75;
  wire [9:0] _sub_x_data_in_index77;
  wire [9:0] _sub_x_data_in_index79;
  wire [9:0] _sub_x_data_in_index81;
  wire [9:0] _sub_x_data_in_index83;
  wire [9:0] _sub_x_data_in_index85;
  wire [9:0] _sub_x_data_in_index87;
  wire [9:0] _sub_x_data_in_index89;
  wire [9:0] _sub_x_data_in_index91;
  wire [9:0] _sub_x_data_in_index93;
  wire [9:0] _sub_x_data_in_index97;
  wire [9:0] _sub_x_data_in_index99;
  wire [9:0] _sub_x_data_in_index101;
  wire [9:0] _sub_x_data_in_index103;
  wire [9:0] _sub_x_data_in_index105;
  wire [9:0] _sub_x_data_in_index107;
  wire [9:0] _sub_x_data_in_index109;
  wire [9:0] _sub_x_data_in_index111;
  wire [9:0] _sub_x_data_in_index113;
  wire [9:0] _sub_x_data_in_index115;
  wire [9:0] _sub_x_data_in_index117;
  wire [9:0] _sub_x_data_in_index119;
  wire [9:0] _sub_x_data_in_index121;
  wire [9:0] _sub_x_data_in_index123;
  wire [9:0] _sub_x_data_in_index125;
  wire [9:0] _sub_x_data_in_index129;
  wire [9:0] _sub_x_data_in_index131;
  wire [9:0] _sub_x_data_in_index133;
  wire [9:0] _sub_x_data_in_index135;
  wire [9:0] _sub_x_data_in_index137;
  wire [9:0] _sub_x_data_in_index139;
  wire [9:0] _sub_x_data_in_index141;
  wire [9:0] _sub_x_data_in_index143;
  wire [9:0] _sub_x_data_in_index145;
  wire [9:0] _sub_x_data_in_index147;
  wire [9:0] _sub_x_data_in_index149;
  wire [9:0] _sub_x_data_in_index151;
  wire [9:0] _sub_x_data_in_index153;
  wire [9:0] _sub_x_data_in_index155;
  wire [9:0] _sub_x_data_in_index157;
  wire [9:0] _sub_x_data_in_index161;
  wire [9:0] _sub_x_data_in_index163;
  wire [9:0] _sub_x_data_in_index165;
  wire [9:0] _sub_x_data_in_index167;
  wire [9:0] _sub_x_data_in_index169;
  wire [9:0] _sub_x_data_in_index171;
  wire [9:0] _sub_x_data_in_index173;
  wire [9:0] _sub_x_data_in_index175;
  wire [9:0] _sub_x_data_in_index177;
  wire [9:0] _sub_x_data_in_index179;
  wire [9:0] _sub_x_data_in_index181;
  wire [9:0] _sub_x_data_in_index183;
  wire [9:0] _sub_x_data_in_index185;
  wire [9:0] _sub_x_data_in_index187;
  wire [9:0] _sub_x_data_in_index189;
  wire [9:0] _sub_x_data_in_index193;
  wire [9:0] _sub_x_data_in_index195;
  wire [9:0] _sub_x_data_in_index197;
  wire [9:0] _sub_x_data_in_index199;
  wire [9:0] _sub_x_data_in_index201;
  wire [9:0] _sub_x_data_in_index203;
  wire [9:0] _sub_x_data_in_index205;
  wire [9:0] _sub_x_data_in_index207;
  wire [9:0] _sub_x_data_in_index209;
  wire [9:0] _sub_x_data_in_index211;
  wire [9:0] _sub_x_data_in_index213;
  wire [9:0] _sub_x_data_in_index215;
  wire [9:0] _sub_x_data_in_index217;
  wire [9:0] _sub_x_data_in_index219;
  wire [9:0] _sub_x_data_in_index221;
  wire [9:0] _sub_x_data_in_index225;
  wire [9:0] _sub_x_data_in_index227;
  wire [9:0] _sub_x_data_in_index229;
  wire [9:0] _sub_x_data_in_index231;
  wire [9:0] _sub_x_data_in_index233;
  wire [9:0] _sub_x_data_in_index235;
  wire [9:0] _sub_x_data_in_index237;
  wire [9:0] _sub_x_data_in_index239;
  wire [9:0] _sub_x_data_in_index241;
  wire [9:0] _sub_x_data_in_index243;
  wire [9:0] _sub_x_data_in_index245;
  wire [9:0] _sub_x_data_in_index247;
  wire [9:0] _sub_x_data_in_index249;
  wire [9:0] _sub_x_data_in_index251;
  wire [9:0] _sub_x_data_in_index253;
  wire [9:0] _sub_x_data_in_index257;
  wire [9:0] _sub_x_data_in_index259;
  wire [9:0] _sub_x_data_in_index261;
  wire [9:0] _sub_x_data_in_index263;
  wire [9:0] _sub_x_data_in_index265;
  wire [9:0] _sub_x_data_in_index267;
  wire [9:0] _sub_x_data_in_index269;
  wire [9:0] _sub_x_data_in_index271;
  wire [9:0] _sub_x_data_in_index273;
  wire [9:0] _sub_x_data_in_index275;
  wire [9:0] _sub_x_data_in_index277;
  wire [9:0] _sub_x_data_in_index279;
  wire [9:0] _sub_x_data_in_index281;
  wire [9:0] _sub_x_data_in_index283;
  wire [9:0] _sub_x_data_in_index285;
  wire [9:0] _sub_x_data_in_index289;
  wire [9:0] _sub_x_data_in_index291;
  wire [9:0] _sub_x_data_in_index293;
  wire [9:0] _sub_x_data_in_index295;
  wire [9:0] _sub_x_data_in_index297;
  wire [9:0] _sub_x_data_in_index299;
  wire [9:0] _sub_x_data_in_index301;
  wire [9:0] _sub_x_data_in_index303;
  wire [9:0] _sub_x_data_in_index305;
  wire [9:0] _sub_x_data_in_index307;
  wire [9:0] _sub_x_data_in_index309;
  wire [9:0] _sub_x_data_in_index311;
  wire [9:0] _sub_x_data_in_index313;
  wire [9:0] _sub_x_data_in_index315;
  wire [9:0] _sub_x_data_in_index317;
  wire [9:0] _sub_x_data_in_index321;
  wire [9:0] _sub_x_data_in_index323;
  wire [9:0] _sub_x_data_in_index325;
  wire [9:0] _sub_x_data_in_index327;
  wire [9:0] _sub_x_data_in_index329;
  wire [9:0] _sub_x_data_in_index331;
  wire [9:0] _sub_x_data_in_index333;
  wire [9:0] _sub_x_data_in_index335;
  wire [9:0] _sub_x_data_in_index337;
  wire [9:0] _sub_x_data_in_index339;
  wire [9:0] _sub_x_data_in_index341;
  wire [9:0] _sub_x_data_in_index343;
  wire [9:0] _sub_x_data_in_index345;
  wire [9:0] _sub_x_data_in_index347;
  wire [9:0] _sub_x_data_in_index349;
  wire [9:0] _sub_x_data_in_index353;
  wire [9:0] _sub_x_data_in_index355;
  wire [9:0] _sub_x_data_in_index357;
  wire [9:0] _sub_x_data_in_index359;
  wire [9:0] _sub_x_data_in_index361;
  wire [9:0] _sub_x_data_in_index363;
  wire [9:0] _sub_x_data_in_index365;
  wire [9:0] _sub_x_data_in_index367;
  wire [9:0] _sub_x_data_in_index369;
  wire [9:0] _sub_x_data_in_index371;
  wire [9:0] _sub_x_data_in_index373;
  wire [9:0] _sub_x_data_in_index375;
  wire [9:0] _sub_x_data_in_index377;
  wire [9:0] _sub_x_data_in_index379;
  wire [9:0] _sub_x_data_in_index381;
  wire [9:0] _sub_x_data_in_index385;
  wire [9:0] _sub_x_data_in_index387;
  wire [9:0] _sub_x_data_in_index389;
  wire [9:0] _sub_x_data_in_index391;
  wire [9:0] _sub_x_data_in_index393;
  wire [9:0] _sub_x_data_in_index395;
  wire [9:0] _sub_x_data_in_index397;
  wire [9:0] _sub_x_data_in_index399;
  wire [9:0] _sub_x_data_in_index401;
  wire [9:0] _sub_x_data_in_index403;
  wire [9:0] _sub_x_data_in_index405;
  wire [9:0] _sub_x_data_in_index407;
  wire [9:0] _sub_x_data_in_index409;
  wire [9:0] _sub_x_data_in_index411;
  wire [9:0] _sub_x_data_in_index413;
  wire [9:0] _sub_x_data_in_index417;
  wire [9:0] _sub_x_data_in_index419;
  wire [9:0] _sub_x_data_in_index421;
  wire [9:0] _sub_x_data_in_index423;
  wire [9:0] _sub_x_data_in_index425;
  wire [9:0] _sub_x_data_in_index427;
  wire [9:0] _sub_x_data_in_index429;
  wire [9:0] _sub_x_data_in_index431;
  wire [9:0] _sub_x_data_in_index433;
  wire [9:0] _sub_x_data_in_index435;
  wire [9:0] _sub_x_data_in_index437;
  wire [9:0] _sub_x_data_in_index439;
  wire [9:0] _sub_x_data_in_index441;
  wire [9:0] _sub_x_data_in_index443;
  wire [9:0] _sub_x_data_in_index445;
  wire [9:0] _sub_x_data_in_index449;
  wire [9:0] _sub_x_data_in_index451;
  wire [9:0] _sub_x_data_in_index453;
  wire [9:0] _sub_x_data_in_index455;
  wire [9:0] _sub_x_data_in_index457;
  wire [9:0] _sub_x_data_in_index459;
  wire [9:0] _sub_x_data_in_index461;
  wire [9:0] _sub_x_data_in_index463;
  wire [9:0] _sub_x_data_in_index465;
  wire [9:0] _sub_x_data_in_index467;
  wire [9:0] _sub_x_data_in_index469;
  wire [9:0] _sub_x_data_in_index471;
  wire [9:0] _sub_x_data_in_index473;
  wire [9:0] _sub_x_data_in_index475;
  wire [9:0] _sub_x_data_in_index477;
  wire [9:0] _sub_x_sub_array_out;
  wire _sub_x_subs_exe;
  wire _sub_x_p_reset;
  wire _sub_x_m_clock;
  reg _reg_0;
  reg _reg_1;
  reg _reg_2;
  reg _reg_3;
  wire _net_4;
  wire _net_5;
  wire _net_6;
  wire _net_7;
  wire _net_8;
  wire _net_9;
  wire _net_10;
  wire _net_11;
  wire _net_12;
  wire _net_13;
  wire _net_14;
  wire _net_15;
  wire _net_16;
  wire _net_17;
  wire _net_18;
  wire _net_19;
  wire _net_20;
  wire _net_21;
  wire _net_22;
  wire _net_23;
  wire _net_24;
  wire _net_25;
  wire _net_26;
  wire _net_27;
  wire _net_28;
  wire _net_29;
  wire _net_30;
  wire _net_31;
  wire _net_32;
  wire _net_33;
  wire _net_34;
  wire _net_35;
  wire _net_36;
  wire _net_37;
  wire _net_38;
  wire _net_39;
  wire _net_40;
  wire _net_41;
  wire _net_42;
  wire _net_43;
  wire _net_44;
  wire _net_45;
  wire _net_46;
  wire _net_47;
  wire _net_48;
  wire _net_49;
  wire _net_50;
  wire _net_51;
  wire _net_52;
  wire _net_53;
  wire _net_54;
  wire _net_55;
  wire _net_56;
  wire _net_57;
  wire _net_58;
  wire _net_59;
  wire _net_60;
  wire _net_61;
  wire _net_62;
  wire _net_63;
  wire _net_64;
  wire _net_65;
  wire _net_66;
  wire _net_67;
  wire _net_68;
  wire _net_69;
  wire _net_70;
  wire _net_71;
  wire _net_72;
  wire _net_73;
  wire _net_74;
  wire _net_75;
  wire _net_76;
  wire _net_77;
  wire _net_78;
  wire _net_79;
  wire _net_80;
  wire _net_81;
  wire _net_82;
  wire _net_83;
  wire _net_84;
  wire _net_85;
  wire _net_86;
  wire _net_87;
  wire _net_88;
  wire _net_89;
  wire _net_90;
  wire _net_91;
  wire _net_92;
  wire _net_93;
  wire _net_94;
  wire _net_95;
  wire _net_96;
  wire _net_97;
  wire _net_98;
  wire _net_99;
  wire _net_100;
  wire _net_101;
  wire _net_102;
  wire _net_103;
  wire _net_104;
  wire _net_105;
  wire _net_106;
  wire _net_107;
  wire _net_108;
  wire _net_109;
  wire _net_110;
  wire _net_111;
  wire _net_112;
  wire _net_113;
  wire _net_114;
  wire _net_115;
  wire _net_116;
  wire _net_117;
  wire _net_118;
  wire _net_119;
  wire _net_120;
  wire _net_121;
  wire _net_122;
  wire _net_123;
  wire _net_124;
  wire _net_125;
  wire _net_126;
  wire _net_127;
  wire _net_128;
  wire _net_129;
  wire _net_130;
  wire _net_131;
  wire _net_132;
  wire _net_133;
  wire _net_134;
  wire _net_135;
  wire _net_136;
  wire _net_137;
  wire _net_138;
  wire _net_139;
  wire _net_140;
  wire _net_141;
  wire _net_142;
  wire _net_143;
  wire _net_144;
  wire _net_145;
  wire _net_146;
  wire _net_147;
  wire _net_148;
  wire _net_149;
  wire _net_150;
  wire _net_151;
  wire _net_152;
  wire _net_153;
  wire _net_154;
  wire _net_155;
  wire _net_156;
  wire _net_157;
  wire _net_158;
  wire _net_159;
  wire _net_160;
  wire _net_161;
  wire _net_162;
  wire _net_163;
  wire _net_164;
  wire _net_165;
  wire _net_166;
  wire _net_167;
  wire _net_168;
  wire _net_169;
  wire _net_170;
  wire _net_171;
  wire _net_172;
  wire _net_173;
  wire _net_174;
  wire _net_175;
  wire _net_176;
  wire _net_177;
  wire _net_178;
  wire _net_179;
  wire _net_180;
  wire _net_181;
  wire _net_182;
  wire _net_183;
  wire _net_184;
  wire _net_185;
  wire _net_186;
  wire _net_187;
  wire _net_188;
  wire _net_189;
  wire _net_190;
  wire _net_191;
  wire _net_192;
  wire _net_193;
  wire _net_194;
  wire _net_195;
  wire _net_196;
  wire _net_197;
  wire _net_198;
  wire _net_199;
  wire _net_200;
  wire _net_201;
  wire _net_202;
  wire _net_203;
  wire _net_204;
  wire _net_205;
  wire _net_206;
  wire _net_207;
  wire _net_208;
  wire _net_209;
  wire _net_210;
  wire _net_211;
  wire _net_212;
  wire _net_213;
  wire _net_214;
  wire _net_215;
  wire _net_216;
  wire _net_217;
  wire _net_218;
  wire _net_219;
  wire _net_220;
  wire _net_221;
  wire _net_222;
  wire _net_223;
  wire _net_224;
  wire _net_225;
  wire _net_226;
  wire _net_227;
  wire _net_228;
  wire _net_229;
  wire _net_230;
  wire _net_231;
  wire _net_232;
  wire _net_233;
  wire _net_234;
  wire _net_235;
  wire _net_236;
  wire _net_237;
  wire _net_238;
  wire _net_239;
  wire _net_240;
  wire _net_241;
  wire _net_242;
  wire _net_243;
  wire _net_244;
  wire _net_245;
  wire _net_246;
  wire _net_247;
  wire _net_248;
  wire _net_249;
  wire _net_250;
  wire _net_251;
  wire _net_252;
  wire _net_253;
  wire _net_254;
  wire _net_255;
  wire _net_256;
  wire _net_257;
  wire _net_258;
  wire _net_259;
  wire _net_260;
  wire _net_261;
  wire _net_262;
  wire _net_263;
  wire _net_264;
  wire _net_265;
  wire _net_266;
  wire _net_267;
  wire _net_268;
  wire _net_269;
  wire _net_270;
  wire _net_271;
  wire _net_272;
  wire _net_273;
  wire _net_274;
  wire _net_275;
  wire _net_276;
  wire _net_277;
  wire _net_278;
  wire _net_279;
  wire _net_280;
  wire _net_281;
  wire _net_282;
  wire _net_283;
  wire _net_284;
  wire _net_285;
  wire _net_286;
  wire _net_287;
  wire _net_288;
  wire _net_289;
  wire _net_290;
  wire _net_291;
  wire _net_292;
  wire _net_293;
  wire _net_294;
  wire _net_295;
  wire _net_296;
  wire _net_297;
  wire _net_298;
  wire _net_299;
  wire _net_300;
  wire _net_301;
  wire _net_302;
  wire _net_303;
  wire _net_304;
  wire _net_305;
  wire _net_306;
  wire _net_307;
  wire _net_308;
  wire _net_309;
  wire _net_310;
  wire _net_311;
  wire _net_312;
  wire _net_313;
  wire _net_314;
  wire _net_315;
  wire _net_316;
  wire _net_317;
  wire _net_318;
  wire _net_319;
  wire _net_320;
  wire _net_321;
  wire _net_322;
  wire _net_323;
  wire _net_324;
  wire _net_325;
  wire _net_326;
  wire _net_327;
  wire _net_328;
  wire _net_329;
  wire _net_330;
  wire _net_331;
  wire _net_332;
  wire _net_333;
  wire _net_334;
  wire _net_335;
  wire _net_336;
  wire _net_337;
  wire _net_338;
  wire _net_339;
  wire _net_340;
  wire _net_341;
  wire _net_342;
  wire _net_343;
  wire _net_344;
  wire _net_345;
  wire _net_346;
  wire _net_347;
  wire _net_348;
  wire _net_349;
  wire _net_350;
  wire _net_351;
  wire _net_352;
  wire _net_353;
  wire _net_354;
  wire _net_355;
  wire _net_356;
  wire _net_357;
  wire _net_358;
  wire _net_359;
  wire _net_360;
  wire _net_361;
  wire _net_362;
  wire _net_363;
  wire _net_364;
  wire _net_365;
  wire _net_366;
  wire _net_367;
  wire _net_368;
  wire _net_369;
  wire _net_370;
  wire _net_371;
  wire _net_372;
  wire _net_373;
  wire _net_374;
  wire _net_375;
  wire _net_376;
  wire _net_377;
  wire _net_378;
  wire _net_379;
  wire _net_380;
  wire _net_381;
  wire _net_382;
  wire _net_383;
  wire _net_384;
  wire _net_385;
  wire _net_386;
  wire _net_387;
  wire _net_388;
  wire _net_389;
  wire _net_390;
  wire _net_391;
  wire _net_392;
  wire _net_393;
  wire _net_394;
  wire _net_395;
  wire _net_396;
  wire _net_397;
  wire _net_398;
  wire _net_399;
  wire _net_400;
  wire _net_401;
  wire _net_402;
  wire _net_403;
  wire _net_404;
  wire _net_405;
  wire _net_406;
  wire _net_407;
  wire _net_408;
  wire _net_409;
  wire _net_410;
  wire _net_411;
  wire _net_412;
  wire _net_413;
  wire _net_414;
  wire _net_415;
  wire _net_416;
  wire _net_417;
  wire _net_418;
  wire _net_419;
  wire _net_420;
  wire _net_421;
  wire _net_422;
  wire _net_423;
  wire _net_424;
  wire _net_425;
  wire _net_426;
  wire _net_427;
  wire _net_428;
  wire _net_429;
  wire _net_430;
  wire _net_431;
  wire _net_432;
  wire _net_433;
  wire _net_434;
  wire _net_435;
  wire _net_436;
  wire _net_437;
  wire _net_438;
  wire _net_439;
  wire _net_440;
  wire _net_441;
  wire _net_442;
  wire _net_443;
  wire _net_444;
  wire _net_445;
  wire _net_446;
  wire _net_447;
  wire _net_448;
  wire _net_449;
  wire _net_450;
  wire _net_451;
  wire _net_452;
  wire _net_453;
  wire _net_454;
  wire _net_455;
  wire _net_456;
  wire _net_457;
  wire _net_458;
  wire _net_459;
  wire _net_460;
  wire _net_461;
  wire _net_462;
  wire _net_463;
  wire _net_464;
  wire _net_465;
  wire _net_466;
  wire _net_467;
  wire _net_468;
  wire _net_469;
  wire _net_470;
  wire _net_471;
  wire _net_472;
  wire _net_473;
  wire _net_474;
  wire _net_475;
  wire _net_476;
  wire _net_477;
  wire _net_478;
  wire _net_479;
  wire _net_480;
  wire _net_481;
  wire _net_482;
  wire _net_483;
  wire _net_484;
  wire _net_485;
  wire _net_486;
  wire _net_487;
  wire _net_488;
  wire _net_489;
  wire _net_490;
  wire _net_491;
  wire _net_492;
  wire _net_493;
  wire _net_494;
  wire _net_495;
  wire _net_496;
  wire _net_497;
  wire _net_498;
  wire _net_499;
  wire _net_500;
  wire _net_501;
  wire _net_502;
  wire _net_503;
  wire _net_504;
  wire _net_505;
  wire _net_506;
  wire _net_507;
  wire _net_508;
  wire _net_509;
  wire _net_510;
  wire _net_511;
  wire _net_512;
  wire _net_513;
  wire _net_514;
  wire _net_515;
  wire _net_516;
  wire _net_517;
  wire _net_518;
  wire _net_519;
  wire _net_520;
  wire _net_521;
  wire _net_522;
  wire _net_523;
  wire _net_524;
  wire _net_525;
  wire _net_526;
  wire _net_527;
  wire _net_528;
  wire _net_529;
  wire _net_530;
  wire _net_531;
  wire _net_532;
  wire _net_533;
  wire _net_534;
  wire _net_535;
  wire _net_536;
  wire _net_537;
  wire _net_538;
  wire _net_539;
  wire _net_540;
  wire _net_541;
  wire _net_542;
  wire _net_543;
  wire _net_544;
  wire _net_545;
  wire _net_546;
  wire _net_547;
  wire _net_548;
  wire _net_549;
  wire _net_550;
  wire _net_551;
  wire _net_552;
  wire _net_553;
  wire _net_554;
  wire _net_555;
  wire _net_556;
  wire _net_557;
  wire _net_558;
  wire _net_559;
  wire _net_560;
  wire _net_561;
  wire _net_562;
  wire _net_563;
  wire _net_564;
  wire _net_565;
  wire _net_566;
  wire _net_567;
  wire _net_568;
  wire _net_569;
  wire _net_570;
  wire _net_571;
  wire _net_572;
  wire _net_573;
  wire _net_574;
  wire _net_575;
  wire _net_576;
  wire _net_577;
  wire _net_578;
  wire _net_579;
  wire _net_580;
  wire _net_581;
  wire _net_582;
  wire _net_583;
  wire _net_584;
  wire _net_585;
  wire _net_586;
  wire _net_587;
  wire _net_588;
  wire _net_589;
  wire _net_590;
  wire _net_591;
  wire _net_592;
  wire _net_593;
  wire _net_594;
  wire _net_595;
  wire _net_596;
  wire _net_597;
  wire _net_598;
  wire _net_599;
  wire _net_600;
  wire _net_601;
  wire _net_602;
  wire _net_603;
  wire _net_604;
  wire _net_605;
  wire _net_606;
  wire _net_607;
  wire _net_608;
  wire _net_609;
  wire _net_610;
  wire _net_611;
  wire _net_612;
  wire _net_613;
  wire _net_614;
  wire _net_615;
  wire _net_616;
  wire _net_617;
  wire _net_618;
  wire _net_619;
  wire _net_620;
  wire _net_621;
  wire _net_622;
  wire _net_623;
  wire _net_624;
  wire _net_625;
  wire _net_626;
  wire _net_627;
  wire _net_628;
  wire _net_629;
  wire _net_630;
  wire _net_631;
  wire _net_632;
  wire _net_633;
  wire _net_634;
  wire _net_635;
  wire _net_636;
  wire _net_637;
  wire _net_638;
  wire _net_639;
  wire _net_640;
  wire _net_641;
  wire _net_642;
  wire _net_643;
  wire _net_644;
  wire _net_645;
  wire _net_646;
  wire _net_647;
  wire _net_648;
  wire _net_649;
  wire _net_650;
  wire _net_651;
  wire _net_652;
  wire _net_653;
  wire _net_654;
  wire _net_655;
  wire _net_656;
  wire _net_657;
  wire _net_658;
  wire _net_659;
  wire _net_660;
  wire _net_661;
  wire _net_662;
  wire _net_663;
  wire _net_664;
  wire _net_665;
  wire _net_666;
  wire _net_667;
  wire _net_668;
  wire _net_669;
  wire _net_670;
  wire _net_671;
  wire _net_672;
  wire _net_673;
  wire _net_674;
  wire _net_675;
  wire _net_676;
  wire _net_677;
  wire _net_678;
  wire _net_679;
  wire _net_680;
  wire _net_681;
  wire _net_682;
  wire _net_683;
  wire _net_684;
  wire _net_685;
  wire _net_686;
  wire _net_687;
  wire _net_688;
  wire _net_689;
  wire _net_690;
  wire _net_691;
  wire _net_692;
  wire _net_693;
  wire _net_694;
  wire _net_695;
  wire _net_696;
  wire _net_697;
  wire _net_698;
  wire _net_699;
  wire _net_700;
  wire _net_701;
  wire _net_702;
  wire _net_703;
  wire _net_704;
  wire _net_705;
  wire _net_706;
  wire _net_707;
  wire _net_708;
  wire _net_709;
  wire _net_710;
  wire _net_711;
  wire _net_712;
  wire _net_713;
  wire _net_714;
  wire _net_715;
  wire _net_716;
  wire _net_717;
  wire _net_718;
  wire _net_719;
  wire _net_720;
  wire _net_721;
  wire _net_722;
  wire _net_723;
  wire _net_724;
  wire _net_725;
  wire _net_726;
  wire _net_727;
  wire _net_728;
  wire _net_729;
  wire _net_730;
  wire _net_731;
  wire _net_732;
  wire _net_733;
  wire _net_734;
  wire _net_735;
  wire _net_736;
  wire _net_737;
  wire _net_738;
  wire _net_739;
  wire _net_740;
  wire _net_741;
  wire _net_742;
  wire _net_743;
  wire _net_744;
  wire _net_745;
  wire _net_746;
  wire _net_747;
  wire _net_748;
  wire _net_749;
  wire _net_750;
  wire _net_751;
  wire _net_752;
  wire _net_753;
  wire _net_754;
  wire _net_755;
  wire _net_756;
  wire _net_757;
  wire _net_758;
  wire _net_759;
  wire _net_760;
  wire _net_761;
  wire _net_762;
  wire _net_763;
  wire _net_764;
  wire _net_765;
  wire _net_766;
  wire _net_767;
  wire _net_768;
  wire _net_769;
  wire _net_770;
  wire _net_771;
  wire _net_772;
  wire _net_773;
  wire _net_774;
  wire _net_775;
  wire _net_776;
  wire _net_777;
  wire _net_778;
  wire _net_779;
  wire _net_780;
  wire _net_781;
  wire _net_782;
  wire _net_783;
  wire _net_784;
  wire _net_785;
  wire _net_786;
  wire _net_787;
  wire _net_788;
  wire _net_789;
  wire _net_790;
  wire _net_791;
  wire _net_792;
  wire _net_793;
  wire _net_794;
  wire _net_795;
  wire _net_796;
  wire _net_797;
  wire _net_798;
  wire _net_799;
  wire _net_800;
  wire _net_801;
  wire _net_802;
  wire _net_803;
  wire _net_804;
  wire _net_805;
  wire _net_806;
  wire _net_807;
  wire _net_808;
  wire _net_809;
  wire _net_810;
  wire _net_811;
  wire _net_812;
  wire _net_813;
  wire _net_814;
  wire _net_815;
  wire _net_816;
  wire _net_817;
  wire _net_818;
  wire _net_819;
  wire _net_820;
  wire _net_821;
  wire _net_822;
  wire _net_823;
  wire _net_824;
  wire _net_825;
  wire _net_826;
  wire _net_827;
  wire _net_828;
  wire _net_829;
  wire _net_830;
  wire _net_831;
  wire _net_832;
  wire _net_833;
  wire _net_834;
  wire _net_835;
  wire _net_836;
  wire _net_837;
  wire _net_838;
  wire _net_839;
  wire _net_840;
  wire _net_841;
  wire _net_842;
  wire _net_843;
  wire _net_844;
  wire _net_845;
  wire _net_846;
  wire _net_847;
  wire _net_848;
  wire _net_849;
  wire _net_850;
  wire _net_851;
  wire _net_852;
  wire _net_853;
  wire _net_854;
  wire _net_855;
  wire _net_856;
  wire _net_857;
  wire _net_858;
  wire _net_859;
  wire _net_860;
  wire _net_861;
  wire _net_862;
  wire _net_863;
  wire _net_864;
  wire _net_865;
  wire _net_866;
  wire _net_867;
  wire _net_868;
  wire _net_869;
  wire _net_870;
  wire _net_871;
  wire _net_872;
  wire _net_873;
  wire _net_874;
  wire _net_875;
  wire _net_876;
  wire _net_877;
  wire _net_878;
  wire _net_879;
  wire _net_880;
  wire _net_881;
  wire _net_882;
  wire _net_883;
  wire _net_884;
  wire _net_885;
  wire _net_886;
  wire _net_887;
  wire _net_888;
  wire _net_889;
  wire _net_890;
  wire _net_891;
  wire _net_892;
  wire _net_893;
  wire _net_894;
  wire _net_895;
  wire _net_896;
  wire _net_897;
  wire _net_898;
  wire _net_899;
  wire _net_900;
  wire _net_901;
  wire _net_902;
  wire _net_903;
  wire _net_904;
  wire _net_905;
  wire _net_906;
  wire _net_907;
  wire _net_908;
  wire _net_909;
  wire _net_910;
  wire _net_911;
  wire _net_912;
  wire _net_913;
  wire _net_914;
  wire _net_915;
  wire _net_916;
  wire _net_917;
  wire _net_918;
  wire _net_919;
  wire _net_920;
  wire _net_921;
  wire _net_922;
  wire _net_923;
  wire _net_924;
  wire _net_925;
  wire _net_926;
  wire _net_927;
  wire _net_928;
  wire _net_929;
  wire _net_930;
  wire _net_931;
  wire _net_932;
  wire _net_933;
  wire _net_934;
  wire _net_935;
  wire _net_936;
  wire _net_937;
  wire _net_938;
  wire _net_939;
  wire _net_940;
  wire _net_941;
  wire _net_942;
  wire _net_943;
  wire _net_944;
  wire _net_945;
  wire _net_946;
  wire _net_947;
  wire _net_948;
  wire _net_949;
  wire _net_950;
  wire _net_951;
  wire _net_952;
  wire _net_953;
  wire _net_954;
  wire _net_955;
  wire _net_956;
  wire _net_957;
  wire _net_958;
  wire _net_959;
  wire _net_960;
  wire _net_961;
  wire _net_962;
  wire _net_963;
  wire _net_964;
  wire _net_965;
  wire _net_966;
  wire _net_967;
  wire _net_968;
  wire _net_969;
  wire _net_970;
  wire _net_971;
  wire _net_972;
  wire _net_973;
  wire _net_974;
  wire _net_975;
  wire _net_976;
  wire _net_977;
  wire _net_978;
  wire _net_979;
  wire _net_980;
  wire _net_981;
  wire _net_982;
  wire _net_983;
  wire _net_984;
  wire _net_985;
  wire _net_986;
  wire _net_987;
  wire _net_988;
  wire _net_989;
  wire _net_990;
  wire _net_991;
  wire _net_992;
  wire _net_993;
  wire _net_994;
  wire _net_995;
  wire _net_996;
  wire _net_997;
  wire _net_998;
  wire _net_999;
  wire _net_1000;
  wire _net_1001;
  wire _net_1002;
  wire _net_1003;
  wire _net_1004;
  wire _net_1005;
  wire _net_1006;
  wire _net_1007;
  wire _net_1008;
  wire _net_1009;
  wire _net_1010;
  wire _net_1011;
  wire _net_1012;
  wire _net_1013;
  wire _net_1014;
  wire _net_1015;
  wire _net_1016;
  wire _net_1017;
  wire _net_1018;
  wire _net_1019;
  wire _net_1020;
  wire _net_1021;
  wire _net_1022;
  wire _net_1023;
  wire _net_1024;
  wire _net_1025;
  wire _net_1026;
  wire _net_1027;
  wire _net_1028;
  wire _net_1029;
  wire _net_1030;
  wire _net_1031;
  wire _net_1032;
  wire _net_1033;
  wire _net_1034;
  wire _net_1035;
  wire _net_1036;
  wire _net_1037;
  wire _net_1038;
  wire _net_1039;
  wire _net_1040;
  wire _net_1041;
  wire _net_1042;
  wire _net_1043;
  wire _net_1044;
  wire _net_1045;
  wire _net_1046;
  wire _net_1047;
  wire _net_1048;
  wire _net_1049;
  wire _net_1050;
  wire _net_1051;
  wire _net_1052;
  wire _net_1053;
  wire _net_1054;
  wire _net_1055;
  wire _net_1056;
  wire _net_1057;
  wire _net_1058;
  wire _net_1059;
  wire _net_1060;
  wire _net_1061;
  wire _net_1062;
  wire _net_1063;
  wire _net_1064;
  wire _net_1065;
  wire _net_1066;
  wire _net_1067;
  wire _net_1068;
  wire _net_1069;
  wire _net_1070;
  wire _net_1071;
  wire _net_1072;
  wire _net_1073;
  wire _net_1074;
  wire _net_1075;
  wire _net_1076;
  wire _net_1077;
  wire _net_1078;
  wire _net_1079;
  wire _net_1080;
  wire _net_1081;
  wire _net_1082;
  wire _net_1083;
  wire _net_1084;
  wire _net_1085;
  wire _net_1086;
  wire _net_1087;
  wire _net_1088;
  wire _net_1089;
  wire _net_1090;
  wire _net_1091;
  wire _net_1092;
  wire _net_1093;
  wire _net_1094;
  wire _net_1095;
  wire _net_1096;
  wire _net_1097;
  wire _net_1098;
  wire _net_1099;
  wire _net_1100;
  wire _net_1101;
  wire _net_1102;
  wire _net_1103;
  wire _net_1104;
  wire _net_1105;
  wire _net_1106;
  wire _net_1107;
  wire _net_1108;
  wire _net_1109;
  wire _net_1110;
  wire _net_1111;
  wire _net_1112;
  wire _net_1113;
  wire _net_1114;
  wire _net_1115;
  wire _net_1116;
  wire _net_1117;
  wire _net_1118;
  wire _net_1119;
  wire _net_1120;
  wire _net_1121;
  wire _net_1122;
  wire _net_1123;
  wire _net_1124;
  wire _net_1125;
  wire _net_1126;
  wire _net_1127;
  wire _net_1128;
  wire _net_1129;
  wire _net_1130;
  wire _net_1131;
  wire _net_1132;
  wire _net_1133;
  wire _net_1134;
  wire _net_1135;
  wire _net_1136;
  wire _net_1137;
  wire _net_1138;
  wire _net_1139;
  wire _net_1140;
  wire _net_1141;
  wire _net_1142;
  wire _net_1143;
  wire _net_1144;
  wire _net_1145;
  wire _net_1146;
  wire _net_1147;
  wire _net_1148;
  wire _net_1149;
  wire _net_1150;
  wire _net_1151;
  wire _net_1152;
  wire _net_1153;
  wire _net_1154;
  wire _net_1155;
  wire _net_1156;
  wire _net_1157;
  wire _net_1158;
  wire _net_1159;
  wire _net_1160;
  wire _net_1161;
  wire _net_1162;
  wire _net_1163;
  wire _net_1164;
  wire _net_1165;
  wire _net_1166;
  wire _net_1167;
  wire _net_1168;
  wire _net_1169;
  wire _net_1170;
  wire _net_1171;
  wire _net_1172;
  wire _net_1173;
  wire _net_1174;
  wire _net_1175;
  wire _net_1176;
  wire _net_1177;
  wire _net_1178;
  wire _net_1179;
  wire _net_1180;
  wire _net_1181;
  wire _net_1182;
  wire _net_1183;
  wire _net_1184;
  wire _net_1185;
  wire _net_1186;
  wire _net_1187;
  wire _net_1188;
  wire _net_1189;
  wire _net_1190;
  wire _net_1191;
  wire _net_1192;
  wire _net_1193;
  wire _net_1194;
  wire _net_1195;
  wire _net_1196;
  wire _net_1197;
  wire _net_1198;
  wire _net_1199;
  wire _net_1200;
  wire _net_1201;
  wire _net_1202;
  wire _net_1203;
  wire _net_1204;
  wire _net_1205;
  wire _net_1206;
  wire _net_1207;
  wire _net_1208;
  wire _net_1209;
  wire _net_1210;
  wire _net_1211;
  wire _net_1212;
  wire _net_1213;
  wire _net_1214;
  wire _net_1215;
  wire _net_1216;
  wire _net_1217;
  wire _net_1218;
  wire _net_1219;
  wire _net_1220;
  wire _net_1221;
  wire _net_1222;
  wire _net_1223;
  wire _net_1224;
  wire _net_1225;
  wire _net_1226;
  wire _net_1227;
  wire _net_1228;
  wire _net_1229;
  wire _net_1230;
  wire _net_1231;
  wire _net_1232;
  wire _net_1233;
  wire _net_1234;
  wire _net_1235;
  wire _net_1236;
  wire _net_1237;
  wire _net_1238;
  wire _net_1239;
  wire _net_1240;
  wire _net_1241;
  wire _net_1242;
  wire _net_1243;
  wire _net_1244;
  wire _net_1245;
  wire _net_1246;
  wire _net_1247;
  wire _net_1248;
  wire _net_1249;
  wire _net_1250;
  wire _net_1251;
  wire _net_1252;
  wire _net_1253;
  wire _net_1254;
  wire _net_1255;
  wire _net_1256;
  wire _net_1257;
  wire _net_1258;
  wire _net_1259;
  wire _net_1260;
  wire _net_1261;
  wire _net_1262;
  wire _net_1263;
  wire _net_1264;
  wire _net_1265;
  wire _net_1266;
  wire _net_1267;
  wire _net_1268;
  wire _net_1269;
  wire _net_1271;
  wire _reg_1_goto;
  wire _net_1272;
  wire _reg_2_goin;
  wire _net_1273;
  wire _net_1275;
  wire _net_1276;
  wire _net_1277;
  wire _net_1278;
  wire _net_1279;
  wire _net_1280;
  wire _net_1281;
  wire _net_1282;
  wire _net_1283;
  wire _net_1284;
  wire _net_1285;
  wire _net_1286;
  wire _net_1287;
  wire _net_1288;
  wire _net_1289;
  wire _net_1290;
  wire _net_1291;
  wire _net_1292;
  wire _net_1293;
  wire _net_1294;
  wire _net_1295;
  wire _net_1296;
  wire _net_1297;
  wire _net_1298;
  wire _net_1299;
  wire _net_1300;
  wire _net_1301;
  wire _net_1302;
  wire _net_1303;
  wire _net_1304;
  wire _net_1305;
  wire _net_1306;
  wire _net_1307;
  wire _net_1308;
  wire _net_1309;
  wire _net_1310;
  wire _net_1311;
  wire _net_1312;
  wire _net_1313;
  wire _net_1314;
  wire _net_1315;
  wire _net_1316;
  wire _net_1317;
  wire _net_1318;
  wire _net_1319;
  wire _net_1320;
  wire _net_1321;
  wire _net_1322;
  wire _net_1323;
  wire _net_1324;
  wire _net_1325;
  wire _net_1326;
  wire _net_1327;
  wire _net_1328;
  wire _net_1329;
  wire _net_1330;
  wire _net_1331;
  wire _net_1332;
  wire _net_1333;
  wire _net_1334;
  wire _net_1335;
  wire _net_1336;
  wire _net_1337;
  wire _net_1338;
  wire _net_1339;
  wire _net_1340;
  wire _net_1341;
  wire _net_1342;
  wire _net_1343;
  wire _net_1344;
  wire _net_1345;
  wire _net_1346;
  wire _net_1347;
  wire _net_1348;
  wire _net_1349;
  wire _net_1350;
  wire _net_1351;
  wire _net_1352;
  wire _net_1353;
  wire _net_1354;
  wire _net_1355;
  wire _net_1356;
  wire _net_1357;
  wire _net_1358;
  wire _net_1359;
  wire _net_1360;
  wire _net_1361;
  wire _net_1362;
  wire _net_1363;
  wire _net_1364;
  wire _net_1365;
  wire _net_1366;
  wire _net_1367;
  wire _net_1368;
  wire _net_1369;
  wire _net_1370;
  wire _net_1371;
  wire _net_1372;
  wire _net_1373;
  wire _net_1374;
  wire _net_1375;
  wire _net_1376;
  wire _net_1377;
  wire _net_1378;
  wire _net_1379;
  wire _net_1380;
  wire _net_1381;
  wire _net_1382;
  wire _net_1383;
  wire _net_1384;
  wire _net_1385;
  wire _net_1386;
  wire _net_1387;
  wire _net_1388;
  wire _net_1389;
  wire _net_1390;
  wire _net_1391;
  wire _net_1392;
  wire _net_1393;
  wire _net_1394;
  wire _net_1395;
  wire _net_1396;
  wire _net_1397;
  wire _net_1398;
  wire _net_1399;
  wire _net_1400;
  wire _net_1401;
  wire _net_1402;
  wire _net_1403;
  wire _net_1404;
  wire _net_1405;
  wire _net_1406;
  wire _net_1407;
  wire _net_1408;
  wire _net_1409;
  wire _net_1410;
  wire _net_1411;
  wire _net_1412;
  wire _net_1413;
  wire _net_1414;
  wire _net_1415;
  wire _net_1416;
  wire _net_1417;
  wire _net_1418;
  wire _net_1419;
  wire _net_1420;
  wire _net_1421;
  wire _net_1422;
  wire _net_1423;
  wire _net_1424;
  wire _net_1425;
  wire _net_1426;
  wire _net_1427;
  wire _net_1428;
  wire _net_1429;
  wire _net_1430;
  wire _net_1431;
  wire _net_1432;
  wire _net_1433;
  wire _net_1434;
  wire _net_1435;
  wire _net_1436;
  wire _net_1437;
  wire _net_1438;
  wire _net_1439;
  wire _net_1440;
  wire _net_1441;
  wire _net_1442;
  wire _net_1443;
  wire _net_1444;
  wire _net_1445;
  wire _net_1446;
  wire _net_1447;
  wire _net_1448;
  wire _net_1449;
  wire _net_1450;
  wire _net_1451;
  wire _net_1452;
  wire _net_1453;
  wire _net_1454;
  wire _net_1455;
  wire _net_1456;
  wire _net_1457;
  wire _net_1458;
  wire _net_1459;
  wire _net_1460;
  wire _net_1461;
  wire _net_1462;
  wire _net_1463;
  wire _net_1464;
  wire _net_1465;
  wire _net_1466;
  wire _net_1467;
  wire _net_1468;
  wire _net_1469;
  wire _net_1470;
  wire _net_1471;
  wire _net_1472;
  wire _net_1473;
  wire _net_1474;
  wire _net_1475;
  wire _net_1476;
  wire _net_1477;
  wire _net_1478;
  wire _net_1479;
  wire _net_1480;
  wire _net_1481;
  wire _net_1482;
  wire _net_1483;
  wire _net_1484;
  wire _net_1485;
  wire _net_1486;
  wire _net_1487;
  wire _net_1488;
  wire _net_1489;
  wire _net_1490;
  wire _net_1491;
  wire _net_1492;
  wire _net_1493;
  wire _net_1494;
  wire _net_1495;
  wire _net_1496;
  wire _net_1497;
  wire _net_1498;
  wire _net_1499;
  wire _net_1500;
  wire _net_1501;
  wire _net_1502;
  wire _net_1503;
  wire _net_1504;
  wire _net_1505;
  wire _net_1506;
  wire _net_1507;
  wire _net_1508;
  wire _net_1509;
  wire _net_1510;
  wire _net_1511;
  wire _net_1512;
  wire _net_1513;
  wire _net_1514;
  wire _net_1515;
  wire _net_1516;
  wire _net_1517;
  wire _net_1518;
  wire _net_1519;
  wire _net_1520;
  wire _net_1521;
  wire _net_1522;
  wire _net_1523;
  wire _net_1524;
  wire _net_1525;
  wire _net_1526;
  wire _net_1527;
  wire _net_1528;
  wire _net_1529;
  wire _net_1530;
  wire _net_1531;
  wire _net_1532;
  wire _net_1533;
  wire _net_1534;
  wire _net_1535;
  wire _net_1536;
  wire _net_1537;
  wire _net_1538;
  wire _net_1539;
  wire _net_1540;
  wire _net_1541;
  wire _net_1542;
  wire _net_1543;
  wire _net_1544;
  wire _net_1545;
  wire _net_1546;
  wire _net_1547;
  wire _net_1548;
  wire _net_1549;
  wire _net_1550;
  wire _net_1551;
  wire _net_1552;
  wire _net_1553;
  wire _net_1554;
  wire _net_1555;
  wire _net_1556;
  wire _net_1557;
  wire _net_1558;
  wire _net_1559;
  wire _net_1560;
  wire _net_1561;
  wire _net_1562;
  wire _net_1563;
  wire _net_1564;
  wire _net_1565;
  wire _net_1566;
  wire _net_1567;
  wire _net_1568;
  wire _net_1569;
  wire _net_1570;
  wire _net_1571;
  wire _net_1572;
  wire _net_1573;
  wire _net_1574;
  wire _net_1575;
  wire _net_1576;
  wire _net_1577;
  wire _net_1578;
  wire _net_1579;
  wire _net_1580;
  wire _net_1581;
  wire _net_1582;
  wire _net_1583;
  wire _net_1584;
  wire _net_1585;
  wire _net_1586;
  wire _net_1587;
  wire _net_1588;
  wire _net_1589;
  wire _net_1590;
  wire _net_1591;
  wire _net_1592;
  wire _net_1593;
  wire _net_1594;
  wire _net_1595;
  wire _net_1596;
  wire _net_1597;
  wire _net_1598;
  wire _net_1599;
  wire _net_1600;
  wire _net_1601;
  wire _net_1602;
  wire _net_1603;
  wire _net_1604;
  wire _net_1605;
  wire _net_1606;
  wire _net_1607;
  wire _net_1608;
  wire _net_1609;
  wire _net_1610;
  wire _net_1611;
  wire _net_1612;
  wire _net_1613;
  wire _net_1614;
  wire _net_1615;
  wire _net_1616;
  wire _net_1617;
  wire _net_1618;
  wire _net_1619;
  wire _net_1620;
  wire _net_1621;
  wire _net_1622;
  wire _net_1623;
  wire _net_1624;
  wire _net_1625;
  wire _net_1626;
  wire _net_1627;
  wire _net_1628;
  wire _net_1629;
  wire _net_1630;
  wire _net_1631;
  wire _net_1632;
  wire _net_1633;
  wire _net_1634;
  wire _net_1635;
  wire _net_1636;
  wire _net_1637;
  wire _net_1638;
  wire _net_1639;
  wire _net_1640;
  wire _net_1641;
  wire _net_1642;
  wire _net_1643;
  wire _net_1644;
  wire _net_1645;
  wire _net_1646;
  wire _net_1647;
  wire _net_1648;
  wire _net_1649;
  wire _net_1650;
  wire _net_1651;
  wire _net_1652;
  wire _net_1653;
  wire _net_1654;
  wire _net_1655;
  wire _net_1656;
  wire _net_1657;
  wire _net_1658;
  wire _net_1659;
  wire _net_1660;
  wire _net_1661;
  wire _net_1662;
  wire _net_1663;
  wire _net_1664;
  wire _net_1665;
  wire _net_1666;
  wire _net_1667;
  wire _net_1668;
  wire _net_1669;
  wire _net_1670;
  wire _net_1671;
  wire _net_1672;
  wire _net_1673;
  wire _net_1674;
  wire _net_1675;
  wire _net_1676;
  wire _net_1677;
  wire _net_1678;
  wire _net_1679;
  wire _net_1680;
  wire _net_1681;
  wire _net_1682;
  wire _net_1683;
  wire _net_1684;
  wire _net_1685;
  wire _net_1686;
  wire _net_1687;
  wire _net_1688;
  wire _net_1689;
  wire _net_1690;
  wire _net_1691;
  wire _net_1692;
  wire _net_1693;
  wire _net_1694;
  wire _net_1695;
  wire _net_1696;
  wire _net_1697;
  wire _net_1698;
  wire _net_1699;
  wire _net_1700;
  wire _net_1701;
  wire _net_1702;
  wire _net_1703;
  wire _net_1704;
  wire _net_1705;
  wire _net_1706;
  wire _net_1707;
  wire _net_1708;
  wire _net_1709;
  wire _net_1710;
  wire _net_1711;
  wire _net_1712;
  wire _net_1713;
  wire _net_1714;
  wire _net_1715;
  wire _net_1716;
  wire _net_1717;
  wire _net_1718;
  wire _net_1719;
  wire _net_1720;
  wire _net_1721;
  wire _net_1722;
  wire _net_1723;
  wire _net_1724;
  wire _net_1725;
  wire _net_1726;
  wire _net_1727;
  wire _net_1728;
  wire _net_1729;
  wire _net_1730;
  wire _net_1731;
  wire _net_1732;
  wire _net_1733;
  wire _net_1734;
  wire _net_1735;
  wire _net_1736;
  wire _net_1737;
  wire _net_1738;
  wire _net_1739;
  wire _net_1740;
  wire _net_1741;
  wire _net_1742;
  wire _net_1743;
  wire _net_1744;
  wire _net_1745;
  wire _net_1746;
  wire _net_1747;
  wire _net_1748;
  wire _net_1749;
  wire _net_1750;
  wire _net_1751;
  wire _net_1752;
  wire _net_1753;
  wire _net_1754;
  wire _net_1755;
  wire _net_1756;
  wire _net_1757;
  wire _net_1758;
  wire _net_1759;
  wire _net_1760;
  wire _net_1761;
  wire _net_1762;
  wire _net_1763;
  wire _net_1764;
  wire _net_1765;
  wire _net_1766;
  wire _net_1767;
  wire _net_1768;
  wire _net_1769;
  wire _net_1770;
  wire _net_1771;
  wire _net_1772;
  wire _net_1773;
  wire _net_1774;
  wire _net_1775;
  wire _net_1776;
  wire _net_1777;
  wire _net_1778;
  wire _net_1779;
  wire _net_1780;
  wire _net_1781;
  wire _net_1782;
  wire _net_1783;
  wire _net_1784;
  wire _net_1785;
  wire _net_1786;
  wire _net_1787;
  wire _net_1788;
  wire _net_1789;
  wire _net_1790;
  wire _net_1791;
  wire _net_1792;
  wire _net_1793;
  wire _net_1794;
  wire _net_1795;
  wire _net_1796;
  wire _net_1797;
  wire _net_1798;
  wire _net_1799;
  wire _net_1800;
  wire _net_1801;
  wire _net_1802;
  wire _net_1803;
  wire _net_1804;
  wire _net_1805;
  wire _net_1806;
  wire _net_1807;
  wire _net_1808;
  wire _net_1809;
  wire _net_1810;
  wire _net_1811;
  wire _net_1812;
  wire _net_1813;
  wire _net_1814;
  wire _net_1815;
  wire _net_1816;
  wire _net_1817;
  wire _net_1818;
  wire _net_1819;
  wire _net_1820;
  wire _net_1821;
  wire _net_1822;
  wire _net_1823;
  wire _net_1824;
  wire _net_1825;
  wire _net_1826;
  wire _net_1827;
  wire _net_1828;
  wire _net_1829;
  wire _net_1830;
  wire _net_1831;
  wire _net_1832;
  wire _net_1833;
  wire _net_1834;
  wire _net_1835;
  wire _net_1836;
  wire _net_1837;
  wire _net_1838;
  wire _net_1839;
  wire _net_1840;
  wire _net_1841;
  wire _net_1842;
  wire _net_1843;
  wire _net_1844;
  wire _net_1845;
  wire _net_1846;
  wire _net_1847;
  wire _net_1848;
  wire _net_1849;
  wire _net_1850;
  wire _net_1851;
  wire _net_1852;
  wire _net_1853;
  wire _net_1854;
  wire _net_1855;
  wire _net_1856;
  wire _net_1857;
  wire _net_1858;
  wire _net_1859;
  wire _net_1860;
  wire _net_1861;
  wire _net_1862;
  wire _net_1863;
  wire _net_1864;
  wire _net_1865;
  wire _net_1866;
  wire _net_1867;
  wire _net_1868;
  wire _net_1869;
  wire _net_1870;
  wire _net_1871;
  wire _net_1872;
  wire _net_1873;
  wire _net_1874;
  wire _net_1875;
  wire _net_1876;
  wire _net_1877;
  wire _net_1878;
  wire _net_1879;
  wire _net_1880;
  wire _net_1881;
  wire _net_1882;
  wire _net_1883;
  wire _net_1884;
  wire _net_1885;
  wire _net_1886;
  wire _net_1887;
  wire _net_1888;
  wire _net_1889;
  wire _net_1890;
  wire _net_1891;
  wire _net_1892;
  wire _net_1893;
  wire _net_1894;
  wire _net_1895;
  wire _net_1896;
  wire _net_1897;
  wire _net_1898;
  wire _net_1899;
  wire _net_1900;
  wire _net_1901;
  wire _net_1902;
  wire _net_1903;
  wire _net_1904;
  wire _net_1905;
  wire _net_1906;
  wire _net_1907;
  wire _net_1908;
  wire _net_1909;
  wire _net_1910;
  wire _net_1911;
  wire _net_1912;
  wire _net_1913;
  wire _net_1914;
  wire _net_1915;
  wire _net_1916;
  wire _net_1917;
  wire _net_1918;
  wire _net_1919;
  wire _net_1920;
  wire _net_1921;
  wire _net_1922;
  wire _net_1923;
  wire _net_1924;
  wire _net_1925;
  wire _net_1926;
  wire _net_1927;
  wire _net_1928;
  wire _net_1929;
  wire _net_1930;
  wire _net_1931;
  wire _net_1932;
  wire _net_1933;
  wire _net_1934;
  wire _net_1935;
  wire _net_1936;
  wire _net_1937;
  wire _net_1938;
  wire _net_1939;
  wire _net_1940;
  wire _net_1941;
  wire _net_1942;
  wire _net_1943;
  wire _net_1944;
  wire _net_1945;
  wire _net_1946;
  wire _net_1947;
  wire _net_1948;
  wire _net_1949;
  wire _net_1950;
  wire _net_1951;
  wire _net_1952;
  wire _net_1953;
  wire _net_1954;
  wire _net_1955;
  wire _net_1956;
  wire _net_1957;
  wire _net_1958;
  wire _net_1959;
  wire _net_1960;
  wire _net_1961;
  wire _net_1962;
  wire _net_1963;
  wire _net_1964;
  wire _net_1965;
  wire _net_1966;
  wire _net_1967;
  wire _net_1968;
  wire _net_1969;
  wire _net_1970;
  wire _net_1971;
  wire _net_1972;
  wire _net_1973;
  wire _net_1974;
  wire _net_1975;
  wire _net_1976;
  wire _net_1977;
  wire _net_1978;
  wire _net_1979;
  wire _net_1980;
  wire _net_1981;
  wire _net_1982;
  wire _net_1983;
  wire _net_1984;
  wire _net_1985;
  wire _net_1986;
  wire _net_1987;
  wire _net_1988;
  wire _net_1989;
  wire _net_1990;
  wire _net_1991;
  wire _net_1992;
  wire _net_1993;
  wire _net_1994;
  wire _net_1995;
  wire _net_1996;
  wire _net_1997;
  wire _net_1998;
  wire _net_1999;
  wire _net_2000;
  wire _net_2001;
  wire _net_2002;
  wire _net_2003;
  wire _net_2004;
  wire _net_2005;
  wire _net_2006;
  wire _net_2007;
  wire _net_2008;
  wire _net_2009;
  wire _net_2010;
  wire _net_2011;
  wire _net_2012;
  wire _net_2013;
  wire _net_2014;
  wire _net_2015;
  wire _net_2016;
  wire _net_2017;
  wire _net_2018;
  wire _net_2019;
  wire _net_2020;
  wire _net_2021;
  wire _net_2022;
  wire _net_2023;
  wire _net_2024;
  wire _net_2025;
  wire _net_2026;
  wire _net_2027;
  wire _net_2028;
  wire _net_2029;
  wire _net_2030;
  wire _net_2031;
  wire _net_2032;
  wire _net_2033;
  wire _net_2034;
  wire _net_2035;
  wire _net_2036;
  wire _net_2037;
  wire _net_2038;
  wire _net_2039;
  wire _net_2040;
  wire _net_2041;
  wire _net_2042;
  wire _net_2043;
  wire _net_2044;
  wire _net_2045;
  wire _net_2046;
  wire _net_2047;
  wire _net_2048;
  wire _net_2049;
  wire _net_2050;
  wire _net_2051;
  wire _net_2052;
  wire _net_2053;
  wire _net_2054;
  wire _net_2055;
  wire _net_2056;
  wire _net_2057;
  wire _net_2058;
  wire _net_2059;
  wire _net_2060;
  wire _net_2061;
  wire _net_2062;
  wire _net_2063;
  wire _net_2064;
  wire _net_2065;
  wire _net_2066;
  wire _net_2067;
  wire _net_2068;
  wire _net_2069;
  wire _net_2070;
  wire _net_2071;
  wire _net_2072;
  wire _net_2073;
  wire _net_2074;
  wire _net_2075;
  wire _net_2076;
  wire _net_2077;
  wire _net_2078;
  wire _net_2079;
  wire _net_2080;
  wire _net_2081;
  wire _net_2082;
  wire _net_2083;
  wire _net_2084;
  wire _net_2085;
  wire _net_2086;
  wire _net_2087;
  wire _net_2088;
  wire _net_2089;
  wire _net_2090;
  wire _net_2091;
  wire _net_2092;
  wire _net_2093;
  wire _net_2094;
  wire _net_2095;
  wire _net_2096;
  wire _net_2097;
  wire _net_2098;
  wire _net_2099;
  wire _net_2100;
  wire _net_2101;
  wire _net_2102;
  wire _net_2103;
  wire _net_2104;
  wire _net_2105;
  wire _net_2106;
  wire _net_2107;
  wire _net_2108;
  wire _net_2109;
  wire _net_2110;
  wire _net_2111;
  wire _net_2112;
  wire _net_2113;
  wire _net_2114;
  wire _net_2115;
  wire _net_2116;
  wire _net_2117;
  wire _net_2118;
  wire _net_2119;
  wire _net_2120;
  wire _net_2121;
  wire _net_2122;
  wire _net_2123;
  wire _net_2124;
  wire _net_2125;
  wire _net_2126;
  wire _net_2127;
  wire _net_2128;
  wire _net_2129;
  wire _net_2130;
  wire _net_2131;
  wire _net_2132;
  wire _net_2133;
  wire _net_2134;
  wire _net_2135;
  wire _net_2136;
  wire _net_2137;
  wire _net_2138;
  wire _net_2139;
  wire _net_2140;
  wire _net_2141;
  wire _net_2142;
  wire _net_2143;
  wire _net_2144;
  wire _net_2145;
  wire _net_2146;
  wire _net_2147;
  wire _net_2148;
  wire _net_2149;
  wire _net_2150;
  wire _net_2151;
  wire _net_2152;
  wire _net_2153;
  wire _net_2154;
  wire _net_2155;
  wire _net_2156;
  wire _net_2157;
  wire _net_2158;
  wire _net_2159;
  wire _net_2160;
  wire _net_2161;
  wire _net_2162;
  wire _net_2163;
  wire _net_2164;
  wire _net_2165;
  wire _net_2166;
  wire _net_2167;
  wire _net_2168;
  wire _net_2169;
  wire _net_2170;
  wire _net_2171;
  wire _net_2172;
  wire _net_2173;
  wire _net_2174;
  wire _net_2175;
  wire _net_2176;
  wire _net_2177;
  wire _net_2178;
  wire _net_2179;
  wire _net_2180;
  wire _net_2181;
  wire _net_2182;
  wire _net_2183;
  wire _net_2184;
  wire _net_2185;
  wire _net_2186;
  wire _net_2187;
  wire _net_2188;
  wire _net_2189;
  wire _net_2190;
  wire _net_2191;
  wire _net_2192;
  wire _net_2193;
  wire _net_2194;
  wire _net_2195;
  wire _net_2196;
  wire _net_2197;
  wire _net_2198;
  wire _net_2199;
  wire _net_2200;
  wire _net_2201;
  wire _net_2202;
  wire _net_2203;
  wire _net_2204;
  wire _net_2205;
  wire _net_2206;
  wire _net_2207;
  wire _net_2208;
  wire _net_2209;
  wire _net_2210;
  wire _net_2211;
  wire _net_2212;
  wire _net_2213;
  wire _net_2214;
  wire _net_2215;
  wire _net_2216;
  wire _net_2217;
  wire _net_2218;
  wire _net_2219;
  wire _net_2220;
  wire _net_2221;
  wire _net_2222;
  wire _net_2223;
  wire _net_2224;
  wire _net_2225;
  wire _net_2226;
  wire _net_2227;
  wire _net_2228;
  wire _net_2229;
  wire _net_2230;
  wire _net_2231;
  wire _net_2232;
  wire _net_2233;
  wire _net_2234;
  wire _net_2235;
  wire _net_2236;
  wire _net_2237;
  wire _net_2238;
  wire _net_2239;
  wire _net_2240;
  wire _net_2241;
  wire _net_2242;
  wire _net_2243;
  wire _net_2244;
  wire _net_2245;
  wire _net_2246;
  wire _net_2247;
  wire _net_2248;
  wire _net_2249;
  wire _net_2250;
  wire _net_2251;
  wire _net_2252;
  wire _net_2253;
  wire _net_2254;
  wire _net_2255;
  wire _net_2256;
  wire _net_2257;
  wire _net_2258;
  wire _net_2259;
  wire _net_2260;
  wire _net_2261;
  wire _net_2262;
  wire _net_2263;
  wire _net_2264;
  wire _net_2265;
  wire _net_2266;
  wire _net_2267;
  wire _net_2268;
  wire _net_2269;
  wire _net_2270;
  wire _net_2271;
  wire _net_2272;
  wire _net_2273;
  wire _net_2274;
  wire _net_2275;
  wire _net_2276;
  wire _net_2277;
  wire _net_2278;
  wire _net_2279;
  wire _net_2280;
  wire _net_2281;
  wire _net_2282;
  wire _net_2283;
  wire _net_2284;
  wire _net_2285;
  wire _net_2286;
  wire _net_2287;
  wire _net_2288;
  wire _net_2289;
  wire _net_2290;
  wire _net_2291;
  wire _net_2292;
  wire _net_2293;
  wire _net_2294;
  wire _net_2295;
  wire _net_2296;
  wire _net_2297;
  wire _net_2298;
  wire _net_2299;
  wire _net_2300;
  wire _net_2301;
  wire _net_2302;
  wire _net_2303;
  wire _net_2304;
  wire _net_2305;
  wire _net_2306;
  wire _net_2307;
  wire _net_2308;
  wire _net_2309;
  wire _net_2310;
  wire _net_2311;
  wire _net_2312;
  wire _net_2313;
  wire _net_2314;
  wire _net_2315;
  wire _net_2316;
  wire _net_2317;
  wire _net_2318;
  wire _net_2319;
  wire _net_2320;
  wire _net_2321;
  wire _net_2322;
  wire _net_2323;
  wire _net_2324;
  wire _net_2325;
  wire _net_2326;
  wire _net_2327;
  wire _net_2328;
  wire _net_2329;
  wire _net_2330;
  wire _net_2331;
  wire _net_2332;
  wire _net_2333;
  wire _net_2334;
  wire _net_2335;
  wire _net_2336;
  wire _net_2337;
  wire _net_2338;
  wire _net_2339;
  wire _net_2340;
  wire _net_2341;
  wire _net_2342;
  wire _net_2343;
  wire _net_2344;
  wire _net_2345;
  wire _net_2346;
  wire _net_2347;
  wire _net_2348;
  wire _net_2349;
  wire _net_2350;
  wire _net_2351;
  wire _net_2352;
  wire _net_2353;
  wire _net_2354;
  wire _net_2355;
  wire _net_2356;
  wire _net_2357;
  wire _net_2358;
  wire _net_2359;
  wire _net_2360;
  wire _net_2361;
  wire _net_2362;
  wire _net_2363;
  wire _net_2364;
  wire _net_2365;
  wire _net_2366;
  wire _net_2367;
  wire _net_2368;
  wire _net_2369;
  wire _net_2370;
  wire _net_2371;
  wire _net_2372;
  wire _net_2373;
  wire _net_2374;
  wire _net_2375;
  wire _net_2376;
  wire _net_2377;
  wire _net_2378;
  wire _net_2379;
  wire _net_2380;
  wire _net_2381;
  wire _net_2382;
  wire _net_2383;
  wire _net_2384;
  wire _net_2385;
  wire _net_2386;
  wire _net_2387;
  wire _net_2388;
  wire _net_2389;
  wire _net_2390;
  wire _net_2391;
  wire _net_2392;
  wire _net_2393;
  wire _net_2394;
  wire _net_2395;
  wire _net_2396;
  wire _net_2397;
  wire _net_2398;
  wire _net_2399;
  wire _net_2400;
  wire _net_2401;
  wire _net_2402;
  wire _net_2403;
  wire _net_2404;
  wire _net_2405;
  wire _net_2406;
  wire _net_2407;
  wire _net_2408;
  wire _net_2409;
  wire _net_2410;
  wire _net_2411;
  wire _net_2412;
  wire _net_2413;
  wire _net_2414;
  wire _net_2415;
  wire _net_2416;
  wire _net_2417;
  wire _net_2418;
  wire _net_2419;
  wire _net_2420;
  wire _net_2421;
  wire _net_2422;
  wire _net_2423;
  wire _net_2424;
  wire _net_2425;
  wire _net_2426;
  wire _net_2427;
  wire _net_2428;
  wire _net_2429;
  wire _net_2430;
  wire _net_2431;
  wire _net_2432;
  wire _net_2433;
  wire _net_2434;
  wire _net_2435;
  wire _net_2436;
  wire _net_2437;
  wire _net_2438;
  wire _net_2439;
  wire _net_2440;
  wire _net_2441;
  wire _net_2442;
  wire _net_2443;
  wire _net_2444;
  wire _net_2445;
  wire _net_2446;
  wire _net_2447;
  wire _net_2448;
  wire _net_2449;
  wire _net_2450;
  wire _net_2451;
  wire _net_2452;
  wire _net_2453;
  wire _net_2454;
  wire _net_2455;
  wire _net_2456;
  wire _net_2457;
  wire _net_2458;
  wire _net_2459;
  wire _net_2460;
  wire _net_2461;
  wire _net_2462;
  wire _net_2463;
  wire _net_2464;
  wire _net_2465;
  wire _net_2466;
  wire _net_2467;
  wire _net_2468;
  wire _net_2469;
  wire _net_2470;
  wire _net_2471;
  wire _net_2472;
  wire _net_2473;
  wire _net_2474;
  wire _net_2475;
  wire _net_2476;
  wire _net_2477;
  wire _net_2478;
  wire _net_2479;
  wire _net_2480;
  wire _net_2481;
  wire _net_2482;
  wire _net_2483;
  wire _net_2484;
  wire _net_2485;
  wire _net_2486;
  wire _net_2487;
  wire _net_2488;
  wire _net_2489;
  wire _net_2490;
  wire _net_2491;
  wire _net_2492;
  wire _net_2493;
  wire _net_2494;
  wire _net_2495;
  wire _net_2496;
  wire _net_2497;
  wire _net_2498;
  wire _net_2499;
  wire _net_2500;
  wire _net_2501;
  wire _net_2502;
  wire _net_2503;
  wire _net_2504;
  wire _net_2505;
  wire _net_2506;
  wire _net_2507;
  wire _net_2508;
  wire _net_2509;
  wire _net_2510;
  wire _net_2511;
  wire _net_2512;
  wire _net_2513;
  wire _net_2514;
  wire _net_2515;
  wire _net_2516;
  wire _net_2517;
  wire _net_2518;
  wire _net_2519;
  wire _net_2520;
  wire _net_2521;
  wire _net_2522;
  wire _net_2523;
  wire _net_2524;
  wire _net_2525;
  wire _net_2526;
  wire _net_2527;
  wire _net_2528;
  wire _net_2529;
  wire _net_2530;
  wire _net_2531;
  wire _net_2532;
  wire _net_2533;
  wire _net_2534;
  wire _net_2535;
  wire _net_2536;
  wire _net_2537;
  wire _net_2538;
  wire _net_2539;
  wire _net_2540;
  wire _net_2541;
  wire _net_2542;
  wire _net_2543;
  wire _net_2544;
  reg _reg_2545;
  reg _reg_2546;
  wire _net_2549;
  wire _net_2550;
  wire _net_2551;
  wire _net_2552;
  wire _net_2553;
  wire _net_2554;
  wire _net_2555;
  wire _net_2556;
  wire _net_2557;
  wire _net_2558;
  wire _net_2559;
  wire _net_2560;
  wire _net_2561;
  wire _net_2562;
  wire _net_2563;
  wire _net_2564;
  wire _net_2565;
  wire _net_2566;
  wire _net_2567;
  wire _net_2568;
  wire _net_2569;
  wire _net_2570;
  wire _net_2571;
  wire _net_2572;
  wire _net_2573;
  wire _net_2574;
  wire _net_2575;
  wire _net_2576;
  wire _net_2577;
  wire _net_2578;
  wire _net_2579;
  wire _net_2580;
  wire _net_2581;
  wire _net_2582;
  wire _net_2583;
  wire _net_2584;
  wire _net_2585;
  wire _net_2586;
  wire _net_2587;
  wire _net_2588;
  wire _net_2589;
  wire _net_2590;
  wire _net_2591;
  wire _net_2592;
  wire _net_2593;
  wire _net_2594;
  wire _net_2595;
  wire _net_2596;
  wire _net_2597;
  wire _net_2598;
  wire _net_2599;
  wire _net_2600;
  wire _net_2601;
  wire _net_2602;
  wire _net_2603;
  wire _net_2604;
  wire _net_2605;
  wire _net_2606;
  wire _net_2607;
  wire _net_2608;
  wire _net_2609;
  wire _net_2610;
  wire _net_2611;
  wire _net_2612;
  wire _net_2613;
  wire _net_2614;
  wire _net_2615;
  wire _net_2616;
  wire _net_2617;
  wire _net_2618;
  wire _net_2619;
  wire _net_2620;
  wire _net_2621;
  wire _net_2622;
  wire _net_2623;
  wire _net_2624;
  wire _net_2625;
  wire _net_2626;
  wire _net_2627;
  wire _net_2628;
  wire _net_2629;
  wire _net_2630;
  wire _net_2631;
  wire _net_2632;
  wire _net_2633;
  wire _net_2634;
  wire _net_2635;
  wire _net_2636;
  wire _net_2637;
  wire _net_2638;
  wire _net_2639;
  wire _net_2640;
  wire _net_2641;
  wire _net_2642;
  wire _net_2643;
  wire _net_2644;
  wire _net_2645;
  wire _net_2646;
  wire _net_2647;
  wire _net_2648;
  wire _net_2649;
  wire _net_2650;
  wire _net_2651;
  wire _net_2652;
  wire _net_2653;
  wire _net_2654;
  wire _net_2655;
  wire _net_2656;
  wire _net_2657;
  wire _net_2658;
  wire _net_2659;
  wire _net_2660;
  wire _net_2661;
  wire _net_2662;
  wire _net_2663;
  wire _net_2664;
  wire _net_2665;
  wire _net_2666;
  wire _net_2667;
  wire _net_2668;
  wire _net_2669;
  wire _net_2670;
  wire _net_2671;
  wire _net_2672;
  wire _net_2673;
  wire _net_2674;
  wire _net_2675;
  wire _net_2676;
  wire _net_2677;
  wire _net_2678;
  wire _net_2679;
  wire _net_2680;
  wire _net_2681;
  wire _net_2682;
  wire _net_2683;
  wire _net_2684;
  wire _net_2685;
  wire _net_2686;
  wire _net_2687;
  wire _net_2688;
  wire _net_2689;
  wire _net_2690;
  wire _net_2691;
  wire _net_2692;
  wire _net_2693;
  wire _net_2694;
  wire _net_2695;
  wire _net_2696;
  wire _net_2697;
  wire _net_2698;
  wire _net_2699;
  wire _net_2700;
  wire _net_2701;
  wire _net_2702;
  wire _net_2703;
  wire _net_2704;
  wire _net_2705;
  wire _net_2706;
  wire _net_2707;
  wire _net_2708;
  wire _net_2709;
  wire _net_2710;
  wire _net_2711;
  wire _net_2712;
  wire _net_2713;
  wire _net_2714;
  wire _net_2715;
  wire _net_2716;
  wire _net_2717;
  wire _net_2718;
  wire _net_2719;
  wire _net_2720;
  wire _net_2721;
  wire _net_2722;
  wire _net_2723;
  wire _net_2724;
  wire _net_2725;
  wire _net_2726;
  wire _net_2727;
  wire _net_2728;
  wire _net_2729;
  wire _net_2730;
  wire _net_2731;
  wire _net_2732;
  wire _net_2733;
  wire _net_2734;
  wire _net_2735;
  wire _net_2736;
  wire _net_2737;
  wire _net_2738;
  wire _net_2739;
  wire _net_2740;
  wire _net_2741;
  wire _net_2742;
  wire _net_2743;
  wire _net_2744;
  wire _net_2745;
  wire _net_2746;
  wire _net_2747;
  wire _net_2748;
  wire _net_2749;
  wire _net_2750;
  wire _net_2751;
  wire _net_2752;
  wire _net_2753;
  wire _net_2754;
  wire _net_2755;
  wire _net_2756;
  wire _net_2757;
  wire _net_2758;
  wire _net_2759;
  wire _net_2760;
  wire _net_2761;
  wire _net_2762;
  wire _net_2763;
  wire _net_2764;
  wire _net_2765;
  wire _net_2766;
  wire _net_2767;
  wire _net_2768;
  wire _net_2769;
  wire _net_2770;
  wire _net_2771;
  wire _net_2772;
  wire _net_2773;
  wire _net_2774;
  wire _net_2775;
  wire _net_2776;
  wire _net_2777;
  wire _net_2778;
  wire _net_2779;
  wire _net_2780;
  wire _net_2781;
  wire _net_2782;
  wire _net_2783;
  wire _net_2784;
  wire _net_2785;
  wire _net_2786;
  wire _net_2787;
  wire _net_2788;
  wire _net_2789;
  wire _net_2790;
  wire _net_2791;
  wire _net_2792;
  wire _net_2793;
  wire _net_2794;
  wire _net_2795;
  wire _net_2796;
  wire _net_2797;
  wire _net_2798;
  wire _net_2799;
  wire _net_2800;
  wire _net_2801;
  wire _net_2802;
  wire _net_2803;
  wire _net_2804;
  wire _net_2805;
  wire _net_2806;
  wire _net_2807;
  wire _net_2808;
  wire _net_2809;
  wire _net_2810;
  wire _net_2811;
  wire _net_2812;
  wire _net_2813;
  wire _net_2814;
  wire _net_2815;
  wire _net_2816;
  wire _net_2817;
  wire _net_2818;
  wire _net_2819;
  wire _net_2820;
  wire _net_2821;
  wire _net_2822;
  wire _net_2823;
  wire _net_2824;
  wire _net_2825;
  wire _net_2826;
  wire _net_2827;
  wire _net_2828;
  wire _net_2829;
  wire _net_2830;
  wire _net_2831;
  wire _net_2832;
  wire _net_2833;
  wire _net_2834;
  wire _net_2835;
  wire _net_2836;
  wire _net_2837;
  wire _net_2838;
  wire _net_2839;
  wire _net_2840;
  wire _net_2841;
  wire _net_2842;
  wire _net_2843;
  wire _net_2844;
  wire _net_2845;
  wire _net_2846;
  wire _net_2847;
  wire _net_2848;
  wire _net_2849;
  wire _net_2850;
  wire _net_2851;
  wire _net_2852;
  wire _net_2853;
  wire _net_2854;
  wire _net_2855;
  wire _net_2856;
  wire _net_2857;
  wire _net_2858;
  wire _net_2859;
  wire _net_2860;
  wire _net_2861;
  wire _net_2862;
  wire _net_2863;
  wire _net_2864;
  wire _net_2865;
  wire _net_2866;
  wire _net_2867;
  wire _net_2868;
  wire _net_2869;
  wire _net_2870;
  wire _net_2871;
  wire _net_2872;
  wire _net_2873;
  wire _net_2874;
  wire _net_2875;
  wire _net_2876;
  wire _net_2877;
  wire _net_2878;
  wire _net_2879;
  wire _net_2880;
  wire _net_2881;
  wire _net_2882;
  wire _net_2883;
  wire _net_2884;
  wire _net_2885;
  wire _net_2886;
  wire _net_2887;
  wire _net_2888;
  wire _net_2889;
  wire _net_2890;
  wire _net_2891;
  wire _net_2892;
  wire _net_2893;
  wire _net_2894;
  wire _net_2895;
  wire _net_2896;
  wire _net_2897;
  wire _net_2898;
  wire _net_2899;
  wire _net_2900;
  wire _net_2901;
  wire _net_2902;
  wire _net_2903;
  wire _net_2904;
  wire _net_2905;
  wire _net_2906;
  wire _net_2907;
  wire _net_2908;
  wire _net_2909;
  wire _net_2910;
  wire _net_2911;
  wire _net_2912;
  wire _net_2913;
  wire _net_2914;
  wire _net_2915;
  wire _net_2916;
  wire _net_2917;
  wire _net_2918;
  wire _net_2919;
  wire _net_2920;
  wire _net_2921;
  wire _net_2922;
  wire _net_2923;
  wire _net_2924;
  wire _net_2925;
  wire _net_2926;
  wire _net_2927;
  wire _net_2928;
  wire _net_2929;
  wire _net_2930;
  wire _net_2931;
  wire _net_2932;
  wire _net_2933;
  wire _net_2934;
  wire _net_2935;
  wire _net_2936;
  wire _net_2937;
  wire _net_2938;
  wire _net_2939;
  wire _net_2940;
  wire _net_2941;
  wire _net_2942;
  wire _net_2943;
  wire _net_2944;
  wire _net_2945;
  wire _net_2946;
  wire _net_2947;
  wire _net_2948;
  wire _net_2949;
  wire _net_2950;
  wire _net_2951;
  wire _net_2952;
  wire _net_2953;
  wire _net_2954;
  wire _net_2955;
  wire _net_2956;
  wire _net_2957;
  wire _net_2958;
  wire _net_2959;
  wire _net_2960;
  wire _net_2961;
  wire _net_2962;
  wire _net_2963;
  wire _net_2964;
  wire _net_2965;
  wire _net_2966;
  wire _net_2967;
  wire _net_2968;
  wire _net_2969;
  wire _net_2970;
  wire _net_2971;
  wire _net_2972;
  wire _net_2973;
  wire _net_2974;
  wire _net_2975;
  wire _net_2976;
  wire _net_2977;
  wire _net_2978;
  wire _net_2979;
  wire _net_2980;
  wire _net_2981;
  wire _net_2982;
  wire _net_2983;
  wire _net_2984;
  wire _net_2985;
  wire _net_2986;
  wire _net_2987;
  wire _net_2988;
  wire _net_2989;
  wire _net_2990;
  wire _net_2991;
  wire _net_2992;
  wire _net_2993;
  wire _net_2994;
  wire _net_2995;
  wire _net_2996;
  wire _net_2997;
  wire _net_2998;
  wire _net_2999;
  wire _net_3000;
  wire _net_3001;
  wire _net_3002;
  wire _net_3003;
  wire _net_3004;
  wire _net_3005;
  wire _net_3006;
  wire _net_3007;
  wire _net_3008;
  wire _net_3009;
  wire _net_3010;
  wire _net_3011;
  wire _net_3012;
  wire _net_3013;
  wire _net_3014;
  wire _net_3015;
  wire _net_3016;
  wire _net_3017;
  wire _net_3018;
  wire _net_3019;
  wire _net_3020;
  wire _net_3021;
  wire _net_3022;
  wire _net_3023;
  wire _net_3024;
  wire _net_3025;
  wire _net_3026;
  wire _net_3027;
  wire _net_3028;
  wire _net_3029;
  wire _net_3030;
  wire _net_3031;
  wire _net_3032;
  wire _net_3033;
  wire _net_3034;
  wire _net_3035;
  wire _net_3036;
  wire _net_3037;
  wire _net_3038;
  wire _net_3039;
  wire _net_3040;
  wire _net_3041;
  wire _net_3042;
  wire _net_3043;
  wire _net_3044;
  wire _net_3045;
  wire _net_3046;
  wire _net_3047;
  wire _net_3048;
  wire _net_3049;
  wire _net_3050;
  wire _net_3051;
  wire _net_3052;
  wire _net_3053;
  wire _net_3054;
  wire _net_3055;
  wire _net_3056;
  wire _net_3057;
  wire _net_3058;
  wire _net_3059;
  wire _net_3060;
  wire _net_3061;
  wire _net_3062;
  wire _net_3063;
  wire _net_3064;
  wire _net_3065;
  wire _net_3066;
  wire _net_3067;
  wire _net_3068;
  wire _net_3069;
  wire _net_3070;
  wire _net_3071;
  wire _net_3072;
  wire _net_3073;
  wire _net_3074;
  wire _net_3075;
  wire _net_3076;
  wire _net_3077;
  wire _net_3078;
  wire _net_3079;
  wire _net_3080;
  wire _net_3081;
  wire _net_3082;
  wire _net_3083;
  wire _net_3084;
  wire _net_3085;
  wire _net_3086;
  wire _net_3087;
  wire _net_3088;
  wire _net_3089;
  wire _net_3090;
  wire _net_3091;
  wire _net_3092;
  wire _net_3093;
  wire _net_3094;
  wire _net_3095;
  wire _net_3096;
  wire _net_3097;
  wire _net_3098;
  wire _net_3099;
  wire _net_3100;
  wire _net_3101;
  wire _net_3102;
  wire _net_3103;
  wire _net_3104;
  wire _net_3105;
  wire _net_3106;
  wire _net_3107;
  wire _net_3108;
  wire _net_3109;
  wire _net_3110;
  wire _net_3111;
  wire _net_3112;
  wire _net_3113;
  wire _net_3114;
  wire _net_3115;
  wire _net_3116;
  wire _net_3117;
  wire _net_3118;
  wire _net_3119;
  wire _net_3120;
  wire _net_3121;
  wire _net_3122;
  wire _net_3123;
  wire _net_3124;
  wire _net_3125;
  wire _net_3126;
  wire _net_3127;
  wire _net_3128;
  wire _net_3129;
  wire _net_3130;
  wire _net_3131;
  wire _net_3132;
  wire _net_3133;
  wire _net_3134;
  wire _net_3135;
  wire _net_3136;
  wire _net_3137;
  wire _net_3138;
  wire _net_3139;
  wire _net_3140;
  wire _net_3141;
  wire _net_3142;
  wire _net_3143;
  wire _net_3144;
  wire _net_3145;
  wire _net_3146;
  wire _net_3147;
  wire _net_3148;
  wire _net_3149;
  wire _net_3150;
  wire _net_3151;
  wire _net_3152;
  wire _net_3153;
  wire _net_3154;
  wire _net_3155;
  wire _net_3156;
  wire _net_3157;
  wire _net_3158;
  wire _net_3159;
  wire _net_3160;
  wire _net_3161;
  wire _net_3162;
  wire _net_3163;
  wire _net_3164;
  wire _net_3165;
  wire _net_3166;
  wire _net_3167;
  wire _net_3168;
  wire _net_3169;
  wire _net_3170;
  wire _net_3171;
  wire _net_3172;
  wire _net_3173;
  wire _net_3174;
  wire _net_3175;
  wire _net_3176;
  wire _net_3177;
  wire _net_3178;
  wire _net_3179;
  wire _net_3180;
  wire _net_3181;
  wire _net_3182;
  wire _net_3183;
  wire _net_3184;
  wire _net_3185;
  wire _net_3186;
  wire _net_3187;
  wire _net_3188;
  wire _net_3189;
  wire _net_3190;
  wire _net_3191;
  wire _net_3192;
  wire _net_3193;
  wire _net_3194;
  wire _net_3195;
  wire _net_3196;
  wire _net_3197;
  wire _net_3198;
  wire _net_3199;
  wire _net_3200;
  wire _net_3201;
  wire _net_3202;
  wire _net_3203;
  wire _net_3204;
  wire _net_3205;
  wire _net_3206;
  wire _net_3207;
  wire _net_3208;
  wire _net_3209;
  wire _net_3210;
  wire _net_3211;
  wire _net_3212;
  wire _net_3213;
  wire _net_3214;
  wire _net_3215;
  wire _net_3216;
  wire _net_3217;
  wire _net_3218;
  wire _net_3219;
  wire _net_3220;
  wire _net_3221;
  wire _net_3222;
  wire _net_3223;
  wire _net_3224;
  wire _net_3225;
  wire _net_3226;
  wire _net_3227;
  wire _net_3228;
  wire _net_3229;
  wire _net_3230;
  wire _net_3231;
  wire _net_3232;
  wire _net_3233;
  wire _net_3234;
  wire _net_3235;
  wire _net_3236;
  wire _net_3237;
  wire _net_3238;
  wire _net_3239;
  wire _net_3240;
  wire _net_3241;
  wire _net_3242;
  wire _net_3243;
  wire _net_3244;
  wire _net_3245;
  wire _net_3246;
  wire _net_3247;
  wire _net_3248;
  wire _net_3249;
  wire _net_3250;
  wire _net_3251;
  wire _net_3252;
  wire _net_3253;
  wire _net_3254;
  wire _net_3255;
  wire _net_3256;
  wire _net_3257;
  wire _net_3258;
  wire _net_3259;
  wire _net_3260;
  wire _net_3261;
  wire _net_3262;
  wire _net_3263;
  wire _net_3264;
  wire _net_3265;
  wire _net_3266;
  wire _net_3267;
  wire _net_3268;
  wire _net_3269;
  wire _net_3270;
  wire _net_3271;
  wire _net_3272;
  wire _net_3273;
  wire _net_3274;
  wire _net_3275;
  wire _net_3276;
  wire _net_3277;
  wire _net_3278;
  wire _net_3279;
  wire _net_3280;
  wire _net_3281;
  wire _net_3282;
  wire _net_3283;
  wire _net_3284;
  wire _net_3285;
  wire _net_3286;
  wire _net_3287;
  wire _net_3288;
  wire _net_3289;
  wire _net_3290;
  wire _net_3291;
  wire _net_3292;
  wire _net_3293;
  wire _net_3294;
  wire _net_3295;
  wire _net_3296;
  wire _net_3297;
  wire _net_3298;
  wire _net_3299;
  wire _net_3300;
  wire _net_3301;
  wire _net_3302;
  wire _net_3303;
  wire _net_3304;
  wire _net_3305;
  wire _net_3306;
  wire _net_3307;
  wire _net_3308;
  wire _net_3309;
  wire _net_3310;
  wire _net_3311;
  wire _net_3312;
  wire _net_3313;
  wire _net_3314;
  wire _net_3315;
  wire _net_3316;
  wire _net_3317;
  wire _net_3318;
  wire _net_3319;
  wire _net_3320;
  wire _net_3321;
  wire _net_3322;
  wire _net_3323;
  wire _net_3324;
  wire _net_3325;
  wire _net_3326;
  wire _net_3327;
  wire _net_3328;
  wire _net_3329;
  wire _net_3330;
  wire _net_3331;
  wire _net_3332;
  wire _net_3333;
  wire _net_3334;
  wire _net_3335;
  wire _net_3336;
  wire _net_3337;
  wire _net_3338;
  wire _net_3339;
  wire _net_3340;
  wire _net_3341;
  wire _net_3342;
  wire _net_3343;
  wire _net_3344;
  wire _net_3345;
  wire _net_3346;
  wire _net_3347;
  wire _net_3348;
  wire _net_3349;
  wire _net_3350;
  wire _net_3351;
  wire _net_3352;
  wire _net_3353;
  wire _net_3354;
  wire _net_3355;
  wire _net_3356;
  wire _net_3357;
  wire _net_3358;
  wire _net_3359;
  wire _net_3360;
  wire _net_3361;
  wire _net_3362;
  wire _net_3363;
  wire _net_3364;
  wire _net_3365;
  wire _net_3366;
  wire _net_3367;
  wire _net_3368;
  wire _net_3369;
  wire _net_3370;
  wire _net_3371;
  wire _net_3372;
  wire _net_3373;
  wire _net_3374;
  wire _net_3375;
  wire _net_3376;
  wire _net_3377;
  wire _net_3378;
  wire _net_3379;
  wire _net_3380;
  wire _net_3381;
  wire _net_3382;
  wire _net_3383;
  wire _net_3384;
  wire _net_3385;
  wire _net_3386;
  wire _net_3387;
  wire _net_3388;
  wire _net_3389;
  wire _net_3390;
  wire _net_3391;
  wire _net_3392;
  wire _net_3393;
  wire _net_3394;
  wire _net_3395;
  wire _net_3396;
  wire _net_3398;
subs sub_x (.m_clock(m_clock), .p_reset( p_reset), .subs_exe(_sub_x_subs_exe), .sub_array_out(_sub_x_sub_array_out), .data_in33(_sub_x_data_in33), .data_in35(_sub_x_data_in35), .data_in37(_sub_x_data_in37), .data_in39(_sub_x_data_in39), .data_in41(_sub_x_data_in41), .data_in43(_sub_x_data_in43), .data_in45(_sub_x_data_in45), .data_in47(_sub_x_data_in47), .data_in49(_sub_x_data_in49), .data_in51(_sub_x_data_in51), .data_in53(_sub_x_data_in53), .data_in55(_sub_x_data_in55), .data_in57(_sub_x_data_in57), .data_in59(_sub_x_data_in59), .data_in61(_sub_x_data_in61), .data_in65(_sub_x_data_in65), .data_in67(_sub_x_data_in67), .data_in69(_sub_x_data_in69), .data_in71(_sub_x_data_in71), .data_in73(_sub_x_data_in73), .data_in75(_sub_x_data_in75), .data_in77(_sub_x_data_in77), .data_in79(_sub_x_data_in79), .data_in81(_sub_x_data_in81), .data_in83(_sub_x_data_in83), .data_in85(_sub_x_data_in85), .data_in87(_sub_x_data_in87), .data_in89(_sub_x_data_in89), .data_in91(_sub_x_data_in91), .data_in93(_sub_x_data_in93), .data_in97(_sub_x_data_in97), .data_in99(_sub_x_data_in99), .data_in101(_sub_x_data_in101), .data_in103(_sub_x_data_in103), .data_in105(_sub_x_data_in105), .data_in107(_sub_x_data_in107), .data_in109(_sub_x_data_in109), .data_in111(_sub_x_data_in111), .data_in113(_sub_x_data_in113), .data_in115(_sub_x_data_in115), .data_in117(_sub_x_data_in117), .data_in119(_sub_x_data_in119), .data_in121(_sub_x_data_in121), .data_in123(_sub_x_data_in123), .data_in125(_sub_x_data_in125), .data_in129(_sub_x_data_in129), .data_in131(_sub_x_data_in131), .data_in133(_sub_x_data_in133), .data_in135(_sub_x_data_in135), .data_in137(_sub_x_data_in137), .data_in139(_sub_x_data_in139), .data_in141(_sub_x_data_in141), .data_in143(_sub_x_data_in143), .data_in145(_sub_x_data_in145), .data_in147(_sub_x_data_in147), .data_in149(_sub_x_data_in149), .data_in151(_sub_x_data_in151), .data_in153(_sub_x_data_in153), .data_in155(_sub_x_data_in155), .data_in157(_sub_x_data_in157), .data_in161(_sub_x_data_in161), .data_in163(_sub_x_data_in163), .data_in165(_sub_x_data_in165), .data_in167(_sub_x_data_in167), .data_in169(_sub_x_data_in169), .data_in171(_sub_x_data_in171), .data_in173(_sub_x_data_in173), .data_in175(_sub_x_data_in175), .data_in177(_sub_x_data_in177), .data_in179(_sub_x_data_in179), .data_in181(_sub_x_data_in181), .data_in183(_sub_x_data_in183), .data_in185(_sub_x_data_in185), .data_in187(_sub_x_data_in187), .data_in189(_sub_x_data_in189), .data_in193(_sub_x_data_in193), .data_in195(_sub_x_data_in195), .data_in197(_sub_x_data_in197), .data_in199(_sub_x_data_in199), .data_in201(_sub_x_data_in201), .data_in203(_sub_x_data_in203), .data_in205(_sub_x_data_in205), .data_in207(_sub_x_data_in207), .data_in209(_sub_x_data_in209), .data_in211(_sub_x_data_in211), .data_in213(_sub_x_data_in213), .data_in215(_sub_x_data_in215), .data_in217(_sub_x_data_in217), .data_in219(_sub_x_data_in219), .data_in221(_sub_x_data_in221), .data_in225(_sub_x_data_in225), .data_in227(_sub_x_data_in227), .data_in229(_sub_x_data_in229), .data_in231(_sub_x_data_in231), .data_in233(_sub_x_data_in233), .data_in235(_sub_x_data_in235), .data_in237(_sub_x_data_in237), .data_in239(_sub_x_data_in239), .data_in241(_sub_x_data_in241), .data_in243(_sub_x_data_in243), .data_in245(_sub_x_data_in245), .data_in247(_sub_x_data_in247), .data_in249(_sub_x_data_in249), .data_in251(_sub_x_data_in251), .data_in253(_sub_x_data_in253), .data_in257(_sub_x_data_in257), .data_in259(_sub_x_data_in259), .data_in261(_sub_x_data_in261), .data_in263(_sub_x_data_in263), .data_in265(_sub_x_data_in265), .data_in267(_sub_x_data_in267), .data_in269(_sub_x_data_in269), .data_in271(_sub_x_data_in271), .data_in273(_sub_x_data_in273), .data_in275(_sub_x_data_in275), .data_in277(_sub_x_data_in277), .data_in279(_sub_x_data_in279), .data_in281(_sub_x_data_in281), .data_in283(_sub_x_data_in283), .data_in285(_sub_x_data_in285), .data_in289(_sub_x_data_in289), .data_in291(_sub_x_data_in291), .data_in293(_sub_x_data_in293), .data_in295(_sub_x_data_in295), .data_in297(_sub_x_data_in297), .data_in299(_sub_x_data_in299), .data_in301(_sub_x_data_in301), .data_in303(_sub_x_data_in303), .data_in305(_sub_x_data_in305), .data_in307(_sub_x_data_in307), .data_in309(_sub_x_data_in309), .data_in311(_sub_x_data_in311), .data_in313(_sub_x_data_in313), .data_in315(_sub_x_data_in315), .data_in317(_sub_x_data_in317), .data_in321(_sub_x_data_in321), .data_in323(_sub_x_data_in323), .data_in325(_sub_x_data_in325), .data_in327(_sub_x_data_in327), .data_in329(_sub_x_data_in329), .data_in331(_sub_x_data_in331), .data_in333(_sub_x_data_in333), .data_in335(_sub_x_data_in335), .data_in337(_sub_x_data_in337), .data_in339(_sub_x_data_in339), .data_in341(_sub_x_data_in341), .data_in343(_sub_x_data_in343), .data_in345(_sub_x_data_in345), .data_in347(_sub_x_data_in347), .data_in349(_sub_x_data_in349), .data_in353(_sub_x_data_in353), .data_in355(_sub_x_data_in355), .data_in357(_sub_x_data_in357), .data_in359(_sub_x_data_in359), .data_in361(_sub_x_data_in361), .data_in363(_sub_x_data_in363), .data_in365(_sub_x_data_in365), .data_in367(_sub_x_data_in367), .data_in369(_sub_x_data_in369), .data_in371(_sub_x_data_in371), .data_in373(_sub_x_data_in373), .data_in375(_sub_x_data_in375), .data_in377(_sub_x_data_in377), .data_in379(_sub_x_data_in379), .data_in381(_sub_x_data_in381), .data_in385(_sub_x_data_in385), .data_in387(_sub_x_data_in387), .data_in389(_sub_x_data_in389), .data_in391(_sub_x_data_in391), .data_in393(_sub_x_data_in393), .data_in395(_sub_x_data_in395), .data_in397(_sub_x_data_in397), .data_in399(_sub_x_data_in399), .data_in401(_sub_x_data_in401), .data_in403(_sub_x_data_in403), .data_in405(_sub_x_data_in405), .data_in407(_sub_x_data_in407), .data_in409(_sub_x_data_in409), .data_in411(_sub_x_data_in411), .data_in413(_sub_x_data_in413), .data_in417(_sub_x_data_in417), .data_in419(_sub_x_data_in419), .data_in421(_sub_x_data_in421), .data_in423(_sub_x_data_in423), .data_in425(_sub_x_data_in425), .data_in427(_sub_x_data_in427), .data_in429(_sub_x_data_in429), .data_in431(_sub_x_data_in431), .data_in433(_sub_x_data_in433), .data_in435(_sub_x_data_in435), .data_in437(_sub_x_data_in437), .data_in439(_sub_x_data_in439), .data_in441(_sub_x_data_in441), .data_in443(_sub_x_data_in443), .data_in445(_sub_x_data_in445), .data_in449(_sub_x_data_in449), .data_in451(_sub_x_data_in451), .data_in453(_sub_x_data_in453), .data_in455(_sub_x_data_in455), .data_in457(_sub_x_data_in457), .data_in459(_sub_x_data_in459), .data_in461(_sub_x_data_in461), .data_in463(_sub_x_data_in463), .data_in465(_sub_x_data_in465), .data_in467(_sub_x_data_in467), .data_in469(_sub_x_data_in469), .data_in471(_sub_x_data_in471), .data_in473(_sub_x_data_in473), .data_in475(_sub_x_data_in475), .data_in477(_sub_x_data_in477), .data_in_index33(_sub_x_data_in_index33), .data_in_index35(_sub_x_data_in_index35), .data_in_index37(_sub_x_data_in_index37), .data_in_index39(_sub_x_data_in_index39), .data_in_index41(_sub_x_data_in_index41), .data_in_index43(_sub_x_data_in_index43), .data_in_index45(_sub_x_data_in_index45), .data_in_index47(_sub_x_data_in_index47), .data_in_index49(_sub_x_data_in_index49), .data_in_index51(_sub_x_data_in_index51), .data_in_index53(_sub_x_data_in_index53), .data_in_index55(_sub_x_data_in_index55), .data_in_index57(_sub_x_data_in_index57), .data_in_index59(_sub_x_data_in_index59), .data_in_index61(_sub_x_data_in_index61), .data_in_index65(_sub_x_data_in_index65), .data_in_index67(_sub_x_data_in_index67), .data_in_index69(_sub_x_data_in_index69), .data_in_index71(_sub_x_data_in_index71), .data_in_index73(_sub_x_data_in_index73), .data_in_index75(_sub_x_data_in_index75), .data_in_index77(_sub_x_data_in_index77), .data_in_index79(_sub_x_data_in_index79), .data_in_index81(_sub_x_data_in_index81), .data_in_index83(_sub_x_data_in_index83), .data_in_index85(_sub_x_data_in_index85), .data_in_index87(_sub_x_data_in_index87), .data_in_index89(_sub_x_data_in_index89), .data_in_index91(_sub_x_data_in_index91), .data_in_index93(_sub_x_data_in_index93), .data_in_index97(_sub_x_data_in_index97), .data_in_index99(_sub_x_data_in_index99), .data_in_index101(_sub_x_data_in_index101), .data_in_index103(_sub_x_data_in_index103), .data_in_index105(_sub_x_data_in_index105), .data_in_index107(_sub_x_data_in_index107), .data_in_index109(_sub_x_data_in_index109), .data_in_index111(_sub_x_data_in_index111), .data_in_index113(_sub_x_data_in_index113), .data_in_index115(_sub_x_data_in_index115), .data_in_index117(_sub_x_data_in_index117), .data_in_index119(_sub_x_data_in_index119), .data_in_index121(_sub_x_data_in_index121), .data_in_index123(_sub_x_data_in_index123), .data_in_index125(_sub_x_data_in_index125), .data_in_index129(_sub_x_data_in_index129), .data_in_index131(_sub_x_data_in_index131), .data_in_index133(_sub_x_data_in_index133), .data_in_index135(_sub_x_data_in_index135), .data_in_index137(_sub_x_data_in_index137), .data_in_index139(_sub_x_data_in_index139), .data_in_index141(_sub_x_data_in_index141), .data_in_index143(_sub_x_data_in_index143), .data_in_index145(_sub_x_data_in_index145), .data_in_index147(_sub_x_data_in_index147), .data_in_index149(_sub_x_data_in_index149), .data_in_index151(_sub_x_data_in_index151), .data_in_index153(_sub_x_data_in_index153), .data_in_index155(_sub_x_data_in_index155), .data_in_index157(_sub_x_data_in_index157), .data_in_index161(_sub_x_data_in_index161), .data_in_index163(_sub_x_data_in_index163), .data_in_index165(_sub_x_data_in_index165), .data_in_index167(_sub_x_data_in_index167), .data_in_index169(_sub_x_data_in_index169), .data_in_index171(_sub_x_data_in_index171), .data_in_index173(_sub_x_data_in_index173), .data_in_index175(_sub_x_data_in_index175), .data_in_index177(_sub_x_data_in_index177), .data_in_index179(_sub_x_data_in_index179), .data_in_index181(_sub_x_data_in_index181), .data_in_index183(_sub_x_data_in_index183), .data_in_index185(_sub_x_data_in_index185), .data_in_index187(_sub_x_data_in_index187), .data_in_index189(_sub_x_data_in_index189), .data_in_index193(_sub_x_data_in_index193), .data_in_index195(_sub_x_data_in_index195), .data_in_index197(_sub_x_data_in_index197), .data_in_index199(_sub_x_data_in_index199), .data_in_index201(_sub_x_data_in_index201), .data_in_index203(_sub_x_data_in_index203), .data_in_index205(_sub_x_data_in_index205), .data_in_index207(_sub_x_data_in_index207), .data_in_index209(_sub_x_data_in_index209), .data_in_index211(_sub_x_data_in_index211), .data_in_index213(_sub_x_data_in_index213), .data_in_index215(_sub_x_data_in_index215), .data_in_index217(_sub_x_data_in_index217), .data_in_index219(_sub_x_data_in_index219), .data_in_index221(_sub_x_data_in_index221), .data_in_index225(_sub_x_data_in_index225), .data_in_index227(_sub_x_data_in_index227), .data_in_index229(_sub_x_data_in_index229), .data_in_index231(_sub_x_data_in_index231), .data_in_index233(_sub_x_data_in_index233), .data_in_index235(_sub_x_data_in_index235), .data_in_index237(_sub_x_data_in_index237), .data_in_index239(_sub_x_data_in_index239), .data_in_index241(_sub_x_data_in_index241), .data_in_index243(_sub_x_data_in_index243), .data_in_index245(_sub_x_data_in_index245), .data_in_index247(_sub_x_data_in_index247), .data_in_index249(_sub_x_data_in_index249), .data_in_index251(_sub_x_data_in_index251), .data_in_index253(_sub_x_data_in_index253), .data_in_index257(_sub_x_data_in_index257), .data_in_index259(_sub_x_data_in_index259), .data_in_index261(_sub_x_data_in_index261), .data_in_index263(_sub_x_data_in_index263), .data_in_index265(_sub_x_data_in_index265), .data_in_index267(_sub_x_data_in_index267), .data_in_index269(_sub_x_data_in_index269), .data_in_index271(_sub_x_data_in_index271), .data_in_index273(_sub_x_data_in_index273), .data_in_index275(_sub_x_data_in_index275), .data_in_index277(_sub_x_data_in_index277), .data_in_index279(_sub_x_data_in_index279), .data_in_index281(_sub_x_data_in_index281), .data_in_index283(_sub_x_data_in_index283), .data_in_index285(_sub_x_data_in_index285), .data_in_index289(_sub_x_data_in_index289), .data_in_index291(_sub_x_data_in_index291), .data_in_index293(_sub_x_data_in_index293), .data_in_index295(_sub_x_data_in_index295), .data_in_index297(_sub_x_data_in_index297), .data_in_index299(_sub_x_data_in_index299), .data_in_index301(_sub_x_data_in_index301), .data_in_index303(_sub_x_data_in_index303), .data_in_index305(_sub_x_data_in_index305), .data_in_index307(_sub_x_data_in_index307), .data_in_index309(_sub_x_data_in_index309), .data_in_index311(_sub_x_data_in_index311), .data_in_index313(_sub_x_data_in_index313), .data_in_index315(_sub_x_data_in_index315), .data_in_index317(_sub_x_data_in_index317), .data_in_index321(_sub_x_data_in_index321), .data_in_index323(_sub_x_data_in_index323), .data_in_index325(_sub_x_data_in_index325), .data_in_index327(_sub_x_data_in_index327), .data_in_index329(_sub_x_data_in_index329), .data_in_index331(_sub_x_data_in_index331), .data_in_index333(_sub_x_data_in_index333), .data_in_index335(_sub_x_data_in_index335), .data_in_index337(_sub_x_data_in_index337), .data_in_index339(_sub_x_data_in_index339), .data_in_index341(_sub_x_data_in_index341), .data_in_index343(_sub_x_data_in_index343), .data_in_index345(_sub_x_data_in_index345), .data_in_index347(_sub_x_data_in_index347), .data_in_index349(_sub_x_data_in_index349), .data_in_index353(_sub_x_data_in_index353), .data_in_index355(_sub_x_data_in_index355), .data_in_index357(_sub_x_data_in_index357), .data_in_index359(_sub_x_data_in_index359), .data_in_index361(_sub_x_data_in_index361), .data_in_index363(_sub_x_data_in_index363), .data_in_index365(_sub_x_data_in_index365), .data_in_index367(_sub_x_data_in_index367), .data_in_index369(_sub_x_data_in_index369), .data_in_index371(_sub_x_data_in_index371), .data_in_index373(_sub_x_data_in_index373), .data_in_index375(_sub_x_data_in_index375), .data_in_index377(_sub_x_data_in_index377), .data_in_index379(_sub_x_data_in_index379), .data_in_index381(_sub_x_data_in_index381), .data_in_index385(_sub_x_data_in_index385), .data_in_index387(_sub_x_data_in_index387), .data_in_index389(_sub_x_data_in_index389), .data_in_index391(_sub_x_data_in_index391), .data_in_index393(_sub_x_data_in_index393), .data_in_index395(_sub_x_data_in_index395), .data_in_index397(_sub_x_data_in_index397), .data_in_index399(_sub_x_data_in_index399), .data_in_index401(_sub_x_data_in_index401), .data_in_index403(_sub_x_data_in_index403), .data_in_index405(_sub_x_data_in_index405), .data_in_index407(_sub_x_data_in_index407), .data_in_index409(_sub_x_data_in_index409), .data_in_index411(_sub_x_data_in_index411), .data_in_index413(_sub_x_data_in_index413), .data_in_index417(_sub_x_data_in_index417), .data_in_index419(_sub_x_data_in_index419), .data_in_index421(_sub_x_data_in_index421), .data_in_index423(_sub_x_data_in_index423), .data_in_index425(_sub_x_data_in_index425), .data_in_index427(_sub_x_data_in_index427), .data_in_index429(_sub_x_data_in_index429), .data_in_index431(_sub_x_data_in_index431), .data_in_index433(_sub_x_data_in_index433), .data_in_index435(_sub_x_data_in_index435), .data_in_index437(_sub_x_data_in_index437), .data_in_index439(_sub_x_data_in_index439), .data_in_index441(_sub_x_data_in_index441), .data_in_index443(_sub_x_data_in_index443), .data_in_index445(_sub_x_data_in_index445), .data_in_index449(_sub_x_data_in_index449), .data_in_index451(_sub_x_data_in_index451), .data_in_index453(_sub_x_data_in_index453), .data_in_index455(_sub_x_data_in_index455), .data_in_index457(_sub_x_data_in_index457), .data_in_index459(_sub_x_data_in_index459), .data_in_index461(_sub_x_data_in_index461), .data_in_index463(_sub_x_data_in_index463), .data_in_index465(_sub_x_data_in_index465), .data_in_index467(_sub_x_data_in_index467), .data_in_index469(_sub_x_data_in_index469), .data_in_index471(_sub_x_data_in_index471), .data_in_index473(_sub_x_data_in_index473), .data_in_index475(_sub_x_data_in_index475), .data_in_index477(_sub_x_data_in_index477));
add_all add_all_x (.m_clock(m_clock), .p_reset( p_reset), .out_data(_add_all_x_out_data), .out_do(_add_all_x_out_do), .in_do(_add_all_x_in_do), .dig_t0(_add_all_x_dig_t0), .dig_t1(_add_all_x_dig_t1), .dig_t2(_add_all_x_dig_t2), .dig_t3(_add_all_x_dig_t3), .dig_t4(_add_all_x_dig_t4), .dig_t5(_add_all_x_dig_t5), .dig_t6(_add_all_x_dig_t6), .dig_t7(_add_all_x_dig_t7), .dig_t8(_add_all_x_dig_t8), .dig_t9(_add_all_x_dig_t9), .dig_t10(_add_all_x_dig_t10), .dig_t11(_add_all_x_dig_t11), .dig_t12(_add_all_x_dig_t12), .dig_t13(_add_all_x_dig_t13), .dig_t14(_add_all_x_dig_t14), .dig_t15(_add_all_x_dig_t15), .dig_t16(_add_all_x_dig_t16), .dig_t17(_add_all_x_dig_t17), .dig_t18(_add_all_x_dig_t18), .dig_t19(_add_all_x_dig_t19), .dig_t20(_add_all_x_dig_t20), .dig_t21(_add_all_x_dig_t21), .dig_t22(_add_all_x_dig_t22), .dig_t23(_add_all_x_dig_t23), .dig_t24(_add_all_x_dig_t24), .dig_t25(_add_all_x_dig_t25), .dig_t26(_add_all_x_dig_t26), .dig_t27(_add_all_x_dig_t27), .dig_t28(_add_all_x_dig_t28), .dig_t29(_add_all_x_dig_t29), .dig_t30(_add_all_x_dig_t30), .dig_t31(_add_all_x_dig_t31), .dig_t32(_add_all_x_dig_t32), .dig_t33(_add_all_x_dig_t33), .dig_t34(_add_all_x_dig_t34), .dig_t35(_add_all_x_dig_t35), .dig_t36(_add_all_x_dig_t36), .dig_t37(_add_all_x_dig_t37), .dig_t38(_add_all_x_dig_t38), .dig_t39(_add_all_x_dig_t39), .dig_t40(_add_all_x_dig_t40), .dig_t41(_add_all_x_dig_t41), .dig_t42(_add_all_x_dig_t42), .dig_t43(_add_all_x_dig_t43), .dig_t44(_add_all_x_dig_t44), .dig_t45(_add_all_x_dig_t45), .dig_t46(_add_all_x_dig_t46), .dig_t47(_add_all_x_dig_t47), .dig_t48(_add_all_x_dig_t48), .dig_t49(_add_all_x_dig_t49), .dig_t50(_add_all_x_dig_t50), .dig_t51(_add_all_x_dig_t51), .dig_t52(_add_all_x_dig_t52), .dig_t53(_add_all_x_dig_t53), .dig_t54(_add_all_x_dig_t54), .dig_t55(_add_all_x_dig_t55), .dig_t56(_add_all_x_dig_t56), .dig_t57(_add_all_x_dig_t57), .dig_t58(_add_all_x_dig_t58), .dig_t59(_add_all_x_dig_t59), .dig_t60(_add_all_x_dig_t60), .dig_t61(_add_all_x_dig_t61), .dig_t62(_add_all_x_dig_t62), .dig_t63(_add_all_x_dig_t63), .dig_t64(_add_all_x_dig_t64), .dig_t65(_add_all_x_dig_t65), .dig_t66(_add_all_x_dig_t66), .dig_t67(_add_all_x_dig_t67), .dig_t68(_add_all_x_dig_t68), .dig_t69(_add_all_x_dig_t69), .dig_t70(_add_all_x_dig_t70), .dig_t71(_add_all_x_dig_t71), .dig_t72(_add_all_x_dig_t72), .dig_t73(_add_all_x_dig_t73), .dig_t74(_add_all_x_dig_t74), .dig_t75(_add_all_x_dig_t75), .dig_t76(_add_all_x_dig_t76), .dig_t77(_add_all_x_dig_t77), .dig_t78(_add_all_x_dig_t78), .dig_t79(_add_all_x_dig_t79), .dig_t80(_add_all_x_dig_t80), .dig_t81(_add_all_x_dig_t81), .dig_t82(_add_all_x_dig_t82), .dig_t83(_add_all_x_dig_t83), .dig_t84(_add_all_x_dig_t84), .dig_t85(_add_all_x_dig_t85), .dig_t86(_add_all_x_dig_t86), .dig_t87(_add_all_x_dig_t87), .dig_t88(_add_all_x_dig_t88), .dig_t89(_add_all_x_dig_t89), .dig_t90(_add_all_x_dig_t90), .dig_t91(_add_all_x_dig_t91), .dig_t92(_add_all_x_dig_t92), .dig_t93(_add_all_x_dig_t93), .dig_t94(_add_all_x_dig_t94), .dig_t95(_add_all_x_dig_t95), .dig_t96(_add_all_x_dig_t96), .dig_t97(_add_all_x_dig_t97), .dig_t98(_add_all_x_dig_t98), .dig_t99(_add_all_x_dig_t99), .dig_t100(_add_all_x_dig_t100), .dig_t101(_add_all_x_dig_t101), .dig_t102(_add_all_x_dig_t102), .dig_t103(_add_all_x_dig_t103), .dig_t104(_add_all_x_dig_t104), .dig_t105(_add_all_x_dig_t105), .dig_t106(_add_all_x_dig_t106), .dig_t107(_add_all_x_dig_t107), .dig_t108(_add_all_x_dig_t108), .dig_t109(_add_all_x_dig_t109), .dig_t110(_add_all_x_dig_t110), .dig_t111(_add_all_x_dig_t111), .dig_t112(_add_all_x_dig_t112), .dig_t113(_add_all_x_dig_t113), .dig_t114(_add_all_x_dig_t114), .dig_t115(_add_all_x_dig_t115), .dig_t116(_add_all_x_dig_t116), .dig_t117(_add_all_x_dig_t117), .dig_t118(_add_all_x_dig_t118), .dig_t119(_add_all_x_dig_t119), .dig_t120(_add_all_x_dig_t120), .dig_t121(_add_all_x_dig_t121), .dig_t122(_add_all_x_dig_t122), .dig_t123(_add_all_x_dig_t123), .dig_t124(_add_all_x_dig_t124), .dig_t125(_add_all_x_dig_t125), .dig_t126(_add_all_x_dig_t126), .dig_t127(_add_all_x_dig_t127), .dig_t128(_add_all_x_dig_t128), .dig_t129(_add_all_x_dig_t129), .dig_t130(_add_all_x_dig_t130), .dig_t131(_add_all_x_dig_t131), .dig_t132(_add_all_x_dig_t132), .dig_t133(_add_all_x_dig_t133), .dig_t134(_add_all_x_dig_t134), .dig_t135(_add_all_x_dig_t135), .dig_t136(_add_all_x_dig_t136), .dig_t137(_add_all_x_dig_t137), .dig_t138(_add_all_x_dig_t138), .dig_t139(_add_all_x_dig_t139), .dig_t140(_add_all_x_dig_t140), .dig_t141(_add_all_x_dig_t141), .dig_t142(_add_all_x_dig_t142), .dig_t143(_add_all_x_dig_t143), .dig_t144(_add_all_x_dig_t144), .dig_t145(_add_all_x_dig_t145), .dig_t146(_add_all_x_dig_t146), .dig_t147(_add_all_x_dig_t147), .dig_t148(_add_all_x_dig_t148), .dig_t149(_add_all_x_dig_t149), .dig_t150(_add_all_x_dig_t150), .dig_t151(_add_all_x_dig_t151), .dig_t152(_add_all_x_dig_t152), .dig_t153(_add_all_x_dig_t153), .dig_t154(_add_all_x_dig_t154), .dig_t155(_add_all_x_dig_t155), .dig_t156(_add_all_x_dig_t156), .dig_t157(_add_all_x_dig_t157), .dig_t158(_add_all_x_dig_t158), .dig_t159(_add_all_x_dig_t159), .dig_t160(_add_all_x_dig_t160), .dig_t161(_add_all_x_dig_t161), .dig_t162(_add_all_x_dig_t162), .dig_t163(_add_all_x_dig_t163), .dig_t164(_add_all_x_dig_t164), .dig_t165(_add_all_x_dig_t165), .dig_t166(_add_all_x_dig_t166), .dig_t167(_add_all_x_dig_t167), .dig_t168(_add_all_x_dig_t168), .dig_t169(_add_all_x_dig_t169), .dig_t170(_add_all_x_dig_t170), .dig_t171(_add_all_x_dig_t171), .dig_t172(_add_all_x_dig_t172), .dig_t173(_add_all_x_dig_t173), .dig_t174(_add_all_x_dig_t174), .dig_t175(_add_all_x_dig_t175), .dig_t176(_add_all_x_dig_t176), .dig_t177(_add_all_x_dig_t177), .dig_t178(_add_all_x_dig_t178), .dig_t179(_add_all_x_dig_t179), .dig_t180(_add_all_x_dig_t180), .dig_t181(_add_all_x_dig_t181), .dig_t182(_add_all_x_dig_t182), .dig_t183(_add_all_x_dig_t183), .dig_t184(_add_all_x_dig_t184), .dig_t185(_add_all_x_dig_t185), .dig_t186(_add_all_x_dig_t186), .dig_t187(_add_all_x_dig_t187), .dig_t188(_add_all_x_dig_t188), .dig_t189(_add_all_x_dig_t189), .dig_t190(_add_all_x_dig_t190), .dig_t191(_add_all_x_dig_t191), .dig_t192(_add_all_x_dig_t192), .dig_t193(_add_all_x_dig_t193), .dig_t194(_add_all_x_dig_t194), .dig_t195(_add_all_x_dig_t195), .dig_t196(_add_all_x_dig_t196), .dig_t197(_add_all_x_dig_t197), .dig_t198(_add_all_x_dig_t198), .dig_t199(_add_all_x_dig_t199), .dig_t200(_add_all_x_dig_t200), .dig_t201(_add_all_x_dig_t201), .dig_t202(_add_all_x_dig_t202), .dig_t203(_add_all_x_dig_t203), .dig_t204(_add_all_x_dig_t204), .dig_t205(_add_all_x_dig_t205), .dig_t206(_add_all_x_dig_t206), .dig_t207(_add_all_x_dig_t207), .dig_t208(_add_all_x_dig_t208), .dig_t209(_add_all_x_dig_t209), .sg_out33(_add_all_x_sg_out33), .sg_out34(_add_all_x_sg_out34), .sg_out35(_add_all_x_sg_out35), .sg_out36(_add_all_x_sg_out36), .sg_out37(_add_all_x_sg_out37), .sg_out38(_add_all_x_sg_out38), .sg_out39(_add_all_x_sg_out39), .sg_out40(_add_all_x_sg_out40), .sg_out41(_add_all_x_sg_out41), .sg_out42(_add_all_x_sg_out42), .sg_out43(_add_all_x_sg_out43), .sg_out44(_add_all_x_sg_out44), .sg_out45(_add_all_x_sg_out45), .sg_out46(_add_all_x_sg_out46), .sg_out47(_add_all_x_sg_out47), .sg_out48(_add_all_x_sg_out48), .sg_out49(_add_all_x_sg_out49), .sg_out50(_add_all_x_sg_out50), .sg_out51(_add_all_x_sg_out51), .sg_out52(_add_all_x_sg_out52), .sg_out53(_add_all_x_sg_out53), .sg_out54(_add_all_x_sg_out54), .sg_out55(_add_all_x_sg_out55), .sg_out56(_add_all_x_sg_out56), .sg_out57(_add_all_x_sg_out57), .sg_out58(_add_all_x_sg_out58), .sg_out59(_add_all_x_sg_out59), .sg_out60(_add_all_x_sg_out60), .sg_out61(_add_all_x_sg_out61), .sg_out62(_add_all_x_sg_out62), .sg_out65(_add_all_x_sg_out65), .sg_out66(_add_all_x_sg_out66), .sg_out67(_add_all_x_sg_out67), .sg_out68(_add_all_x_sg_out68), .sg_out69(_add_all_x_sg_out69), .sg_out70(_add_all_x_sg_out70), .sg_out71(_add_all_x_sg_out71), .sg_out72(_add_all_x_sg_out72), .sg_out73(_add_all_x_sg_out73), .sg_out74(_add_all_x_sg_out74), .sg_out75(_add_all_x_sg_out75), .sg_out76(_add_all_x_sg_out76), .sg_out77(_add_all_x_sg_out77), .sg_out78(_add_all_x_sg_out78), .sg_out79(_add_all_x_sg_out79), .sg_out80(_add_all_x_sg_out80), .sg_out81(_add_all_x_sg_out81), .sg_out82(_add_all_x_sg_out82), .sg_out83(_add_all_x_sg_out83), .sg_out84(_add_all_x_sg_out84), .sg_out85(_add_all_x_sg_out85), .sg_out86(_add_all_x_sg_out86), .sg_out87(_add_all_x_sg_out87), .sg_out88(_add_all_x_sg_out88), .sg_out89(_add_all_x_sg_out89), .sg_out90(_add_all_x_sg_out90), .sg_out91(_add_all_x_sg_out91), .sg_out92(_add_all_x_sg_out92), .sg_out93(_add_all_x_sg_out93), .sg_out94(_add_all_x_sg_out94), .sg_out97(_add_all_x_sg_out97), .sg_out98(_add_all_x_sg_out98), .sg_out99(_add_all_x_sg_out99), .sg_out100(_add_all_x_sg_out100), .sg_out101(_add_all_x_sg_out101), .sg_out102(_add_all_x_sg_out102), .sg_out103(_add_all_x_sg_out103), .sg_out104(_add_all_x_sg_out104), .sg_out105(_add_all_x_sg_out105), .sg_out106(_add_all_x_sg_out106), .sg_out107(_add_all_x_sg_out107), .sg_out108(_add_all_x_sg_out108), .sg_out109(_add_all_x_sg_out109), .sg_out110(_add_all_x_sg_out110), .sg_out111(_add_all_x_sg_out111), .sg_out112(_add_all_x_sg_out112), .sg_out113(_add_all_x_sg_out113), .sg_out114(_add_all_x_sg_out114), .sg_out115(_add_all_x_sg_out115), .sg_out116(_add_all_x_sg_out116), .sg_out117(_add_all_x_sg_out117), .sg_out118(_add_all_x_sg_out118), .sg_out119(_add_all_x_sg_out119), .sg_out120(_add_all_x_sg_out120), .sg_out121(_add_all_x_sg_out121), .sg_out122(_add_all_x_sg_out122), .sg_out123(_add_all_x_sg_out123), .sg_out124(_add_all_x_sg_out124), .sg_out125(_add_all_x_sg_out125), .sg_out126(_add_all_x_sg_out126), .sg_out129(_add_all_x_sg_out129), .sg_out130(_add_all_x_sg_out130), .sg_out131(_add_all_x_sg_out131), .sg_out132(_add_all_x_sg_out132), .sg_out133(_add_all_x_sg_out133), .sg_out134(_add_all_x_sg_out134), .sg_out135(_add_all_x_sg_out135), .sg_out136(_add_all_x_sg_out136), .sg_out137(_add_all_x_sg_out137), .sg_out138(_add_all_x_sg_out138), .sg_out139(_add_all_x_sg_out139), .sg_out140(_add_all_x_sg_out140), .sg_out141(_add_all_x_sg_out141), .sg_out142(_add_all_x_sg_out142), .sg_out143(_add_all_x_sg_out143), .sg_out144(_add_all_x_sg_out144), .sg_out145(_add_all_x_sg_out145), .sg_out146(_add_all_x_sg_out146), .sg_out147(_add_all_x_sg_out147), .sg_out148(_add_all_x_sg_out148), .sg_out149(_add_all_x_sg_out149), .sg_out150(_add_all_x_sg_out150), .sg_out151(_add_all_x_sg_out151), .sg_out152(_add_all_x_sg_out152), .sg_out153(_add_all_x_sg_out153), .sg_out154(_add_all_x_sg_out154), .sg_out155(_add_all_x_sg_out155), .sg_out156(_add_all_x_sg_out156), .sg_out157(_add_all_x_sg_out157), .sg_out158(_add_all_x_sg_out158), .sg_out161(_add_all_x_sg_out161), .sg_out162(_add_all_x_sg_out162), .sg_out163(_add_all_x_sg_out163), .sg_out164(_add_all_x_sg_out164), .sg_out165(_add_all_x_sg_out165), .sg_out166(_add_all_x_sg_out166), .sg_out167(_add_all_x_sg_out167), .sg_out168(_add_all_x_sg_out168), .sg_out169(_add_all_x_sg_out169), .sg_out170(_add_all_x_sg_out170), .sg_out171(_add_all_x_sg_out171), .sg_out172(_add_all_x_sg_out172), .sg_out173(_add_all_x_sg_out173), .sg_out174(_add_all_x_sg_out174), .sg_out175(_add_all_x_sg_out175), .sg_out176(_add_all_x_sg_out176), .sg_out177(_add_all_x_sg_out177), .sg_out178(_add_all_x_sg_out178), .sg_out179(_add_all_x_sg_out179), .sg_out180(_add_all_x_sg_out180), .sg_out181(_add_all_x_sg_out181), .sg_out182(_add_all_x_sg_out182), .sg_out183(_add_all_x_sg_out183), .sg_out184(_add_all_x_sg_out184), .sg_out185(_add_all_x_sg_out185), .sg_out186(_add_all_x_sg_out186), .sg_out187(_add_all_x_sg_out187), .sg_out188(_add_all_x_sg_out188), .sg_out189(_add_all_x_sg_out189), .sg_out190(_add_all_x_sg_out190), .sg_out193(_add_all_x_sg_out193), .sg_out194(_add_all_x_sg_out194), .sg_out195(_add_all_x_sg_out195), .sg_out196(_add_all_x_sg_out196), .sg_out197(_add_all_x_sg_out197), .sg_out198(_add_all_x_sg_out198), .sg_out199(_add_all_x_sg_out199), .sg_out200(_add_all_x_sg_out200), .sg_out201(_add_all_x_sg_out201), .sg_out202(_add_all_x_sg_out202), .sg_out203(_add_all_x_sg_out203), .sg_out204(_add_all_x_sg_out204), .sg_out205(_add_all_x_sg_out205), .sg_out206(_add_all_x_sg_out206), .sg_out207(_add_all_x_sg_out207), .sg_out208(_add_all_x_sg_out208), .sg_out209(_add_all_x_sg_out209), .sg_out210(_add_all_x_sg_out210), .sg_out211(_add_all_x_sg_out211), .sg_out212(_add_all_x_sg_out212), .sg_out213(_add_all_x_sg_out213), .sg_out214(_add_all_x_sg_out214), .sg_out215(_add_all_x_sg_out215), .sg_out216(_add_all_x_sg_out216), .sg_out217(_add_all_x_sg_out217), .sg_out218(_add_all_x_sg_out218), .sg_out219(_add_all_x_sg_out219), .sg_out220(_add_all_x_sg_out220), .sg_out221(_add_all_x_sg_out221), .sg_out222(_add_all_x_sg_out222), .sg_out225(_add_all_x_sg_out225), .sg_out226(_add_all_x_sg_out226), .sg_out227(_add_all_x_sg_out227), .sg_out228(_add_all_x_sg_out228), .sg_out229(_add_all_x_sg_out229), .sg_out230(_add_all_x_sg_out230), .sg_out231(_add_all_x_sg_out231), .sg_out232(_add_all_x_sg_out232), .sg_out233(_add_all_x_sg_out233), .sg_out234(_add_all_x_sg_out234), .sg_out235(_add_all_x_sg_out235), .sg_out236(_add_all_x_sg_out236), .sg_out237(_add_all_x_sg_out237), .sg_out238(_add_all_x_sg_out238), .sg_out239(_add_all_x_sg_out239), .sg_out240(_add_all_x_sg_out240), .sg_out241(_add_all_x_sg_out241), .sg_out242(_add_all_x_sg_out242), .sg_out243(_add_all_x_sg_out243), .sg_out244(_add_all_x_sg_out244), .sg_out245(_add_all_x_sg_out245), .sg_out246(_add_all_x_sg_out246), .sg_out247(_add_all_x_sg_out247), .sg_out248(_add_all_x_sg_out248), .sg_out249(_add_all_x_sg_out249), .sg_out250(_add_all_x_sg_out250), .sg_out251(_add_all_x_sg_out251), .sg_out252(_add_all_x_sg_out252), .sg_out253(_add_all_x_sg_out253), .sg_out254(_add_all_x_sg_out254), .sg_out257(_add_all_x_sg_out257), .sg_out258(_add_all_x_sg_out258), .sg_out259(_add_all_x_sg_out259), .sg_out260(_add_all_x_sg_out260), .sg_out261(_add_all_x_sg_out261), .sg_out262(_add_all_x_sg_out262), .sg_out263(_add_all_x_sg_out263), .sg_out264(_add_all_x_sg_out264), .sg_out265(_add_all_x_sg_out265), .sg_out266(_add_all_x_sg_out266), .sg_out267(_add_all_x_sg_out267), .sg_out268(_add_all_x_sg_out268), .sg_out269(_add_all_x_sg_out269), .sg_out270(_add_all_x_sg_out270), .sg_out271(_add_all_x_sg_out271), .sg_out272(_add_all_x_sg_out272), .sg_out273(_add_all_x_sg_out273), .sg_out274(_add_all_x_sg_out274), .sg_out275(_add_all_x_sg_out275), .sg_out276(_add_all_x_sg_out276), .sg_out277(_add_all_x_sg_out277), .sg_out278(_add_all_x_sg_out278), .sg_out279(_add_all_x_sg_out279), .sg_out280(_add_all_x_sg_out280), .sg_out281(_add_all_x_sg_out281), .sg_out282(_add_all_x_sg_out282), .sg_out283(_add_all_x_sg_out283), .sg_out284(_add_all_x_sg_out284), .sg_out285(_add_all_x_sg_out285), .sg_out286(_add_all_x_sg_out286), .sg_out289(_add_all_x_sg_out289), .sg_out290(_add_all_x_sg_out290), .sg_out291(_add_all_x_sg_out291), .sg_out292(_add_all_x_sg_out292), .sg_out293(_add_all_x_sg_out293), .sg_out294(_add_all_x_sg_out294), .sg_out295(_add_all_x_sg_out295), .sg_out296(_add_all_x_sg_out296), .sg_out297(_add_all_x_sg_out297), .sg_out298(_add_all_x_sg_out298), .sg_out299(_add_all_x_sg_out299), .sg_out300(_add_all_x_sg_out300), .sg_out301(_add_all_x_sg_out301), .sg_out302(_add_all_x_sg_out302), .sg_out303(_add_all_x_sg_out303), .sg_out304(_add_all_x_sg_out304), .sg_out305(_add_all_x_sg_out305), .sg_out306(_add_all_x_sg_out306), .sg_out307(_add_all_x_sg_out307), .sg_out308(_add_all_x_sg_out308), .sg_out309(_add_all_x_sg_out309), .sg_out310(_add_all_x_sg_out310), .sg_out311(_add_all_x_sg_out311), .sg_out312(_add_all_x_sg_out312), .sg_out313(_add_all_x_sg_out313), .sg_out314(_add_all_x_sg_out314), .sg_out315(_add_all_x_sg_out315), .sg_out316(_add_all_x_sg_out316), .sg_out317(_add_all_x_sg_out317), .sg_out318(_add_all_x_sg_out318), .sg_out321(_add_all_x_sg_out321), .sg_out322(_add_all_x_sg_out322), .sg_out323(_add_all_x_sg_out323), .sg_out324(_add_all_x_sg_out324), .sg_out325(_add_all_x_sg_out325), .sg_out326(_add_all_x_sg_out326), .sg_out327(_add_all_x_sg_out327), .sg_out328(_add_all_x_sg_out328), .sg_out329(_add_all_x_sg_out329), .sg_out330(_add_all_x_sg_out330), .sg_out331(_add_all_x_sg_out331), .sg_out332(_add_all_x_sg_out332), .sg_out333(_add_all_x_sg_out333), .sg_out334(_add_all_x_sg_out334), .sg_out335(_add_all_x_sg_out335), .sg_out336(_add_all_x_sg_out336), .sg_out337(_add_all_x_sg_out337), .sg_out338(_add_all_x_sg_out338), .sg_out339(_add_all_x_sg_out339), .sg_out340(_add_all_x_sg_out340), .sg_out341(_add_all_x_sg_out341), .sg_out342(_add_all_x_sg_out342), .sg_out343(_add_all_x_sg_out343), .sg_out344(_add_all_x_sg_out344), .sg_out345(_add_all_x_sg_out345), .sg_out346(_add_all_x_sg_out346), .sg_out347(_add_all_x_sg_out347), .sg_out348(_add_all_x_sg_out348), .sg_out349(_add_all_x_sg_out349), .sg_out350(_add_all_x_sg_out350), .sg_out353(_add_all_x_sg_out353), .sg_out354(_add_all_x_sg_out354), .sg_out355(_add_all_x_sg_out355), .sg_out356(_add_all_x_sg_out356), .sg_out357(_add_all_x_sg_out357), .sg_out358(_add_all_x_sg_out358), .sg_out359(_add_all_x_sg_out359), .sg_out360(_add_all_x_sg_out360), .sg_out361(_add_all_x_sg_out361), .sg_out362(_add_all_x_sg_out362), .sg_out363(_add_all_x_sg_out363), .sg_out364(_add_all_x_sg_out364), .sg_out365(_add_all_x_sg_out365), .sg_out366(_add_all_x_sg_out366), .sg_out367(_add_all_x_sg_out367), .sg_out368(_add_all_x_sg_out368), .sg_out369(_add_all_x_sg_out369), .sg_out370(_add_all_x_sg_out370), .sg_out371(_add_all_x_sg_out371), .sg_out372(_add_all_x_sg_out372), .sg_out373(_add_all_x_sg_out373), .sg_out374(_add_all_x_sg_out374), .sg_out375(_add_all_x_sg_out375), .sg_out376(_add_all_x_sg_out376), .sg_out377(_add_all_x_sg_out377), .sg_out378(_add_all_x_sg_out378), .sg_out379(_add_all_x_sg_out379), .sg_out380(_add_all_x_sg_out380), .sg_out381(_add_all_x_sg_out381), .sg_out382(_add_all_x_sg_out382), .sg_out385(_add_all_x_sg_out385), .sg_out386(_add_all_x_sg_out386), .sg_out387(_add_all_x_sg_out387), .sg_out388(_add_all_x_sg_out388), .sg_out389(_add_all_x_sg_out389), .sg_out390(_add_all_x_sg_out390), .sg_out391(_add_all_x_sg_out391), .sg_out392(_add_all_x_sg_out392), .sg_out393(_add_all_x_sg_out393), .sg_out394(_add_all_x_sg_out394), .sg_out395(_add_all_x_sg_out395), .sg_out396(_add_all_x_sg_out396), .sg_out397(_add_all_x_sg_out397), .sg_out398(_add_all_x_sg_out398), .sg_out399(_add_all_x_sg_out399), .sg_out400(_add_all_x_sg_out400), .sg_out401(_add_all_x_sg_out401), .sg_out402(_add_all_x_sg_out402), .sg_out403(_add_all_x_sg_out403), .sg_out404(_add_all_x_sg_out404), .sg_out405(_add_all_x_sg_out405), .sg_out406(_add_all_x_sg_out406), .sg_out407(_add_all_x_sg_out407), .sg_out408(_add_all_x_sg_out408), .sg_out409(_add_all_x_sg_out409), .sg_out410(_add_all_x_sg_out410), .sg_out411(_add_all_x_sg_out411), .sg_out412(_add_all_x_sg_out412), .sg_out413(_add_all_x_sg_out413), .sg_out414(_add_all_x_sg_out414), .sg_out417(_add_all_x_sg_out417), .sg_out418(_add_all_x_sg_out418), .sg_out419(_add_all_x_sg_out419), .sg_out420(_add_all_x_sg_out420), .sg_out421(_add_all_x_sg_out421), .sg_out422(_add_all_x_sg_out422), .sg_out423(_add_all_x_sg_out423), .sg_out424(_add_all_x_sg_out424), .sg_out425(_add_all_x_sg_out425), .sg_out426(_add_all_x_sg_out426), .sg_out427(_add_all_x_sg_out427), .sg_out428(_add_all_x_sg_out428), .sg_out429(_add_all_x_sg_out429), .sg_out430(_add_all_x_sg_out430), .sg_out431(_add_all_x_sg_out431), .sg_out432(_add_all_x_sg_out432), .sg_out433(_add_all_x_sg_out433), .sg_out434(_add_all_x_sg_out434), .sg_out435(_add_all_x_sg_out435), .sg_out436(_add_all_x_sg_out436), .sg_out437(_add_all_x_sg_out437), .sg_out438(_add_all_x_sg_out438), .sg_out439(_add_all_x_sg_out439), .sg_out440(_add_all_x_sg_out440), .sg_out441(_add_all_x_sg_out441), .sg_out442(_add_all_x_sg_out442), .sg_out443(_add_all_x_sg_out443), .sg_out444(_add_all_x_sg_out444), .sg_out445(_add_all_x_sg_out445), .sg_out446(_add_all_x_sg_out446), .sg_out449(_add_all_x_sg_out449), .sg_out450(_add_all_x_sg_out450), .sg_out451(_add_all_x_sg_out451), .sg_out452(_add_all_x_sg_out452), .sg_out453(_add_all_x_sg_out453), .sg_out454(_add_all_x_sg_out454), .sg_out455(_add_all_x_sg_out455), .sg_out456(_add_all_x_sg_out456), .sg_out457(_add_all_x_sg_out457), .sg_out458(_add_all_x_sg_out458), .sg_out459(_add_all_x_sg_out459), .sg_out460(_add_all_x_sg_out460), .sg_out461(_add_all_x_sg_out461), .sg_out462(_add_all_x_sg_out462), .sg_out463(_add_all_x_sg_out463), .sg_out464(_add_all_x_sg_out464), .sg_out465(_add_all_x_sg_out465), .sg_out466(_add_all_x_sg_out466), .sg_out467(_add_all_x_sg_out467), .sg_out468(_add_all_x_sg_out468), .sg_out469(_add_all_x_sg_out469), .sg_out470(_add_all_x_sg_out470), .sg_out471(_add_all_x_sg_out471), .sg_out472(_add_all_x_sg_out472), .sg_out473(_add_all_x_sg_out473), .sg_out474(_add_all_x_sg_out474), .sg_out475(_add_all_x_sg_out475), .sg_out476(_add_all_x_sg_out476), .sg_out477(_add_all_x_sg_out477), .sg_out478(_add_all_x_sg_out478), .sg_in33(_add_all_x_sg_in33), .sg_in34(_add_all_x_sg_in34), .sg_in35(_add_all_x_sg_in35), .sg_in36(_add_all_x_sg_in36), .sg_in37(_add_all_x_sg_in37), .sg_in38(_add_all_x_sg_in38), .sg_in39(_add_all_x_sg_in39), .sg_in40(_add_all_x_sg_in40), .sg_in41(_add_all_x_sg_in41), .sg_in42(_add_all_x_sg_in42), .sg_in43(_add_all_x_sg_in43), .sg_in44(_add_all_x_sg_in44), .sg_in45(_add_all_x_sg_in45), .sg_in46(_add_all_x_sg_in46), .sg_in47(_add_all_x_sg_in47), .sg_in48(_add_all_x_sg_in48), .sg_in49(_add_all_x_sg_in49), .sg_in50(_add_all_x_sg_in50), .sg_in51(_add_all_x_sg_in51), .sg_in52(_add_all_x_sg_in52), .sg_in53(_add_all_x_sg_in53), .sg_in54(_add_all_x_sg_in54), .sg_in55(_add_all_x_sg_in55), .sg_in56(_add_all_x_sg_in56), .sg_in57(_add_all_x_sg_in57), .sg_in58(_add_all_x_sg_in58), .sg_in59(_add_all_x_sg_in59), .sg_in60(_add_all_x_sg_in60), .sg_in61(_add_all_x_sg_in61), .sg_in62(_add_all_x_sg_in62), .sg_in65(_add_all_x_sg_in65), .sg_in66(_add_all_x_sg_in66), .sg_in67(_add_all_x_sg_in67), .sg_in68(_add_all_x_sg_in68), .sg_in69(_add_all_x_sg_in69), .sg_in70(_add_all_x_sg_in70), .sg_in71(_add_all_x_sg_in71), .sg_in72(_add_all_x_sg_in72), .sg_in73(_add_all_x_sg_in73), .sg_in74(_add_all_x_sg_in74), .sg_in75(_add_all_x_sg_in75), .sg_in76(_add_all_x_sg_in76), .sg_in77(_add_all_x_sg_in77), .sg_in78(_add_all_x_sg_in78), .sg_in79(_add_all_x_sg_in79), .sg_in80(_add_all_x_sg_in80), .sg_in81(_add_all_x_sg_in81), .sg_in82(_add_all_x_sg_in82), .sg_in83(_add_all_x_sg_in83), .sg_in84(_add_all_x_sg_in84), .sg_in85(_add_all_x_sg_in85), .sg_in86(_add_all_x_sg_in86), .sg_in87(_add_all_x_sg_in87), .sg_in88(_add_all_x_sg_in88), .sg_in89(_add_all_x_sg_in89), .sg_in90(_add_all_x_sg_in90), .sg_in91(_add_all_x_sg_in91), .sg_in92(_add_all_x_sg_in92), .sg_in93(_add_all_x_sg_in93), .sg_in94(_add_all_x_sg_in94), .sg_in97(_add_all_x_sg_in97), .sg_in98(_add_all_x_sg_in98), .sg_in99(_add_all_x_sg_in99), .sg_in100(_add_all_x_sg_in100), .sg_in101(_add_all_x_sg_in101), .sg_in102(_add_all_x_sg_in102), .sg_in103(_add_all_x_sg_in103), .sg_in104(_add_all_x_sg_in104), .sg_in105(_add_all_x_sg_in105), .sg_in106(_add_all_x_sg_in106), .sg_in107(_add_all_x_sg_in107), .sg_in108(_add_all_x_sg_in108), .sg_in109(_add_all_x_sg_in109), .sg_in110(_add_all_x_sg_in110), .sg_in111(_add_all_x_sg_in111), .sg_in112(_add_all_x_sg_in112), .sg_in113(_add_all_x_sg_in113), .sg_in114(_add_all_x_sg_in114), .sg_in115(_add_all_x_sg_in115), .sg_in116(_add_all_x_sg_in116), .sg_in117(_add_all_x_sg_in117), .sg_in118(_add_all_x_sg_in118), .sg_in119(_add_all_x_sg_in119), .sg_in120(_add_all_x_sg_in120), .sg_in121(_add_all_x_sg_in121), .sg_in122(_add_all_x_sg_in122), .sg_in123(_add_all_x_sg_in123), .sg_in124(_add_all_x_sg_in124), .sg_in125(_add_all_x_sg_in125), .sg_in126(_add_all_x_sg_in126), .sg_in129(_add_all_x_sg_in129), .sg_in130(_add_all_x_sg_in130), .sg_in131(_add_all_x_sg_in131), .sg_in132(_add_all_x_sg_in132), .sg_in133(_add_all_x_sg_in133), .sg_in134(_add_all_x_sg_in134), .sg_in135(_add_all_x_sg_in135), .sg_in136(_add_all_x_sg_in136), .sg_in137(_add_all_x_sg_in137), .sg_in138(_add_all_x_sg_in138), .sg_in139(_add_all_x_sg_in139), .sg_in140(_add_all_x_sg_in140), .sg_in141(_add_all_x_sg_in141), .sg_in142(_add_all_x_sg_in142), .sg_in143(_add_all_x_sg_in143), .sg_in144(_add_all_x_sg_in144), .sg_in145(_add_all_x_sg_in145), .sg_in146(_add_all_x_sg_in146), .sg_in147(_add_all_x_sg_in147), .sg_in148(_add_all_x_sg_in148), .sg_in149(_add_all_x_sg_in149), .sg_in150(_add_all_x_sg_in150), .sg_in151(_add_all_x_sg_in151), .sg_in152(_add_all_x_sg_in152), .sg_in153(_add_all_x_sg_in153), .sg_in154(_add_all_x_sg_in154), .sg_in155(_add_all_x_sg_in155), .sg_in156(_add_all_x_sg_in156), .sg_in157(_add_all_x_sg_in157), .sg_in158(_add_all_x_sg_in158), .sg_in161(_add_all_x_sg_in161), .sg_in162(_add_all_x_sg_in162), .sg_in163(_add_all_x_sg_in163), .sg_in164(_add_all_x_sg_in164), .sg_in165(_add_all_x_sg_in165), .sg_in166(_add_all_x_sg_in166), .sg_in167(_add_all_x_sg_in167), .sg_in168(_add_all_x_sg_in168), .sg_in169(_add_all_x_sg_in169), .sg_in170(_add_all_x_sg_in170), .sg_in171(_add_all_x_sg_in171), .sg_in172(_add_all_x_sg_in172), .sg_in173(_add_all_x_sg_in173), .sg_in174(_add_all_x_sg_in174), .sg_in175(_add_all_x_sg_in175), .sg_in176(_add_all_x_sg_in176), .sg_in177(_add_all_x_sg_in177), .sg_in178(_add_all_x_sg_in178), .sg_in179(_add_all_x_sg_in179), .sg_in180(_add_all_x_sg_in180), .sg_in181(_add_all_x_sg_in181), .sg_in182(_add_all_x_sg_in182), .sg_in183(_add_all_x_sg_in183), .sg_in184(_add_all_x_sg_in184), .sg_in185(_add_all_x_sg_in185), .sg_in186(_add_all_x_sg_in186), .sg_in187(_add_all_x_sg_in187), .sg_in188(_add_all_x_sg_in188), .sg_in189(_add_all_x_sg_in189), .sg_in190(_add_all_x_sg_in190), .sg_in193(_add_all_x_sg_in193), .sg_in194(_add_all_x_sg_in194), .sg_in195(_add_all_x_sg_in195), .sg_in196(_add_all_x_sg_in196), .sg_in197(_add_all_x_sg_in197), .sg_in198(_add_all_x_sg_in198), .sg_in199(_add_all_x_sg_in199), .sg_in200(_add_all_x_sg_in200), .sg_in201(_add_all_x_sg_in201), .sg_in202(_add_all_x_sg_in202), .sg_in203(_add_all_x_sg_in203), .sg_in204(_add_all_x_sg_in204), .sg_in205(_add_all_x_sg_in205), .sg_in206(_add_all_x_sg_in206), .sg_in207(_add_all_x_sg_in207), .sg_in208(_add_all_x_sg_in208), .sg_in209(_add_all_x_sg_in209), .sg_in210(_add_all_x_sg_in210), .sg_in211(_add_all_x_sg_in211), .sg_in212(_add_all_x_sg_in212), .sg_in213(_add_all_x_sg_in213), .sg_in214(_add_all_x_sg_in214), .sg_in215(_add_all_x_sg_in215), .sg_in216(_add_all_x_sg_in216), .sg_in217(_add_all_x_sg_in217), .sg_in218(_add_all_x_sg_in218), .sg_in219(_add_all_x_sg_in219), .sg_in220(_add_all_x_sg_in220), .sg_in221(_add_all_x_sg_in221), .sg_in222(_add_all_x_sg_in222), .sg_in225(_add_all_x_sg_in225), .sg_in226(_add_all_x_sg_in226), .sg_in227(_add_all_x_sg_in227), .sg_in228(_add_all_x_sg_in228), .sg_in229(_add_all_x_sg_in229), .sg_in230(_add_all_x_sg_in230), .sg_in231(_add_all_x_sg_in231), .sg_in232(_add_all_x_sg_in232), .sg_in233(_add_all_x_sg_in233), .sg_in234(_add_all_x_sg_in234), .sg_in235(_add_all_x_sg_in235), .sg_in236(_add_all_x_sg_in236), .sg_in237(_add_all_x_sg_in237), .sg_in238(_add_all_x_sg_in238), .sg_in239(_add_all_x_sg_in239), .sg_in240(_add_all_x_sg_in240), .sg_in241(_add_all_x_sg_in241), .sg_in242(_add_all_x_sg_in242), .sg_in243(_add_all_x_sg_in243), .sg_in244(_add_all_x_sg_in244), .sg_in245(_add_all_x_sg_in245), .sg_in246(_add_all_x_sg_in246), .sg_in247(_add_all_x_sg_in247), .sg_in248(_add_all_x_sg_in248), .sg_in249(_add_all_x_sg_in249), .sg_in250(_add_all_x_sg_in250), .sg_in251(_add_all_x_sg_in251), .sg_in252(_add_all_x_sg_in252), .sg_in253(_add_all_x_sg_in253), .sg_in254(_add_all_x_sg_in254), .sg_in257(_add_all_x_sg_in257), .sg_in258(_add_all_x_sg_in258), .sg_in259(_add_all_x_sg_in259), .sg_in260(_add_all_x_sg_in260), .sg_in261(_add_all_x_sg_in261), .sg_in262(_add_all_x_sg_in262), .sg_in263(_add_all_x_sg_in263), .sg_in264(_add_all_x_sg_in264), .sg_in265(_add_all_x_sg_in265), .sg_in266(_add_all_x_sg_in266), .sg_in267(_add_all_x_sg_in267), .sg_in268(_add_all_x_sg_in268), .sg_in269(_add_all_x_sg_in269), .sg_in270(_add_all_x_sg_in270), .sg_in271(_add_all_x_sg_in271), .sg_in272(_add_all_x_sg_in272), .sg_in273(_add_all_x_sg_in273), .sg_in274(_add_all_x_sg_in274), .sg_in275(_add_all_x_sg_in275), .sg_in276(_add_all_x_sg_in276), .sg_in277(_add_all_x_sg_in277), .sg_in278(_add_all_x_sg_in278), .sg_in279(_add_all_x_sg_in279), .sg_in280(_add_all_x_sg_in280), .sg_in281(_add_all_x_sg_in281), .sg_in282(_add_all_x_sg_in282), .sg_in283(_add_all_x_sg_in283), .sg_in284(_add_all_x_sg_in284), .sg_in285(_add_all_x_sg_in285), .sg_in286(_add_all_x_sg_in286), .sg_in289(_add_all_x_sg_in289), .sg_in290(_add_all_x_sg_in290), .sg_in291(_add_all_x_sg_in291), .sg_in292(_add_all_x_sg_in292), .sg_in293(_add_all_x_sg_in293), .sg_in294(_add_all_x_sg_in294), .sg_in295(_add_all_x_sg_in295), .sg_in296(_add_all_x_sg_in296), .sg_in297(_add_all_x_sg_in297), .sg_in298(_add_all_x_sg_in298), .sg_in299(_add_all_x_sg_in299), .sg_in300(_add_all_x_sg_in300), .sg_in301(_add_all_x_sg_in301), .sg_in302(_add_all_x_sg_in302), .sg_in303(_add_all_x_sg_in303), .sg_in304(_add_all_x_sg_in304), .sg_in305(_add_all_x_sg_in305), .sg_in306(_add_all_x_sg_in306), .sg_in307(_add_all_x_sg_in307), .sg_in308(_add_all_x_sg_in308), .sg_in309(_add_all_x_sg_in309), .sg_in310(_add_all_x_sg_in310), .sg_in311(_add_all_x_sg_in311), .sg_in312(_add_all_x_sg_in312), .sg_in313(_add_all_x_sg_in313), .sg_in314(_add_all_x_sg_in314), .sg_in315(_add_all_x_sg_in315), .sg_in316(_add_all_x_sg_in316), .sg_in317(_add_all_x_sg_in317), .sg_in318(_add_all_x_sg_in318), .sg_in321(_add_all_x_sg_in321), .sg_in322(_add_all_x_sg_in322), .sg_in323(_add_all_x_sg_in323), .sg_in324(_add_all_x_sg_in324), .sg_in325(_add_all_x_sg_in325), .sg_in326(_add_all_x_sg_in326), .sg_in327(_add_all_x_sg_in327), .sg_in328(_add_all_x_sg_in328), .sg_in329(_add_all_x_sg_in329), .sg_in330(_add_all_x_sg_in330), .sg_in331(_add_all_x_sg_in331), .sg_in332(_add_all_x_sg_in332), .sg_in333(_add_all_x_sg_in333), .sg_in334(_add_all_x_sg_in334), .sg_in335(_add_all_x_sg_in335), .sg_in336(_add_all_x_sg_in336), .sg_in337(_add_all_x_sg_in337), .sg_in338(_add_all_x_sg_in338), .sg_in339(_add_all_x_sg_in339), .sg_in340(_add_all_x_sg_in340), .sg_in341(_add_all_x_sg_in341), .sg_in342(_add_all_x_sg_in342), .sg_in343(_add_all_x_sg_in343), .sg_in344(_add_all_x_sg_in344), .sg_in345(_add_all_x_sg_in345), .sg_in346(_add_all_x_sg_in346), .sg_in347(_add_all_x_sg_in347), .sg_in348(_add_all_x_sg_in348), .sg_in349(_add_all_x_sg_in349), .sg_in350(_add_all_x_sg_in350), .sg_in353(_add_all_x_sg_in353), .sg_in354(_add_all_x_sg_in354), .sg_in355(_add_all_x_sg_in355), .sg_in356(_add_all_x_sg_in356), .sg_in357(_add_all_x_sg_in357), .sg_in358(_add_all_x_sg_in358), .sg_in359(_add_all_x_sg_in359), .sg_in360(_add_all_x_sg_in360), .sg_in361(_add_all_x_sg_in361), .sg_in362(_add_all_x_sg_in362), .sg_in363(_add_all_x_sg_in363), .sg_in364(_add_all_x_sg_in364), .sg_in365(_add_all_x_sg_in365), .sg_in366(_add_all_x_sg_in366), .sg_in367(_add_all_x_sg_in367), .sg_in368(_add_all_x_sg_in368), .sg_in369(_add_all_x_sg_in369), .sg_in370(_add_all_x_sg_in370), .sg_in371(_add_all_x_sg_in371), .sg_in372(_add_all_x_sg_in372), .sg_in373(_add_all_x_sg_in373), .sg_in374(_add_all_x_sg_in374), .sg_in375(_add_all_x_sg_in375), .sg_in376(_add_all_x_sg_in376), .sg_in377(_add_all_x_sg_in377), .sg_in378(_add_all_x_sg_in378), .sg_in379(_add_all_x_sg_in379), .sg_in380(_add_all_x_sg_in380), .sg_in381(_add_all_x_sg_in381), .sg_in382(_add_all_x_sg_in382), .sg_in385(_add_all_x_sg_in385), .sg_in386(_add_all_x_sg_in386), .sg_in387(_add_all_x_sg_in387), .sg_in388(_add_all_x_sg_in388), .sg_in389(_add_all_x_sg_in389), .sg_in390(_add_all_x_sg_in390), .sg_in391(_add_all_x_sg_in391), .sg_in392(_add_all_x_sg_in392), .sg_in393(_add_all_x_sg_in393), .sg_in394(_add_all_x_sg_in394), .sg_in395(_add_all_x_sg_in395), .sg_in396(_add_all_x_sg_in396), .sg_in397(_add_all_x_sg_in397), .sg_in398(_add_all_x_sg_in398), .sg_in399(_add_all_x_sg_in399), .sg_in400(_add_all_x_sg_in400), .sg_in401(_add_all_x_sg_in401), .sg_in402(_add_all_x_sg_in402), .sg_in403(_add_all_x_sg_in403), .sg_in404(_add_all_x_sg_in404), .sg_in405(_add_all_x_sg_in405), .sg_in406(_add_all_x_sg_in406), .sg_in407(_add_all_x_sg_in407), .sg_in408(_add_all_x_sg_in408), .sg_in409(_add_all_x_sg_in409), .sg_in410(_add_all_x_sg_in410), .sg_in411(_add_all_x_sg_in411), .sg_in412(_add_all_x_sg_in412), .sg_in413(_add_all_x_sg_in413), .sg_in414(_add_all_x_sg_in414), .sg_in417(_add_all_x_sg_in417), .sg_in418(_add_all_x_sg_in418), .sg_in419(_add_all_x_sg_in419), .sg_in420(_add_all_x_sg_in420), .sg_in421(_add_all_x_sg_in421), .sg_in422(_add_all_x_sg_in422), .sg_in423(_add_all_x_sg_in423), .sg_in424(_add_all_x_sg_in424), .sg_in425(_add_all_x_sg_in425), .sg_in426(_add_all_x_sg_in426), .sg_in427(_add_all_x_sg_in427), .sg_in428(_add_all_x_sg_in428), .sg_in429(_add_all_x_sg_in429), .sg_in430(_add_all_x_sg_in430), .sg_in431(_add_all_x_sg_in431), .sg_in432(_add_all_x_sg_in432), .sg_in433(_add_all_x_sg_in433), .sg_in434(_add_all_x_sg_in434), .sg_in435(_add_all_x_sg_in435), .sg_in436(_add_all_x_sg_in436), .sg_in437(_add_all_x_sg_in437), .sg_in438(_add_all_x_sg_in438), .sg_in439(_add_all_x_sg_in439), .sg_in440(_add_all_x_sg_in440), .sg_in441(_add_all_x_sg_in441), .sg_in442(_add_all_x_sg_in442), .sg_in443(_add_all_x_sg_in443), .sg_in444(_add_all_x_sg_in444), .sg_in445(_add_all_x_sg_in445), .sg_in446(_add_all_x_sg_in446), .sg_in449(_add_all_x_sg_in449), .sg_in450(_add_all_x_sg_in450), .sg_in451(_add_all_x_sg_in451), .sg_in452(_add_all_x_sg_in452), .sg_in453(_add_all_x_sg_in453), .sg_in454(_add_all_x_sg_in454), .sg_in455(_add_all_x_sg_in455), .sg_in456(_add_all_x_sg_in456), .sg_in457(_add_all_x_sg_in457), .sg_in458(_add_all_x_sg_in458), .sg_in459(_add_all_x_sg_in459), .sg_in460(_add_all_x_sg_in460), .sg_in461(_add_all_x_sg_in461), .sg_in462(_add_all_x_sg_in462), .sg_in463(_add_all_x_sg_in463), .sg_in464(_add_all_x_sg_in464), .sg_in465(_add_all_x_sg_in465), .sg_in466(_add_all_x_sg_in466), .sg_in467(_add_all_x_sg_in467), .sg_in468(_add_all_x_sg_in468), .sg_in469(_add_all_x_sg_in469), .sg_in470(_add_all_x_sg_in470), .sg_in471(_add_all_x_sg_in471), .sg_in472(_add_all_x_sg_in472), .sg_in473(_add_all_x_sg_in473), .sg_in474(_add_all_x_sg_in474), .sg_in475(_add_all_x_sg_in475), .sg_in476(_add_all_x_sg_in476), .sg_in477(_add_all_x_sg_in477), .sg_in478(_add_all_x_sg_in478), .data_out_index33(_add_all_x_data_out_index33), .data_out_index34(_add_all_x_data_out_index34), .data_out_index35(_add_all_x_data_out_index35), .data_out_index36(_add_all_x_data_out_index36), .data_out_index37(_add_all_x_data_out_index37), .data_out_index38(_add_all_x_data_out_index38), .data_out_index39(_add_all_x_data_out_index39), .data_out_index40(_add_all_x_data_out_index40), .data_out_index41(_add_all_x_data_out_index41), .data_out_index42(_add_all_x_data_out_index42), .data_out_index43(_add_all_x_data_out_index43), .data_out_index44(_add_all_x_data_out_index44), .data_out_index45(_add_all_x_data_out_index45), .data_out_index46(_add_all_x_data_out_index46), .data_out_index47(_add_all_x_data_out_index47), .data_out_index48(_add_all_x_data_out_index48), .data_out_index49(_add_all_x_data_out_index49), .data_out_index50(_add_all_x_data_out_index50), .data_out_index51(_add_all_x_data_out_index51), .data_out_index52(_add_all_x_data_out_index52), .data_out_index53(_add_all_x_data_out_index53), .data_out_index54(_add_all_x_data_out_index54), .data_out_index55(_add_all_x_data_out_index55), .data_out_index56(_add_all_x_data_out_index56), .data_out_index57(_add_all_x_data_out_index57), .data_out_index58(_add_all_x_data_out_index58), .data_out_index59(_add_all_x_data_out_index59), .data_out_index60(_add_all_x_data_out_index60), .data_out_index61(_add_all_x_data_out_index61), .data_out_index62(_add_all_x_data_out_index62), .data_out_index65(_add_all_x_data_out_index65), .data_out_index66(_add_all_x_data_out_index66), .data_out_index67(_add_all_x_data_out_index67), .data_out_index68(_add_all_x_data_out_index68), .data_out_index69(_add_all_x_data_out_index69), .data_out_index70(_add_all_x_data_out_index70), .data_out_index71(_add_all_x_data_out_index71), .data_out_index72(_add_all_x_data_out_index72), .data_out_index73(_add_all_x_data_out_index73), .data_out_index74(_add_all_x_data_out_index74), .data_out_index75(_add_all_x_data_out_index75), .data_out_index76(_add_all_x_data_out_index76), .data_out_index77(_add_all_x_data_out_index77), .data_out_index78(_add_all_x_data_out_index78), .data_out_index79(_add_all_x_data_out_index79), .data_out_index80(_add_all_x_data_out_index80), .data_out_index81(_add_all_x_data_out_index81), .data_out_index82(_add_all_x_data_out_index82), .data_out_index83(_add_all_x_data_out_index83), .data_out_index84(_add_all_x_data_out_index84), .data_out_index85(_add_all_x_data_out_index85), .data_out_index86(_add_all_x_data_out_index86), .data_out_index87(_add_all_x_data_out_index87), .data_out_index88(_add_all_x_data_out_index88), .data_out_index89(_add_all_x_data_out_index89), .data_out_index90(_add_all_x_data_out_index90), .data_out_index91(_add_all_x_data_out_index91), .data_out_index92(_add_all_x_data_out_index92), .data_out_index93(_add_all_x_data_out_index93), .data_out_index94(_add_all_x_data_out_index94), .data_out_index97(_add_all_x_data_out_index97), .data_out_index98(_add_all_x_data_out_index98), .data_out_index99(_add_all_x_data_out_index99), .data_out_index100(_add_all_x_data_out_index100), .data_out_index101(_add_all_x_data_out_index101), .data_out_index102(_add_all_x_data_out_index102), .data_out_index103(_add_all_x_data_out_index103), .data_out_index104(_add_all_x_data_out_index104), .data_out_index105(_add_all_x_data_out_index105), .data_out_index106(_add_all_x_data_out_index106), .data_out_index107(_add_all_x_data_out_index107), .data_out_index108(_add_all_x_data_out_index108), .data_out_index109(_add_all_x_data_out_index109), .data_out_index110(_add_all_x_data_out_index110), .data_out_index111(_add_all_x_data_out_index111), .data_out_index112(_add_all_x_data_out_index112), .data_out_index113(_add_all_x_data_out_index113), .data_out_index114(_add_all_x_data_out_index114), .data_out_index115(_add_all_x_data_out_index115), .data_out_index116(_add_all_x_data_out_index116), .data_out_index117(_add_all_x_data_out_index117), .data_out_index118(_add_all_x_data_out_index118), .data_out_index119(_add_all_x_data_out_index119), .data_out_index120(_add_all_x_data_out_index120), .data_out_index121(_add_all_x_data_out_index121), .data_out_index122(_add_all_x_data_out_index122), .data_out_index123(_add_all_x_data_out_index123), .data_out_index124(_add_all_x_data_out_index124), .data_out_index125(_add_all_x_data_out_index125), .data_out_index126(_add_all_x_data_out_index126), .data_out_index129(_add_all_x_data_out_index129), .data_out_index130(_add_all_x_data_out_index130), .data_out_index131(_add_all_x_data_out_index131), .data_out_index132(_add_all_x_data_out_index132), .data_out_index133(_add_all_x_data_out_index133), .data_out_index134(_add_all_x_data_out_index134), .data_out_index135(_add_all_x_data_out_index135), .data_out_index136(_add_all_x_data_out_index136), .data_out_index137(_add_all_x_data_out_index137), .data_out_index138(_add_all_x_data_out_index138), .data_out_index139(_add_all_x_data_out_index139), .data_out_index140(_add_all_x_data_out_index140), .data_out_index141(_add_all_x_data_out_index141), .data_out_index142(_add_all_x_data_out_index142), .data_out_index143(_add_all_x_data_out_index143), .data_out_index144(_add_all_x_data_out_index144), .data_out_index145(_add_all_x_data_out_index145), .data_out_index146(_add_all_x_data_out_index146), .data_out_index147(_add_all_x_data_out_index147), .data_out_index148(_add_all_x_data_out_index148), .data_out_index149(_add_all_x_data_out_index149), .data_out_index150(_add_all_x_data_out_index150), .data_out_index151(_add_all_x_data_out_index151), .data_out_index152(_add_all_x_data_out_index152), .data_out_index153(_add_all_x_data_out_index153), .data_out_index154(_add_all_x_data_out_index154), .data_out_index155(_add_all_x_data_out_index155), .data_out_index156(_add_all_x_data_out_index156), .data_out_index157(_add_all_x_data_out_index157), .data_out_index158(_add_all_x_data_out_index158), .data_out_index161(_add_all_x_data_out_index161), .data_out_index162(_add_all_x_data_out_index162), .data_out_index163(_add_all_x_data_out_index163), .data_out_index164(_add_all_x_data_out_index164), .data_out_index165(_add_all_x_data_out_index165), .data_out_index166(_add_all_x_data_out_index166), .data_out_index167(_add_all_x_data_out_index167), .data_out_index168(_add_all_x_data_out_index168), .data_out_index169(_add_all_x_data_out_index169), .data_out_index170(_add_all_x_data_out_index170), .data_out_index171(_add_all_x_data_out_index171), .data_out_index172(_add_all_x_data_out_index172), .data_out_index173(_add_all_x_data_out_index173), .data_out_index174(_add_all_x_data_out_index174), .data_out_index175(_add_all_x_data_out_index175), .data_out_index176(_add_all_x_data_out_index176), .data_out_index177(_add_all_x_data_out_index177), .data_out_index178(_add_all_x_data_out_index178), .data_out_index179(_add_all_x_data_out_index179), .data_out_index180(_add_all_x_data_out_index180), .data_out_index181(_add_all_x_data_out_index181), .data_out_index182(_add_all_x_data_out_index182), .data_out_index183(_add_all_x_data_out_index183), .data_out_index184(_add_all_x_data_out_index184), .data_out_index185(_add_all_x_data_out_index185), .data_out_index186(_add_all_x_data_out_index186), .data_out_index187(_add_all_x_data_out_index187), .data_out_index188(_add_all_x_data_out_index188), .data_out_index189(_add_all_x_data_out_index189), .data_out_index190(_add_all_x_data_out_index190), .data_out_index193(_add_all_x_data_out_index193), .data_out_index194(_add_all_x_data_out_index194), .data_out_index195(_add_all_x_data_out_index195), .data_out_index196(_add_all_x_data_out_index196), .data_out_index197(_add_all_x_data_out_index197), .data_out_index198(_add_all_x_data_out_index198), .data_out_index199(_add_all_x_data_out_index199), .data_out_index200(_add_all_x_data_out_index200), .data_out_index201(_add_all_x_data_out_index201), .data_out_index202(_add_all_x_data_out_index202), .data_out_index203(_add_all_x_data_out_index203), .data_out_index204(_add_all_x_data_out_index204), .data_out_index205(_add_all_x_data_out_index205), .data_out_index206(_add_all_x_data_out_index206), .data_out_index207(_add_all_x_data_out_index207), .data_out_index208(_add_all_x_data_out_index208), .data_out_index209(_add_all_x_data_out_index209), .data_out_index210(_add_all_x_data_out_index210), .data_out_index211(_add_all_x_data_out_index211), .data_out_index212(_add_all_x_data_out_index212), .data_out_index213(_add_all_x_data_out_index213), .data_out_index214(_add_all_x_data_out_index214), .data_out_index215(_add_all_x_data_out_index215), .data_out_index216(_add_all_x_data_out_index216), .data_out_index217(_add_all_x_data_out_index217), .data_out_index218(_add_all_x_data_out_index218), .data_out_index219(_add_all_x_data_out_index219), .data_out_index220(_add_all_x_data_out_index220), .data_out_index221(_add_all_x_data_out_index221), .data_out_index222(_add_all_x_data_out_index222), .data_out_index225(_add_all_x_data_out_index225), .data_out_index226(_add_all_x_data_out_index226), .data_out_index227(_add_all_x_data_out_index227), .data_out_index228(_add_all_x_data_out_index228), .data_out_index229(_add_all_x_data_out_index229), .data_out_index230(_add_all_x_data_out_index230), .data_out_index231(_add_all_x_data_out_index231), .data_out_index232(_add_all_x_data_out_index232), .data_out_index233(_add_all_x_data_out_index233), .data_out_index234(_add_all_x_data_out_index234), .data_out_index235(_add_all_x_data_out_index235), .data_out_index236(_add_all_x_data_out_index236), .data_out_index237(_add_all_x_data_out_index237), .data_out_index238(_add_all_x_data_out_index238), .data_out_index239(_add_all_x_data_out_index239), .data_out_index240(_add_all_x_data_out_index240), .data_out_index241(_add_all_x_data_out_index241), .data_out_index242(_add_all_x_data_out_index242), .data_out_index243(_add_all_x_data_out_index243), .data_out_index244(_add_all_x_data_out_index244), .data_out_index245(_add_all_x_data_out_index245), .data_out_index246(_add_all_x_data_out_index246), .data_out_index247(_add_all_x_data_out_index247), .data_out_index248(_add_all_x_data_out_index248), .data_out_index249(_add_all_x_data_out_index249), .data_out_index250(_add_all_x_data_out_index250), .data_out_index251(_add_all_x_data_out_index251), .data_out_index252(_add_all_x_data_out_index252), .data_out_index253(_add_all_x_data_out_index253), .data_out_index254(_add_all_x_data_out_index254), .data_out_index257(_add_all_x_data_out_index257), .data_out_index258(_add_all_x_data_out_index258), .data_out_index259(_add_all_x_data_out_index259), .data_out_index260(_add_all_x_data_out_index260), .data_out_index261(_add_all_x_data_out_index261), .data_out_index262(_add_all_x_data_out_index262), .data_out_index263(_add_all_x_data_out_index263), .data_out_index264(_add_all_x_data_out_index264), .data_out_index265(_add_all_x_data_out_index265), .data_out_index266(_add_all_x_data_out_index266), .data_out_index267(_add_all_x_data_out_index267), .data_out_index268(_add_all_x_data_out_index268), .data_out_index269(_add_all_x_data_out_index269), .data_out_index270(_add_all_x_data_out_index270), .data_out_index271(_add_all_x_data_out_index271), .data_out_index272(_add_all_x_data_out_index272), .data_out_index273(_add_all_x_data_out_index273), .data_out_index274(_add_all_x_data_out_index274), .data_out_index275(_add_all_x_data_out_index275), .data_out_index276(_add_all_x_data_out_index276), .data_out_index277(_add_all_x_data_out_index277), .data_out_index278(_add_all_x_data_out_index278), .data_out_index279(_add_all_x_data_out_index279), .data_out_index280(_add_all_x_data_out_index280), .data_out_index281(_add_all_x_data_out_index281), .data_out_index282(_add_all_x_data_out_index282), .data_out_index283(_add_all_x_data_out_index283), .data_out_index284(_add_all_x_data_out_index284), .data_out_index285(_add_all_x_data_out_index285), .data_out_index286(_add_all_x_data_out_index286), .data_out_index289(_add_all_x_data_out_index289), .data_out_index290(_add_all_x_data_out_index290), .data_out_index291(_add_all_x_data_out_index291), .data_out_index292(_add_all_x_data_out_index292), .data_out_index293(_add_all_x_data_out_index293), .data_out_index294(_add_all_x_data_out_index294), .data_out_index295(_add_all_x_data_out_index295), .data_out_index296(_add_all_x_data_out_index296), .data_out_index297(_add_all_x_data_out_index297), .data_out_index298(_add_all_x_data_out_index298), .data_out_index299(_add_all_x_data_out_index299), .data_out_index300(_add_all_x_data_out_index300), .data_out_index301(_add_all_x_data_out_index301), .data_out_index302(_add_all_x_data_out_index302), .data_out_index303(_add_all_x_data_out_index303), .data_out_index304(_add_all_x_data_out_index304), .data_out_index305(_add_all_x_data_out_index305), .data_out_index306(_add_all_x_data_out_index306), .data_out_index307(_add_all_x_data_out_index307), .data_out_index308(_add_all_x_data_out_index308), .data_out_index309(_add_all_x_data_out_index309), .data_out_index310(_add_all_x_data_out_index310), .data_out_index311(_add_all_x_data_out_index311), .data_out_index312(_add_all_x_data_out_index312), .data_out_index313(_add_all_x_data_out_index313), .data_out_index314(_add_all_x_data_out_index314), .data_out_index315(_add_all_x_data_out_index315), .data_out_index316(_add_all_x_data_out_index316), .data_out_index317(_add_all_x_data_out_index317), .data_out_index318(_add_all_x_data_out_index318), .data_out_index321(_add_all_x_data_out_index321), .data_out_index322(_add_all_x_data_out_index322), .data_out_index323(_add_all_x_data_out_index323), .data_out_index324(_add_all_x_data_out_index324), .data_out_index325(_add_all_x_data_out_index325), .data_out_index326(_add_all_x_data_out_index326), .data_out_index327(_add_all_x_data_out_index327), .data_out_index328(_add_all_x_data_out_index328), .data_out_index329(_add_all_x_data_out_index329), .data_out_index330(_add_all_x_data_out_index330), .data_out_index331(_add_all_x_data_out_index331), .data_out_index332(_add_all_x_data_out_index332), .data_out_index333(_add_all_x_data_out_index333), .data_out_index334(_add_all_x_data_out_index334), .data_out_index335(_add_all_x_data_out_index335), .data_out_index336(_add_all_x_data_out_index336), .data_out_index337(_add_all_x_data_out_index337), .data_out_index338(_add_all_x_data_out_index338), .data_out_index339(_add_all_x_data_out_index339), .data_out_index340(_add_all_x_data_out_index340), .data_out_index341(_add_all_x_data_out_index341), .data_out_index342(_add_all_x_data_out_index342), .data_out_index343(_add_all_x_data_out_index343), .data_out_index344(_add_all_x_data_out_index344), .data_out_index345(_add_all_x_data_out_index345), .data_out_index346(_add_all_x_data_out_index346), .data_out_index347(_add_all_x_data_out_index347), .data_out_index348(_add_all_x_data_out_index348), .data_out_index349(_add_all_x_data_out_index349), .data_out_index350(_add_all_x_data_out_index350), .data_out_index353(_add_all_x_data_out_index353), .data_out_index354(_add_all_x_data_out_index354), .data_out_index355(_add_all_x_data_out_index355), .data_out_index356(_add_all_x_data_out_index356), .data_out_index357(_add_all_x_data_out_index357), .data_out_index358(_add_all_x_data_out_index358), .data_out_index359(_add_all_x_data_out_index359), .data_out_index360(_add_all_x_data_out_index360), .data_out_index361(_add_all_x_data_out_index361), .data_out_index362(_add_all_x_data_out_index362), .data_out_index363(_add_all_x_data_out_index363), .data_out_index364(_add_all_x_data_out_index364), .data_out_index365(_add_all_x_data_out_index365), .data_out_index366(_add_all_x_data_out_index366), .data_out_index367(_add_all_x_data_out_index367), .data_out_index368(_add_all_x_data_out_index368), .data_out_index369(_add_all_x_data_out_index369), .data_out_index370(_add_all_x_data_out_index370), .data_out_index371(_add_all_x_data_out_index371), .data_out_index372(_add_all_x_data_out_index372), .data_out_index373(_add_all_x_data_out_index373), .data_out_index374(_add_all_x_data_out_index374), .data_out_index375(_add_all_x_data_out_index375), .data_out_index376(_add_all_x_data_out_index376), .data_out_index377(_add_all_x_data_out_index377), .data_out_index378(_add_all_x_data_out_index378), .data_out_index379(_add_all_x_data_out_index379), .data_out_index380(_add_all_x_data_out_index380), .data_out_index381(_add_all_x_data_out_index381), .data_out_index382(_add_all_x_data_out_index382), .data_out_index385(_add_all_x_data_out_index385), .data_out_index386(_add_all_x_data_out_index386), .data_out_index387(_add_all_x_data_out_index387), .data_out_index388(_add_all_x_data_out_index388), .data_out_index389(_add_all_x_data_out_index389), .data_out_index390(_add_all_x_data_out_index390), .data_out_index391(_add_all_x_data_out_index391), .data_out_index392(_add_all_x_data_out_index392), .data_out_index393(_add_all_x_data_out_index393), .data_out_index394(_add_all_x_data_out_index394), .data_out_index395(_add_all_x_data_out_index395), .data_out_index396(_add_all_x_data_out_index396), .data_out_index397(_add_all_x_data_out_index397), .data_out_index398(_add_all_x_data_out_index398), .data_out_index399(_add_all_x_data_out_index399), .data_out_index400(_add_all_x_data_out_index400), .data_out_index401(_add_all_x_data_out_index401), .data_out_index402(_add_all_x_data_out_index402), .data_out_index403(_add_all_x_data_out_index403), .data_out_index404(_add_all_x_data_out_index404), .data_out_index405(_add_all_x_data_out_index405), .data_out_index406(_add_all_x_data_out_index406), .data_out_index407(_add_all_x_data_out_index407), .data_out_index408(_add_all_x_data_out_index408), .data_out_index409(_add_all_x_data_out_index409), .data_out_index410(_add_all_x_data_out_index410), .data_out_index411(_add_all_x_data_out_index411), .data_out_index412(_add_all_x_data_out_index412), .data_out_index413(_add_all_x_data_out_index413), .data_out_index414(_add_all_x_data_out_index414), .data_out_index417(_add_all_x_data_out_index417), .data_out_index418(_add_all_x_data_out_index418), .data_out_index419(_add_all_x_data_out_index419), .data_out_index420(_add_all_x_data_out_index420), .data_out_index421(_add_all_x_data_out_index421), .data_out_index422(_add_all_x_data_out_index422), .data_out_index423(_add_all_x_data_out_index423), .data_out_index424(_add_all_x_data_out_index424), .data_out_index425(_add_all_x_data_out_index425), .data_out_index426(_add_all_x_data_out_index426), .data_out_index427(_add_all_x_data_out_index427), .data_out_index428(_add_all_x_data_out_index428), .data_out_index429(_add_all_x_data_out_index429), .data_out_index430(_add_all_x_data_out_index430), .data_out_index431(_add_all_x_data_out_index431), .data_out_index432(_add_all_x_data_out_index432), .data_out_index433(_add_all_x_data_out_index433), .data_out_index434(_add_all_x_data_out_index434), .data_out_index435(_add_all_x_data_out_index435), .data_out_index436(_add_all_x_data_out_index436), .data_out_index437(_add_all_x_data_out_index437), .data_out_index438(_add_all_x_data_out_index438), .data_out_index439(_add_all_x_data_out_index439), .data_out_index440(_add_all_x_data_out_index440), .data_out_index441(_add_all_x_data_out_index441), .data_out_index442(_add_all_x_data_out_index442), .data_out_index443(_add_all_x_data_out_index443), .data_out_index444(_add_all_x_data_out_index444), .data_out_index445(_add_all_x_data_out_index445), .data_out_index446(_add_all_x_data_out_index446), .data_out_index449(_add_all_x_data_out_index449), .data_out_index450(_add_all_x_data_out_index450), .data_out_index451(_add_all_x_data_out_index451), .data_out_index452(_add_all_x_data_out_index452), .data_out_index453(_add_all_x_data_out_index453), .data_out_index454(_add_all_x_data_out_index454), .data_out_index455(_add_all_x_data_out_index455), .data_out_index456(_add_all_x_data_out_index456), .data_out_index457(_add_all_x_data_out_index457), .data_out_index458(_add_all_x_data_out_index458), .data_out_index459(_add_all_x_data_out_index459), .data_out_index460(_add_all_x_data_out_index460), .data_out_index461(_add_all_x_data_out_index461), .data_out_index462(_add_all_x_data_out_index462), .data_out_index463(_add_all_x_data_out_index463), .data_out_index464(_add_all_x_data_out_index464), .data_out_index465(_add_all_x_data_out_index465), .data_out_index466(_add_all_x_data_out_index466), .data_out_index467(_add_all_x_data_out_index467), .data_out_index468(_add_all_x_data_out_index468), .data_out_index469(_add_all_x_data_out_index469), .data_out_index470(_add_all_x_data_out_index470), .data_out_index471(_add_all_x_data_out_index471), .data_out_index472(_add_all_x_data_out_index472), .data_out_index473(_add_all_x_data_out_index473), .data_out_index474(_add_all_x_data_out_index474), .data_out_index475(_add_all_x_data_out_index475), .data_out_index476(_add_all_x_data_out_index476), .data_out_index477(_add_all_x_data_out_index477), .data_out_index478(_add_all_x_data_out_index478), .data_out33(_add_all_x_data_out33), .data_out34(_add_all_x_data_out34), .data_out35(_add_all_x_data_out35), .data_out36(_add_all_x_data_out36), .data_out37(_add_all_x_data_out37), .data_out38(_add_all_x_data_out38), .data_out39(_add_all_x_data_out39), .data_out40(_add_all_x_data_out40), .data_out41(_add_all_x_data_out41), .data_out42(_add_all_x_data_out42), .data_out43(_add_all_x_data_out43), .data_out44(_add_all_x_data_out44), .data_out45(_add_all_x_data_out45), .data_out46(_add_all_x_data_out46), .data_out47(_add_all_x_data_out47), .data_out48(_add_all_x_data_out48), .data_out49(_add_all_x_data_out49), .data_out50(_add_all_x_data_out50), .data_out51(_add_all_x_data_out51), .data_out52(_add_all_x_data_out52), .data_out53(_add_all_x_data_out53), .data_out54(_add_all_x_data_out54), .data_out55(_add_all_x_data_out55), .data_out56(_add_all_x_data_out56), .data_out57(_add_all_x_data_out57), .data_out58(_add_all_x_data_out58), .data_out59(_add_all_x_data_out59), .data_out60(_add_all_x_data_out60), .data_out61(_add_all_x_data_out61), .data_out62(_add_all_x_data_out62), .data_out65(_add_all_x_data_out65), .data_out66(_add_all_x_data_out66), .data_out67(_add_all_x_data_out67), .data_out68(_add_all_x_data_out68), .data_out69(_add_all_x_data_out69), .data_out70(_add_all_x_data_out70), .data_out71(_add_all_x_data_out71), .data_out72(_add_all_x_data_out72), .data_out73(_add_all_x_data_out73), .data_out74(_add_all_x_data_out74), .data_out75(_add_all_x_data_out75), .data_out76(_add_all_x_data_out76), .data_out77(_add_all_x_data_out77), .data_out78(_add_all_x_data_out78), .data_out79(_add_all_x_data_out79), .data_out80(_add_all_x_data_out80), .data_out81(_add_all_x_data_out81), .data_out82(_add_all_x_data_out82), .data_out83(_add_all_x_data_out83), .data_out84(_add_all_x_data_out84), .data_out85(_add_all_x_data_out85), .data_out86(_add_all_x_data_out86), .data_out87(_add_all_x_data_out87), .data_out88(_add_all_x_data_out88), .data_out89(_add_all_x_data_out89), .data_out90(_add_all_x_data_out90), .data_out91(_add_all_x_data_out91), .data_out92(_add_all_x_data_out92), .data_out93(_add_all_x_data_out93), .data_out94(_add_all_x_data_out94), .data_out97(_add_all_x_data_out97), .data_out98(_add_all_x_data_out98), .data_out99(_add_all_x_data_out99), .data_out100(_add_all_x_data_out100), .data_out101(_add_all_x_data_out101), .data_out102(_add_all_x_data_out102), .data_out103(_add_all_x_data_out103), .data_out104(_add_all_x_data_out104), .data_out105(_add_all_x_data_out105), .data_out106(_add_all_x_data_out106), .data_out107(_add_all_x_data_out107), .data_out108(_add_all_x_data_out108), .data_out109(_add_all_x_data_out109), .data_out110(_add_all_x_data_out110), .data_out111(_add_all_x_data_out111), .data_out112(_add_all_x_data_out112), .data_out113(_add_all_x_data_out113), .data_out114(_add_all_x_data_out114), .data_out115(_add_all_x_data_out115), .data_out116(_add_all_x_data_out116), .data_out117(_add_all_x_data_out117), .data_out118(_add_all_x_data_out118), .data_out119(_add_all_x_data_out119), .data_out120(_add_all_x_data_out120), .data_out121(_add_all_x_data_out121), .data_out122(_add_all_x_data_out122), .data_out123(_add_all_x_data_out123), .data_out124(_add_all_x_data_out124), .data_out125(_add_all_x_data_out125), .data_out126(_add_all_x_data_out126), .data_out129(_add_all_x_data_out129), .data_out130(_add_all_x_data_out130), .data_out131(_add_all_x_data_out131), .data_out132(_add_all_x_data_out132), .data_out133(_add_all_x_data_out133), .data_out134(_add_all_x_data_out134), .data_out135(_add_all_x_data_out135), .data_out136(_add_all_x_data_out136), .data_out137(_add_all_x_data_out137), .data_out138(_add_all_x_data_out138), .data_out139(_add_all_x_data_out139), .data_out140(_add_all_x_data_out140), .data_out141(_add_all_x_data_out141), .data_out142(_add_all_x_data_out142), .data_out143(_add_all_x_data_out143), .data_out144(_add_all_x_data_out144), .data_out145(_add_all_x_data_out145), .data_out146(_add_all_x_data_out146), .data_out147(_add_all_x_data_out147), .data_out148(_add_all_x_data_out148), .data_out149(_add_all_x_data_out149), .data_out150(_add_all_x_data_out150), .data_out151(_add_all_x_data_out151), .data_out152(_add_all_x_data_out152), .data_out153(_add_all_x_data_out153), .data_out154(_add_all_x_data_out154), .data_out155(_add_all_x_data_out155), .data_out156(_add_all_x_data_out156), .data_out157(_add_all_x_data_out157), .data_out158(_add_all_x_data_out158), .data_out161(_add_all_x_data_out161), .data_out162(_add_all_x_data_out162), .data_out163(_add_all_x_data_out163), .data_out164(_add_all_x_data_out164), .data_out165(_add_all_x_data_out165), .data_out166(_add_all_x_data_out166), .data_out167(_add_all_x_data_out167), .data_out168(_add_all_x_data_out168), .data_out169(_add_all_x_data_out169), .data_out170(_add_all_x_data_out170), .data_out171(_add_all_x_data_out171), .data_out172(_add_all_x_data_out172), .data_out173(_add_all_x_data_out173), .data_out174(_add_all_x_data_out174), .data_out175(_add_all_x_data_out175), .data_out176(_add_all_x_data_out176), .data_out177(_add_all_x_data_out177), .data_out178(_add_all_x_data_out178), .data_out179(_add_all_x_data_out179), .data_out180(_add_all_x_data_out180), .data_out181(_add_all_x_data_out181), .data_out182(_add_all_x_data_out182), .data_out183(_add_all_x_data_out183), .data_out184(_add_all_x_data_out184), .data_out185(_add_all_x_data_out185), .data_out186(_add_all_x_data_out186), .data_out187(_add_all_x_data_out187), .data_out188(_add_all_x_data_out188), .data_out189(_add_all_x_data_out189), .data_out190(_add_all_x_data_out190), .data_out193(_add_all_x_data_out193), .data_out194(_add_all_x_data_out194), .data_out195(_add_all_x_data_out195), .data_out196(_add_all_x_data_out196), .data_out197(_add_all_x_data_out197), .data_out198(_add_all_x_data_out198), .data_out199(_add_all_x_data_out199), .data_out200(_add_all_x_data_out200), .data_out201(_add_all_x_data_out201), .data_out202(_add_all_x_data_out202), .data_out203(_add_all_x_data_out203), .data_out204(_add_all_x_data_out204), .data_out205(_add_all_x_data_out205), .data_out206(_add_all_x_data_out206), .data_out207(_add_all_x_data_out207), .data_out208(_add_all_x_data_out208), .data_out209(_add_all_x_data_out209), .data_out210(_add_all_x_data_out210), .data_out211(_add_all_x_data_out211), .data_out212(_add_all_x_data_out212), .data_out213(_add_all_x_data_out213), .data_out214(_add_all_x_data_out214), .data_out215(_add_all_x_data_out215), .data_out216(_add_all_x_data_out216), .data_out217(_add_all_x_data_out217), .data_out218(_add_all_x_data_out218), .data_out219(_add_all_x_data_out219), .data_out220(_add_all_x_data_out220), .data_out221(_add_all_x_data_out221), .data_out222(_add_all_x_data_out222), .data_out225(_add_all_x_data_out225), .data_out226(_add_all_x_data_out226), .data_out227(_add_all_x_data_out227), .data_out228(_add_all_x_data_out228), .data_out229(_add_all_x_data_out229), .data_out230(_add_all_x_data_out230), .data_out231(_add_all_x_data_out231), .data_out232(_add_all_x_data_out232), .data_out233(_add_all_x_data_out233), .data_out234(_add_all_x_data_out234), .data_out235(_add_all_x_data_out235), .data_out236(_add_all_x_data_out236), .data_out237(_add_all_x_data_out237), .data_out238(_add_all_x_data_out238), .data_out239(_add_all_x_data_out239), .data_out240(_add_all_x_data_out240), .data_out241(_add_all_x_data_out241), .data_out242(_add_all_x_data_out242), .data_out243(_add_all_x_data_out243), .data_out244(_add_all_x_data_out244), .data_out245(_add_all_x_data_out245), .data_out246(_add_all_x_data_out246), .data_out247(_add_all_x_data_out247), .data_out248(_add_all_x_data_out248), .data_out249(_add_all_x_data_out249), .data_out250(_add_all_x_data_out250), .data_out251(_add_all_x_data_out251), .data_out252(_add_all_x_data_out252), .data_out253(_add_all_x_data_out253), .data_out254(_add_all_x_data_out254), .data_out257(_add_all_x_data_out257), .data_out258(_add_all_x_data_out258), .data_out259(_add_all_x_data_out259), .data_out260(_add_all_x_data_out260), .data_out261(_add_all_x_data_out261), .data_out262(_add_all_x_data_out262), .data_out263(_add_all_x_data_out263), .data_out264(_add_all_x_data_out264), .data_out265(_add_all_x_data_out265), .data_out266(_add_all_x_data_out266), .data_out267(_add_all_x_data_out267), .data_out268(_add_all_x_data_out268), .data_out269(_add_all_x_data_out269), .data_out270(_add_all_x_data_out270), .data_out271(_add_all_x_data_out271), .data_out272(_add_all_x_data_out272), .data_out273(_add_all_x_data_out273), .data_out274(_add_all_x_data_out274), .data_out275(_add_all_x_data_out275), .data_out276(_add_all_x_data_out276), .data_out277(_add_all_x_data_out277), .data_out278(_add_all_x_data_out278), .data_out279(_add_all_x_data_out279), .data_out280(_add_all_x_data_out280), .data_out281(_add_all_x_data_out281), .data_out282(_add_all_x_data_out282), .data_out283(_add_all_x_data_out283), .data_out284(_add_all_x_data_out284), .data_out285(_add_all_x_data_out285), .data_out286(_add_all_x_data_out286), .data_out289(_add_all_x_data_out289), .data_out290(_add_all_x_data_out290), .data_out291(_add_all_x_data_out291), .data_out292(_add_all_x_data_out292), .data_out293(_add_all_x_data_out293), .data_out294(_add_all_x_data_out294), .data_out295(_add_all_x_data_out295), .data_out296(_add_all_x_data_out296), .data_out297(_add_all_x_data_out297), .data_out298(_add_all_x_data_out298), .data_out299(_add_all_x_data_out299), .data_out300(_add_all_x_data_out300), .data_out301(_add_all_x_data_out301), .data_out302(_add_all_x_data_out302), .data_out303(_add_all_x_data_out303), .data_out304(_add_all_x_data_out304), .data_out305(_add_all_x_data_out305), .data_out306(_add_all_x_data_out306), .data_out307(_add_all_x_data_out307), .data_out308(_add_all_x_data_out308), .data_out309(_add_all_x_data_out309), .data_out310(_add_all_x_data_out310), .data_out311(_add_all_x_data_out311), .data_out312(_add_all_x_data_out312), .data_out313(_add_all_x_data_out313), .data_out314(_add_all_x_data_out314), .data_out315(_add_all_x_data_out315), .data_out316(_add_all_x_data_out316), .data_out317(_add_all_x_data_out317), .data_out318(_add_all_x_data_out318), .data_out321(_add_all_x_data_out321), .data_out322(_add_all_x_data_out322), .data_out323(_add_all_x_data_out323), .data_out324(_add_all_x_data_out324), .data_out325(_add_all_x_data_out325), .data_out326(_add_all_x_data_out326), .data_out327(_add_all_x_data_out327), .data_out328(_add_all_x_data_out328), .data_out329(_add_all_x_data_out329), .data_out330(_add_all_x_data_out330), .data_out331(_add_all_x_data_out331), .data_out332(_add_all_x_data_out332), .data_out333(_add_all_x_data_out333), .data_out334(_add_all_x_data_out334), .data_out335(_add_all_x_data_out335), .data_out336(_add_all_x_data_out336), .data_out337(_add_all_x_data_out337), .data_out338(_add_all_x_data_out338), .data_out339(_add_all_x_data_out339), .data_out340(_add_all_x_data_out340), .data_out341(_add_all_x_data_out341), .data_out342(_add_all_x_data_out342), .data_out343(_add_all_x_data_out343), .data_out344(_add_all_x_data_out344), .data_out345(_add_all_x_data_out345), .data_out346(_add_all_x_data_out346), .data_out347(_add_all_x_data_out347), .data_out348(_add_all_x_data_out348), .data_out349(_add_all_x_data_out349), .data_out350(_add_all_x_data_out350), .data_out353(_add_all_x_data_out353), .data_out354(_add_all_x_data_out354), .data_out355(_add_all_x_data_out355), .data_out356(_add_all_x_data_out356), .data_out357(_add_all_x_data_out357), .data_out358(_add_all_x_data_out358), .data_out359(_add_all_x_data_out359), .data_out360(_add_all_x_data_out360), .data_out361(_add_all_x_data_out361), .data_out362(_add_all_x_data_out362), .data_out363(_add_all_x_data_out363), .data_out364(_add_all_x_data_out364), .data_out365(_add_all_x_data_out365), .data_out366(_add_all_x_data_out366), .data_out367(_add_all_x_data_out367), .data_out368(_add_all_x_data_out368), .data_out369(_add_all_x_data_out369), .data_out370(_add_all_x_data_out370), .data_out371(_add_all_x_data_out371), .data_out372(_add_all_x_data_out372), .data_out373(_add_all_x_data_out373), .data_out374(_add_all_x_data_out374), .data_out375(_add_all_x_data_out375), .data_out376(_add_all_x_data_out376), .data_out377(_add_all_x_data_out377), .data_out378(_add_all_x_data_out378), .data_out379(_add_all_x_data_out379), .data_out380(_add_all_x_data_out380), .data_out381(_add_all_x_data_out381), .data_out382(_add_all_x_data_out382), .data_out385(_add_all_x_data_out385), .data_out386(_add_all_x_data_out386), .data_out387(_add_all_x_data_out387), .data_out388(_add_all_x_data_out388), .data_out389(_add_all_x_data_out389), .data_out390(_add_all_x_data_out390), .data_out391(_add_all_x_data_out391), .data_out392(_add_all_x_data_out392), .data_out393(_add_all_x_data_out393), .data_out394(_add_all_x_data_out394), .data_out395(_add_all_x_data_out395), .data_out396(_add_all_x_data_out396), .data_out397(_add_all_x_data_out397), .data_out398(_add_all_x_data_out398), .data_out399(_add_all_x_data_out399), .data_out400(_add_all_x_data_out400), .data_out401(_add_all_x_data_out401), .data_out402(_add_all_x_data_out402), .data_out403(_add_all_x_data_out403), .data_out404(_add_all_x_data_out404), .data_out405(_add_all_x_data_out405), .data_out406(_add_all_x_data_out406), .data_out407(_add_all_x_data_out407), .data_out408(_add_all_x_data_out408), .data_out409(_add_all_x_data_out409), .data_out410(_add_all_x_data_out410), .data_out411(_add_all_x_data_out411), .data_out412(_add_all_x_data_out412), .data_out413(_add_all_x_data_out413), .data_out414(_add_all_x_data_out414), .data_out417(_add_all_x_data_out417), .data_out418(_add_all_x_data_out418), .data_out419(_add_all_x_data_out419), .data_out420(_add_all_x_data_out420), .data_out421(_add_all_x_data_out421), .data_out422(_add_all_x_data_out422), .data_out423(_add_all_x_data_out423), .data_out424(_add_all_x_data_out424), .data_out425(_add_all_x_data_out425), .data_out426(_add_all_x_data_out426), .data_out427(_add_all_x_data_out427), .data_out428(_add_all_x_data_out428), .data_out429(_add_all_x_data_out429), .data_out430(_add_all_x_data_out430), .data_out431(_add_all_x_data_out431), .data_out432(_add_all_x_data_out432), .data_out433(_add_all_x_data_out433), .data_out434(_add_all_x_data_out434), .data_out435(_add_all_x_data_out435), .data_out436(_add_all_x_data_out436), .data_out437(_add_all_x_data_out437), .data_out438(_add_all_x_data_out438), .data_out439(_add_all_x_data_out439), .data_out440(_add_all_x_data_out440), .data_out441(_add_all_x_data_out441), .data_out442(_add_all_x_data_out442), .data_out443(_add_all_x_data_out443), .data_out444(_add_all_x_data_out444), .data_out445(_add_all_x_data_out445), .data_out446(_add_all_x_data_out446), .data_out449(_add_all_x_data_out449), .data_out450(_add_all_x_data_out450), .data_out451(_add_all_x_data_out451), .data_out452(_add_all_x_data_out452), .data_out453(_add_all_x_data_out453), .data_out454(_add_all_x_data_out454), .data_out455(_add_all_x_data_out455), .data_out456(_add_all_x_data_out456), .data_out457(_add_all_x_data_out457), .data_out458(_add_all_x_data_out458), .data_out459(_add_all_x_data_out459), .data_out460(_add_all_x_data_out460), .data_out461(_add_all_x_data_out461), .data_out462(_add_all_x_data_out462), .data_out463(_add_all_x_data_out463), .data_out464(_add_all_x_data_out464), .data_out465(_add_all_x_data_out465), .data_out466(_add_all_x_data_out466), .data_out467(_add_all_x_data_out467), .data_out468(_add_all_x_data_out468), .data_out469(_add_all_x_data_out469), .data_out470(_add_all_x_data_out470), .data_out471(_add_all_x_data_out471), .data_out472(_add_all_x_data_out472), .data_out473(_add_all_x_data_out473), .data_out474(_add_all_x_data_out474), .data_out475(_add_all_x_data_out475), .data_out476(_add_all_x_data_out476), .data_out477(_add_all_x_data_out477), .data_out478(_add_all_x_data_out478), .data_in_org33(_add_all_x_data_in_org33), .data_in_org34(_add_all_x_data_in_org34), .data_in_org35(_add_all_x_data_in_org35), .data_in_org36(_add_all_x_data_in_org36), .data_in_org37(_add_all_x_data_in_org37), .data_in_org38(_add_all_x_data_in_org38), .data_in_org39(_add_all_x_data_in_org39), .data_in_org40(_add_all_x_data_in_org40), .data_in_org41(_add_all_x_data_in_org41), .data_in_org42(_add_all_x_data_in_org42), .data_in_org43(_add_all_x_data_in_org43), .data_in_org44(_add_all_x_data_in_org44), .data_in_org45(_add_all_x_data_in_org45), .data_in_org46(_add_all_x_data_in_org46), .data_in_org47(_add_all_x_data_in_org47), .data_in_org48(_add_all_x_data_in_org48), .data_in_org49(_add_all_x_data_in_org49), .data_in_org50(_add_all_x_data_in_org50), .data_in_org51(_add_all_x_data_in_org51), .data_in_org52(_add_all_x_data_in_org52), .data_in_org53(_add_all_x_data_in_org53), .data_in_org54(_add_all_x_data_in_org54), .data_in_org55(_add_all_x_data_in_org55), .data_in_org56(_add_all_x_data_in_org56), .data_in_org57(_add_all_x_data_in_org57), .data_in_org58(_add_all_x_data_in_org58), .data_in_org59(_add_all_x_data_in_org59), .data_in_org60(_add_all_x_data_in_org60), .data_in_org61(_add_all_x_data_in_org61), .data_in_org62(_add_all_x_data_in_org62), .data_in_org65(_add_all_x_data_in_org65), .data_in_org66(_add_all_x_data_in_org66), .data_in_org67(_add_all_x_data_in_org67), .data_in_org68(_add_all_x_data_in_org68), .data_in_org69(_add_all_x_data_in_org69), .data_in_org70(_add_all_x_data_in_org70), .data_in_org71(_add_all_x_data_in_org71), .data_in_org72(_add_all_x_data_in_org72), .data_in_org73(_add_all_x_data_in_org73), .data_in_org74(_add_all_x_data_in_org74), .data_in_org75(_add_all_x_data_in_org75), .data_in_org76(_add_all_x_data_in_org76), .data_in_org77(_add_all_x_data_in_org77), .data_in_org78(_add_all_x_data_in_org78), .data_in_org79(_add_all_x_data_in_org79), .data_in_org80(_add_all_x_data_in_org80), .data_in_org81(_add_all_x_data_in_org81), .data_in_org82(_add_all_x_data_in_org82), .data_in_org83(_add_all_x_data_in_org83), .data_in_org84(_add_all_x_data_in_org84), .data_in_org85(_add_all_x_data_in_org85), .data_in_org86(_add_all_x_data_in_org86), .data_in_org87(_add_all_x_data_in_org87), .data_in_org88(_add_all_x_data_in_org88), .data_in_org89(_add_all_x_data_in_org89), .data_in_org90(_add_all_x_data_in_org90), .data_in_org91(_add_all_x_data_in_org91), .data_in_org92(_add_all_x_data_in_org92), .data_in_org93(_add_all_x_data_in_org93), .data_in_org94(_add_all_x_data_in_org94), .data_in_org97(_add_all_x_data_in_org97), .data_in_org98(_add_all_x_data_in_org98), .data_in_org99(_add_all_x_data_in_org99), .data_in_org100(_add_all_x_data_in_org100), .data_in_org101(_add_all_x_data_in_org101), .data_in_org102(_add_all_x_data_in_org102), .data_in_org103(_add_all_x_data_in_org103), .data_in_org104(_add_all_x_data_in_org104), .data_in_org105(_add_all_x_data_in_org105), .data_in_org106(_add_all_x_data_in_org106), .data_in_org107(_add_all_x_data_in_org107), .data_in_org108(_add_all_x_data_in_org108), .data_in_org109(_add_all_x_data_in_org109), .data_in_org110(_add_all_x_data_in_org110), .data_in_org111(_add_all_x_data_in_org111), .data_in_org112(_add_all_x_data_in_org112), .data_in_org113(_add_all_x_data_in_org113), .data_in_org114(_add_all_x_data_in_org114), .data_in_org115(_add_all_x_data_in_org115), .data_in_org116(_add_all_x_data_in_org116), .data_in_org117(_add_all_x_data_in_org117), .data_in_org118(_add_all_x_data_in_org118), .data_in_org119(_add_all_x_data_in_org119), .data_in_org120(_add_all_x_data_in_org120), .data_in_org121(_add_all_x_data_in_org121), .data_in_org122(_add_all_x_data_in_org122), .data_in_org123(_add_all_x_data_in_org123), .data_in_org124(_add_all_x_data_in_org124), .data_in_org125(_add_all_x_data_in_org125), .data_in_org126(_add_all_x_data_in_org126), .data_in_org129(_add_all_x_data_in_org129), .data_in_org130(_add_all_x_data_in_org130), .data_in_org131(_add_all_x_data_in_org131), .data_in_org132(_add_all_x_data_in_org132), .data_in_org133(_add_all_x_data_in_org133), .data_in_org134(_add_all_x_data_in_org134), .data_in_org135(_add_all_x_data_in_org135), .data_in_org136(_add_all_x_data_in_org136), .data_in_org137(_add_all_x_data_in_org137), .data_in_org138(_add_all_x_data_in_org138), .data_in_org139(_add_all_x_data_in_org139), .data_in_org140(_add_all_x_data_in_org140), .data_in_org141(_add_all_x_data_in_org141), .data_in_org142(_add_all_x_data_in_org142), .data_in_org143(_add_all_x_data_in_org143), .data_in_org144(_add_all_x_data_in_org144), .data_in_org145(_add_all_x_data_in_org145), .data_in_org146(_add_all_x_data_in_org146), .data_in_org147(_add_all_x_data_in_org147), .data_in_org148(_add_all_x_data_in_org148), .data_in_org149(_add_all_x_data_in_org149), .data_in_org150(_add_all_x_data_in_org150), .data_in_org151(_add_all_x_data_in_org151), .data_in_org152(_add_all_x_data_in_org152), .data_in_org153(_add_all_x_data_in_org153), .data_in_org154(_add_all_x_data_in_org154), .data_in_org155(_add_all_x_data_in_org155), .data_in_org156(_add_all_x_data_in_org156), .data_in_org157(_add_all_x_data_in_org157), .data_in_org158(_add_all_x_data_in_org158), .data_in_org161(_add_all_x_data_in_org161), .data_in_org162(_add_all_x_data_in_org162), .data_in_org163(_add_all_x_data_in_org163), .data_in_org164(_add_all_x_data_in_org164), .data_in_org165(_add_all_x_data_in_org165), .data_in_org166(_add_all_x_data_in_org166), .data_in_org167(_add_all_x_data_in_org167), .data_in_org168(_add_all_x_data_in_org168), .data_in_org169(_add_all_x_data_in_org169), .data_in_org170(_add_all_x_data_in_org170), .data_in_org171(_add_all_x_data_in_org171), .data_in_org172(_add_all_x_data_in_org172), .data_in_org173(_add_all_x_data_in_org173), .data_in_org174(_add_all_x_data_in_org174), .data_in_org175(_add_all_x_data_in_org175), .data_in_org176(_add_all_x_data_in_org176), .data_in_org177(_add_all_x_data_in_org177), .data_in_org178(_add_all_x_data_in_org178), .data_in_org179(_add_all_x_data_in_org179), .data_in_org180(_add_all_x_data_in_org180), .data_in_org181(_add_all_x_data_in_org181), .data_in_org182(_add_all_x_data_in_org182), .data_in_org183(_add_all_x_data_in_org183), .data_in_org184(_add_all_x_data_in_org184), .data_in_org185(_add_all_x_data_in_org185), .data_in_org186(_add_all_x_data_in_org186), .data_in_org187(_add_all_x_data_in_org187), .data_in_org188(_add_all_x_data_in_org188), .data_in_org189(_add_all_x_data_in_org189), .data_in_org190(_add_all_x_data_in_org190), .data_in_org193(_add_all_x_data_in_org193), .data_in_org194(_add_all_x_data_in_org194), .data_in_org195(_add_all_x_data_in_org195), .data_in_org196(_add_all_x_data_in_org196), .data_in_org197(_add_all_x_data_in_org197), .data_in_org198(_add_all_x_data_in_org198), .data_in_org199(_add_all_x_data_in_org199), .data_in_org200(_add_all_x_data_in_org200), .data_in_org201(_add_all_x_data_in_org201), .data_in_org202(_add_all_x_data_in_org202), .data_in_org203(_add_all_x_data_in_org203), .data_in_org204(_add_all_x_data_in_org204), .data_in_org205(_add_all_x_data_in_org205), .data_in_org206(_add_all_x_data_in_org206), .data_in_org207(_add_all_x_data_in_org207), .data_in_org208(_add_all_x_data_in_org208), .data_in_org209(_add_all_x_data_in_org209), .data_in_org210(_add_all_x_data_in_org210), .data_in_org211(_add_all_x_data_in_org211), .data_in_org212(_add_all_x_data_in_org212), .data_in_org213(_add_all_x_data_in_org213), .data_in_org214(_add_all_x_data_in_org214), .data_in_org215(_add_all_x_data_in_org215), .data_in_org216(_add_all_x_data_in_org216), .data_in_org217(_add_all_x_data_in_org217), .data_in_org218(_add_all_x_data_in_org218), .data_in_org219(_add_all_x_data_in_org219), .data_in_org220(_add_all_x_data_in_org220), .data_in_org221(_add_all_x_data_in_org221), .data_in_org222(_add_all_x_data_in_org222), .data_in_org225(_add_all_x_data_in_org225), .data_in_org226(_add_all_x_data_in_org226), .data_in_org227(_add_all_x_data_in_org227), .data_in_org228(_add_all_x_data_in_org228), .data_in_org229(_add_all_x_data_in_org229), .data_in_org230(_add_all_x_data_in_org230), .data_in_org231(_add_all_x_data_in_org231), .data_in_org232(_add_all_x_data_in_org232), .data_in_org233(_add_all_x_data_in_org233), .data_in_org234(_add_all_x_data_in_org234), .data_in_org235(_add_all_x_data_in_org235), .data_in_org236(_add_all_x_data_in_org236), .data_in_org237(_add_all_x_data_in_org237), .data_in_org238(_add_all_x_data_in_org238), .data_in_org239(_add_all_x_data_in_org239), .data_in_org240(_add_all_x_data_in_org240), .data_in_org241(_add_all_x_data_in_org241), .data_in_org242(_add_all_x_data_in_org242), .data_in_org243(_add_all_x_data_in_org243), .data_in_org244(_add_all_x_data_in_org244), .data_in_org245(_add_all_x_data_in_org245), .data_in_org246(_add_all_x_data_in_org246), .data_in_org247(_add_all_x_data_in_org247), .data_in_org248(_add_all_x_data_in_org248), .data_in_org249(_add_all_x_data_in_org249), .data_in_org250(_add_all_x_data_in_org250), .data_in_org251(_add_all_x_data_in_org251), .data_in_org252(_add_all_x_data_in_org252), .data_in_org253(_add_all_x_data_in_org253), .data_in_org254(_add_all_x_data_in_org254), .data_in_org257(_add_all_x_data_in_org257), .data_in_org258(_add_all_x_data_in_org258), .data_in_org259(_add_all_x_data_in_org259), .data_in_org260(_add_all_x_data_in_org260), .data_in_org261(_add_all_x_data_in_org261), .data_in_org262(_add_all_x_data_in_org262), .data_in_org263(_add_all_x_data_in_org263), .data_in_org264(_add_all_x_data_in_org264), .data_in_org265(_add_all_x_data_in_org265), .data_in_org266(_add_all_x_data_in_org266), .data_in_org267(_add_all_x_data_in_org267), .data_in_org268(_add_all_x_data_in_org268), .data_in_org269(_add_all_x_data_in_org269), .data_in_org270(_add_all_x_data_in_org270), .data_in_org271(_add_all_x_data_in_org271), .data_in_org272(_add_all_x_data_in_org272), .data_in_org273(_add_all_x_data_in_org273), .data_in_org274(_add_all_x_data_in_org274), .data_in_org275(_add_all_x_data_in_org275), .data_in_org276(_add_all_x_data_in_org276), .data_in_org277(_add_all_x_data_in_org277), .data_in_org278(_add_all_x_data_in_org278), .data_in_org279(_add_all_x_data_in_org279), .data_in_org280(_add_all_x_data_in_org280), .data_in_org281(_add_all_x_data_in_org281), .data_in_org282(_add_all_x_data_in_org282), .data_in_org283(_add_all_x_data_in_org283), .data_in_org284(_add_all_x_data_in_org284), .data_in_org285(_add_all_x_data_in_org285), .data_in_org286(_add_all_x_data_in_org286), .data_in_org289(_add_all_x_data_in_org289), .data_in_org290(_add_all_x_data_in_org290), .data_in_org291(_add_all_x_data_in_org291), .data_in_org292(_add_all_x_data_in_org292), .data_in_org293(_add_all_x_data_in_org293), .data_in_org294(_add_all_x_data_in_org294), .data_in_org295(_add_all_x_data_in_org295), .data_in_org296(_add_all_x_data_in_org296), .data_in_org297(_add_all_x_data_in_org297), .data_in_org298(_add_all_x_data_in_org298), .data_in_org299(_add_all_x_data_in_org299), .data_in_org300(_add_all_x_data_in_org300), .data_in_org301(_add_all_x_data_in_org301), .data_in_org302(_add_all_x_data_in_org302), .data_in_org303(_add_all_x_data_in_org303), .data_in_org304(_add_all_x_data_in_org304), .data_in_org305(_add_all_x_data_in_org305), .data_in_org306(_add_all_x_data_in_org306), .data_in_org307(_add_all_x_data_in_org307), .data_in_org308(_add_all_x_data_in_org308), .data_in_org309(_add_all_x_data_in_org309), .data_in_org310(_add_all_x_data_in_org310), .data_in_org311(_add_all_x_data_in_org311), .data_in_org312(_add_all_x_data_in_org312), .data_in_org313(_add_all_x_data_in_org313), .data_in_org314(_add_all_x_data_in_org314), .data_in_org315(_add_all_x_data_in_org315), .data_in_org316(_add_all_x_data_in_org316), .data_in_org317(_add_all_x_data_in_org317), .data_in_org318(_add_all_x_data_in_org318), .data_in_org321(_add_all_x_data_in_org321), .data_in_org322(_add_all_x_data_in_org322), .data_in_org323(_add_all_x_data_in_org323), .data_in_org324(_add_all_x_data_in_org324), .data_in_org325(_add_all_x_data_in_org325), .data_in_org326(_add_all_x_data_in_org326), .data_in_org327(_add_all_x_data_in_org327), .data_in_org328(_add_all_x_data_in_org328), .data_in_org329(_add_all_x_data_in_org329), .data_in_org330(_add_all_x_data_in_org330), .data_in_org331(_add_all_x_data_in_org331), .data_in_org332(_add_all_x_data_in_org332), .data_in_org333(_add_all_x_data_in_org333), .data_in_org334(_add_all_x_data_in_org334), .data_in_org335(_add_all_x_data_in_org335), .data_in_org336(_add_all_x_data_in_org336), .data_in_org337(_add_all_x_data_in_org337), .data_in_org338(_add_all_x_data_in_org338), .data_in_org339(_add_all_x_data_in_org339), .data_in_org340(_add_all_x_data_in_org340), .data_in_org341(_add_all_x_data_in_org341), .data_in_org342(_add_all_x_data_in_org342), .data_in_org343(_add_all_x_data_in_org343), .data_in_org344(_add_all_x_data_in_org344), .data_in_org345(_add_all_x_data_in_org345), .data_in_org346(_add_all_x_data_in_org346), .data_in_org347(_add_all_x_data_in_org347), .data_in_org348(_add_all_x_data_in_org348), .data_in_org349(_add_all_x_data_in_org349), .data_in_org350(_add_all_x_data_in_org350), .data_in_org353(_add_all_x_data_in_org353), .data_in_org354(_add_all_x_data_in_org354), .data_in_org355(_add_all_x_data_in_org355), .data_in_org356(_add_all_x_data_in_org356), .data_in_org357(_add_all_x_data_in_org357), .data_in_org358(_add_all_x_data_in_org358), .data_in_org359(_add_all_x_data_in_org359), .data_in_org360(_add_all_x_data_in_org360), .data_in_org361(_add_all_x_data_in_org361), .data_in_org362(_add_all_x_data_in_org362), .data_in_org363(_add_all_x_data_in_org363), .data_in_org364(_add_all_x_data_in_org364), .data_in_org365(_add_all_x_data_in_org365), .data_in_org366(_add_all_x_data_in_org366), .data_in_org367(_add_all_x_data_in_org367), .data_in_org368(_add_all_x_data_in_org368), .data_in_org369(_add_all_x_data_in_org369), .data_in_org370(_add_all_x_data_in_org370), .data_in_org371(_add_all_x_data_in_org371), .data_in_org372(_add_all_x_data_in_org372), .data_in_org373(_add_all_x_data_in_org373), .data_in_org374(_add_all_x_data_in_org374), .data_in_org375(_add_all_x_data_in_org375), .data_in_org376(_add_all_x_data_in_org376), .data_in_org377(_add_all_x_data_in_org377), .data_in_org378(_add_all_x_data_in_org378), .data_in_org379(_add_all_x_data_in_org379), .data_in_org380(_add_all_x_data_in_org380), .data_in_org381(_add_all_x_data_in_org381), .data_in_org382(_add_all_x_data_in_org382), .data_in_org385(_add_all_x_data_in_org385), .data_in_org386(_add_all_x_data_in_org386), .data_in_org387(_add_all_x_data_in_org387), .data_in_org388(_add_all_x_data_in_org388), .data_in_org389(_add_all_x_data_in_org389), .data_in_org390(_add_all_x_data_in_org390), .data_in_org391(_add_all_x_data_in_org391), .data_in_org392(_add_all_x_data_in_org392), .data_in_org393(_add_all_x_data_in_org393), .data_in_org394(_add_all_x_data_in_org394), .data_in_org395(_add_all_x_data_in_org395), .data_in_org396(_add_all_x_data_in_org396), .data_in_org397(_add_all_x_data_in_org397), .data_in_org398(_add_all_x_data_in_org398), .data_in_org399(_add_all_x_data_in_org399), .data_in_org400(_add_all_x_data_in_org400), .data_in_org401(_add_all_x_data_in_org401), .data_in_org402(_add_all_x_data_in_org402), .data_in_org403(_add_all_x_data_in_org403), .data_in_org404(_add_all_x_data_in_org404), .data_in_org405(_add_all_x_data_in_org405), .data_in_org406(_add_all_x_data_in_org406), .data_in_org407(_add_all_x_data_in_org407), .data_in_org408(_add_all_x_data_in_org408), .data_in_org409(_add_all_x_data_in_org409), .data_in_org410(_add_all_x_data_in_org410), .data_in_org411(_add_all_x_data_in_org411), .data_in_org412(_add_all_x_data_in_org412), .data_in_org413(_add_all_x_data_in_org413), .data_in_org414(_add_all_x_data_in_org414), .data_in_org417(_add_all_x_data_in_org417), .data_in_org418(_add_all_x_data_in_org418), .data_in_org419(_add_all_x_data_in_org419), .data_in_org420(_add_all_x_data_in_org420), .data_in_org421(_add_all_x_data_in_org421), .data_in_org422(_add_all_x_data_in_org422), .data_in_org423(_add_all_x_data_in_org423), .data_in_org424(_add_all_x_data_in_org424), .data_in_org425(_add_all_x_data_in_org425), .data_in_org426(_add_all_x_data_in_org426), .data_in_org427(_add_all_x_data_in_org427), .data_in_org428(_add_all_x_data_in_org428), .data_in_org429(_add_all_x_data_in_org429), .data_in_org430(_add_all_x_data_in_org430), .data_in_org431(_add_all_x_data_in_org431), .data_in_org432(_add_all_x_data_in_org432), .data_in_org433(_add_all_x_data_in_org433), .data_in_org434(_add_all_x_data_in_org434), .data_in_org435(_add_all_x_data_in_org435), .data_in_org436(_add_all_x_data_in_org436), .data_in_org437(_add_all_x_data_in_org437), .data_in_org438(_add_all_x_data_in_org438), .data_in_org439(_add_all_x_data_in_org439), .data_in_org440(_add_all_x_data_in_org440), .data_in_org441(_add_all_x_data_in_org441), .data_in_org442(_add_all_x_data_in_org442), .data_in_org443(_add_all_x_data_in_org443), .data_in_org444(_add_all_x_data_in_org444), .data_in_org445(_add_all_x_data_in_org445), .data_in_org446(_add_all_x_data_in_org446), .data_in_org449(_add_all_x_data_in_org449), .data_in_org450(_add_all_x_data_in_org450), .data_in_org451(_add_all_x_data_in_org451), .data_in_org452(_add_all_x_data_in_org452), .data_in_org453(_add_all_x_data_in_org453), .data_in_org454(_add_all_x_data_in_org454), .data_in_org455(_add_all_x_data_in_org455), .data_in_org456(_add_all_x_data_in_org456), .data_in_org457(_add_all_x_data_in_org457), .data_in_org458(_add_all_x_data_in_org458), .data_in_org459(_add_all_x_data_in_org459), .data_in_org460(_add_all_x_data_in_org460), .data_in_org461(_add_all_x_data_in_org461), .data_in_org462(_add_all_x_data_in_org462), .data_in_org463(_add_all_x_data_in_org463), .data_in_org464(_add_all_x_data_in_org464), .data_in_org465(_add_all_x_data_in_org465), .data_in_org466(_add_all_x_data_in_org466), .data_in_org467(_add_all_x_data_in_org467), .data_in_org468(_add_all_x_data_in_org468), .data_in_org469(_add_all_x_data_in_org469), .data_in_org470(_add_all_x_data_in_org470), .data_in_org471(_add_all_x_data_in_org471), .data_in_org472(_add_all_x_data_in_org472), .data_in_org473(_add_all_x_data_in_org473), .data_in_org474(_add_all_x_data_in_org474), .data_in_org475(_add_all_x_data_in_org475), .data_in_org476(_add_all_x_data_in_org476), .data_in_org477(_add_all_x_data_in_org477), .data_in_org478(_add_all_x_data_in_org478), .data_out_org33(_add_all_x_data_out_org33), .data_out_org34(_add_all_x_data_out_org34), .data_out_org35(_add_all_x_data_out_org35), .data_out_org36(_add_all_x_data_out_org36), .data_out_org37(_add_all_x_data_out_org37), .data_out_org38(_add_all_x_data_out_org38), .data_out_org39(_add_all_x_data_out_org39), .data_out_org40(_add_all_x_data_out_org40), .data_out_org41(_add_all_x_data_out_org41), .data_out_org42(_add_all_x_data_out_org42), .data_out_org43(_add_all_x_data_out_org43), .data_out_org44(_add_all_x_data_out_org44), .data_out_org45(_add_all_x_data_out_org45), .data_out_org46(_add_all_x_data_out_org46), .data_out_org47(_add_all_x_data_out_org47), .data_out_org48(_add_all_x_data_out_org48), .data_out_org49(_add_all_x_data_out_org49), .data_out_org50(_add_all_x_data_out_org50), .data_out_org51(_add_all_x_data_out_org51), .data_out_org52(_add_all_x_data_out_org52), .data_out_org53(_add_all_x_data_out_org53), .data_out_org54(_add_all_x_data_out_org54), .data_out_org55(_add_all_x_data_out_org55), .data_out_org56(_add_all_x_data_out_org56), .data_out_org57(_add_all_x_data_out_org57), .data_out_org58(_add_all_x_data_out_org58), .data_out_org59(_add_all_x_data_out_org59), .data_out_org60(_add_all_x_data_out_org60), .data_out_org61(_add_all_x_data_out_org61), .data_out_org62(_add_all_x_data_out_org62), .data_out_org65(_add_all_x_data_out_org65), .data_out_org66(_add_all_x_data_out_org66), .data_out_org67(_add_all_x_data_out_org67), .data_out_org68(_add_all_x_data_out_org68), .data_out_org69(_add_all_x_data_out_org69), .data_out_org70(_add_all_x_data_out_org70), .data_out_org71(_add_all_x_data_out_org71), .data_out_org72(_add_all_x_data_out_org72), .data_out_org73(_add_all_x_data_out_org73), .data_out_org74(_add_all_x_data_out_org74), .data_out_org75(_add_all_x_data_out_org75), .data_out_org76(_add_all_x_data_out_org76), .data_out_org77(_add_all_x_data_out_org77), .data_out_org78(_add_all_x_data_out_org78), .data_out_org79(_add_all_x_data_out_org79), .data_out_org80(_add_all_x_data_out_org80), .data_out_org81(_add_all_x_data_out_org81), .data_out_org82(_add_all_x_data_out_org82), .data_out_org83(_add_all_x_data_out_org83), .data_out_org84(_add_all_x_data_out_org84), .data_out_org85(_add_all_x_data_out_org85), .data_out_org86(_add_all_x_data_out_org86), .data_out_org87(_add_all_x_data_out_org87), .data_out_org88(_add_all_x_data_out_org88), .data_out_org89(_add_all_x_data_out_org89), .data_out_org90(_add_all_x_data_out_org90), .data_out_org91(_add_all_x_data_out_org91), .data_out_org92(_add_all_x_data_out_org92), .data_out_org93(_add_all_x_data_out_org93), .data_out_org94(_add_all_x_data_out_org94), .data_out_org97(_add_all_x_data_out_org97), .data_out_org98(_add_all_x_data_out_org98), .data_out_org99(_add_all_x_data_out_org99), .data_out_org100(_add_all_x_data_out_org100), .data_out_org101(_add_all_x_data_out_org101), .data_out_org102(_add_all_x_data_out_org102), .data_out_org103(_add_all_x_data_out_org103), .data_out_org104(_add_all_x_data_out_org104), .data_out_org105(_add_all_x_data_out_org105), .data_out_org106(_add_all_x_data_out_org106), .data_out_org107(_add_all_x_data_out_org107), .data_out_org108(_add_all_x_data_out_org108), .data_out_org109(_add_all_x_data_out_org109), .data_out_org110(_add_all_x_data_out_org110), .data_out_org111(_add_all_x_data_out_org111), .data_out_org112(_add_all_x_data_out_org112), .data_out_org113(_add_all_x_data_out_org113), .data_out_org114(_add_all_x_data_out_org114), .data_out_org115(_add_all_x_data_out_org115), .data_out_org116(_add_all_x_data_out_org116), .data_out_org117(_add_all_x_data_out_org117), .data_out_org118(_add_all_x_data_out_org118), .data_out_org119(_add_all_x_data_out_org119), .data_out_org120(_add_all_x_data_out_org120), .data_out_org121(_add_all_x_data_out_org121), .data_out_org122(_add_all_x_data_out_org122), .data_out_org123(_add_all_x_data_out_org123), .data_out_org124(_add_all_x_data_out_org124), .data_out_org125(_add_all_x_data_out_org125), .data_out_org126(_add_all_x_data_out_org126), .data_out_org129(_add_all_x_data_out_org129), .data_out_org130(_add_all_x_data_out_org130), .data_out_org131(_add_all_x_data_out_org131), .data_out_org132(_add_all_x_data_out_org132), .data_out_org133(_add_all_x_data_out_org133), .data_out_org134(_add_all_x_data_out_org134), .data_out_org135(_add_all_x_data_out_org135), .data_out_org136(_add_all_x_data_out_org136), .data_out_org137(_add_all_x_data_out_org137), .data_out_org138(_add_all_x_data_out_org138), .data_out_org139(_add_all_x_data_out_org139), .data_out_org140(_add_all_x_data_out_org140), .data_out_org141(_add_all_x_data_out_org141), .data_out_org142(_add_all_x_data_out_org142), .data_out_org143(_add_all_x_data_out_org143), .data_out_org144(_add_all_x_data_out_org144), .data_out_org145(_add_all_x_data_out_org145), .data_out_org146(_add_all_x_data_out_org146), .data_out_org147(_add_all_x_data_out_org147), .data_out_org148(_add_all_x_data_out_org148), .data_out_org149(_add_all_x_data_out_org149), .data_out_org150(_add_all_x_data_out_org150), .data_out_org151(_add_all_x_data_out_org151), .data_out_org152(_add_all_x_data_out_org152), .data_out_org153(_add_all_x_data_out_org153), .data_out_org154(_add_all_x_data_out_org154), .data_out_org155(_add_all_x_data_out_org155), .data_out_org156(_add_all_x_data_out_org156), .data_out_org157(_add_all_x_data_out_org157), .data_out_org158(_add_all_x_data_out_org158), .data_out_org161(_add_all_x_data_out_org161), .data_out_org162(_add_all_x_data_out_org162), .data_out_org163(_add_all_x_data_out_org163), .data_out_org164(_add_all_x_data_out_org164), .data_out_org165(_add_all_x_data_out_org165), .data_out_org166(_add_all_x_data_out_org166), .data_out_org167(_add_all_x_data_out_org167), .data_out_org168(_add_all_x_data_out_org168), .data_out_org169(_add_all_x_data_out_org169), .data_out_org170(_add_all_x_data_out_org170), .data_out_org171(_add_all_x_data_out_org171), .data_out_org172(_add_all_x_data_out_org172), .data_out_org173(_add_all_x_data_out_org173), .data_out_org174(_add_all_x_data_out_org174), .data_out_org175(_add_all_x_data_out_org175), .data_out_org176(_add_all_x_data_out_org176), .data_out_org177(_add_all_x_data_out_org177), .data_out_org178(_add_all_x_data_out_org178), .data_out_org179(_add_all_x_data_out_org179), .data_out_org180(_add_all_x_data_out_org180), .data_out_org181(_add_all_x_data_out_org181), .data_out_org182(_add_all_x_data_out_org182), .data_out_org183(_add_all_x_data_out_org183), .data_out_org184(_add_all_x_data_out_org184), .data_out_org185(_add_all_x_data_out_org185), .data_out_org186(_add_all_x_data_out_org186), .data_out_org187(_add_all_x_data_out_org187), .data_out_org188(_add_all_x_data_out_org188), .data_out_org189(_add_all_x_data_out_org189), .data_out_org190(_add_all_x_data_out_org190), .data_out_org193(_add_all_x_data_out_org193), .data_out_org194(_add_all_x_data_out_org194), .data_out_org195(_add_all_x_data_out_org195), .data_out_org196(_add_all_x_data_out_org196), .data_out_org197(_add_all_x_data_out_org197), .data_out_org198(_add_all_x_data_out_org198), .data_out_org199(_add_all_x_data_out_org199), .data_out_org200(_add_all_x_data_out_org200), .data_out_org201(_add_all_x_data_out_org201), .data_out_org202(_add_all_x_data_out_org202), .data_out_org203(_add_all_x_data_out_org203), .data_out_org204(_add_all_x_data_out_org204), .data_out_org205(_add_all_x_data_out_org205), .data_out_org206(_add_all_x_data_out_org206), .data_out_org207(_add_all_x_data_out_org207), .data_out_org208(_add_all_x_data_out_org208), .data_out_org209(_add_all_x_data_out_org209), .data_out_org210(_add_all_x_data_out_org210), .data_out_org211(_add_all_x_data_out_org211), .data_out_org212(_add_all_x_data_out_org212), .data_out_org213(_add_all_x_data_out_org213), .data_out_org214(_add_all_x_data_out_org214), .data_out_org215(_add_all_x_data_out_org215), .data_out_org216(_add_all_x_data_out_org216), .data_out_org217(_add_all_x_data_out_org217), .data_out_org218(_add_all_x_data_out_org218), .data_out_org219(_add_all_x_data_out_org219), .data_out_org220(_add_all_x_data_out_org220), .data_out_org221(_add_all_x_data_out_org221), .data_out_org222(_add_all_x_data_out_org222), .data_out_org225(_add_all_x_data_out_org225), .data_out_org226(_add_all_x_data_out_org226), .data_out_org227(_add_all_x_data_out_org227), .data_out_org228(_add_all_x_data_out_org228), .data_out_org229(_add_all_x_data_out_org229), .data_out_org230(_add_all_x_data_out_org230), .data_out_org231(_add_all_x_data_out_org231), .data_out_org232(_add_all_x_data_out_org232), .data_out_org233(_add_all_x_data_out_org233), .data_out_org234(_add_all_x_data_out_org234), .data_out_org235(_add_all_x_data_out_org235), .data_out_org236(_add_all_x_data_out_org236), .data_out_org237(_add_all_x_data_out_org237), .data_out_org238(_add_all_x_data_out_org238), .data_out_org239(_add_all_x_data_out_org239), .data_out_org240(_add_all_x_data_out_org240), .data_out_org241(_add_all_x_data_out_org241), .data_out_org242(_add_all_x_data_out_org242), .data_out_org243(_add_all_x_data_out_org243), .data_out_org244(_add_all_x_data_out_org244), .data_out_org245(_add_all_x_data_out_org245), .data_out_org246(_add_all_x_data_out_org246), .data_out_org247(_add_all_x_data_out_org247), .data_out_org248(_add_all_x_data_out_org248), .data_out_org249(_add_all_x_data_out_org249), .data_out_org250(_add_all_x_data_out_org250), .data_out_org251(_add_all_x_data_out_org251), .data_out_org252(_add_all_x_data_out_org252), .data_out_org253(_add_all_x_data_out_org253), .data_out_org254(_add_all_x_data_out_org254), .data_out_org257(_add_all_x_data_out_org257), .data_out_org258(_add_all_x_data_out_org258), .data_out_org259(_add_all_x_data_out_org259), .data_out_org260(_add_all_x_data_out_org260), .data_out_org261(_add_all_x_data_out_org261), .data_out_org262(_add_all_x_data_out_org262), .data_out_org263(_add_all_x_data_out_org263), .data_out_org264(_add_all_x_data_out_org264), .data_out_org265(_add_all_x_data_out_org265), .data_out_org266(_add_all_x_data_out_org266), .data_out_org267(_add_all_x_data_out_org267), .data_out_org268(_add_all_x_data_out_org268), .data_out_org269(_add_all_x_data_out_org269), .data_out_org270(_add_all_x_data_out_org270), .data_out_org271(_add_all_x_data_out_org271), .data_out_org272(_add_all_x_data_out_org272), .data_out_org273(_add_all_x_data_out_org273), .data_out_org274(_add_all_x_data_out_org274), .data_out_org275(_add_all_x_data_out_org275), .data_out_org276(_add_all_x_data_out_org276), .data_out_org277(_add_all_x_data_out_org277), .data_out_org278(_add_all_x_data_out_org278), .data_out_org279(_add_all_x_data_out_org279), .data_out_org280(_add_all_x_data_out_org280), .data_out_org281(_add_all_x_data_out_org281), .data_out_org282(_add_all_x_data_out_org282), .data_out_org283(_add_all_x_data_out_org283), .data_out_org284(_add_all_x_data_out_org284), .data_out_org285(_add_all_x_data_out_org285), .data_out_org286(_add_all_x_data_out_org286), .data_out_org289(_add_all_x_data_out_org289), .data_out_org290(_add_all_x_data_out_org290), .data_out_org291(_add_all_x_data_out_org291), .data_out_org292(_add_all_x_data_out_org292), .data_out_org293(_add_all_x_data_out_org293), .data_out_org294(_add_all_x_data_out_org294), .data_out_org295(_add_all_x_data_out_org295), .data_out_org296(_add_all_x_data_out_org296), .data_out_org297(_add_all_x_data_out_org297), .data_out_org298(_add_all_x_data_out_org298), .data_out_org299(_add_all_x_data_out_org299), .data_out_org300(_add_all_x_data_out_org300), .data_out_org301(_add_all_x_data_out_org301), .data_out_org302(_add_all_x_data_out_org302), .data_out_org303(_add_all_x_data_out_org303), .data_out_org304(_add_all_x_data_out_org304), .data_out_org305(_add_all_x_data_out_org305), .data_out_org306(_add_all_x_data_out_org306), .data_out_org307(_add_all_x_data_out_org307), .data_out_org308(_add_all_x_data_out_org308), .data_out_org309(_add_all_x_data_out_org309), .data_out_org310(_add_all_x_data_out_org310), .data_out_org311(_add_all_x_data_out_org311), .data_out_org312(_add_all_x_data_out_org312), .data_out_org313(_add_all_x_data_out_org313), .data_out_org314(_add_all_x_data_out_org314), .data_out_org315(_add_all_x_data_out_org315), .data_out_org316(_add_all_x_data_out_org316), .data_out_org317(_add_all_x_data_out_org317), .data_out_org318(_add_all_x_data_out_org318), .data_out_org321(_add_all_x_data_out_org321), .data_out_org322(_add_all_x_data_out_org322), .data_out_org323(_add_all_x_data_out_org323), .data_out_org324(_add_all_x_data_out_org324), .data_out_org325(_add_all_x_data_out_org325), .data_out_org326(_add_all_x_data_out_org326), .data_out_org327(_add_all_x_data_out_org327), .data_out_org328(_add_all_x_data_out_org328), .data_out_org329(_add_all_x_data_out_org329), .data_out_org330(_add_all_x_data_out_org330), .data_out_org331(_add_all_x_data_out_org331), .data_out_org332(_add_all_x_data_out_org332), .data_out_org333(_add_all_x_data_out_org333), .data_out_org334(_add_all_x_data_out_org334), .data_out_org335(_add_all_x_data_out_org335), .data_out_org336(_add_all_x_data_out_org336), .data_out_org337(_add_all_x_data_out_org337), .data_out_org338(_add_all_x_data_out_org338), .data_out_org339(_add_all_x_data_out_org339), .data_out_org340(_add_all_x_data_out_org340), .data_out_org341(_add_all_x_data_out_org341), .data_out_org342(_add_all_x_data_out_org342), .data_out_org343(_add_all_x_data_out_org343), .data_out_org344(_add_all_x_data_out_org344), .data_out_org345(_add_all_x_data_out_org345), .data_out_org346(_add_all_x_data_out_org346), .data_out_org347(_add_all_x_data_out_org347), .data_out_org348(_add_all_x_data_out_org348), .data_out_org349(_add_all_x_data_out_org349), .data_out_org350(_add_all_x_data_out_org350), .data_out_org353(_add_all_x_data_out_org353), .data_out_org354(_add_all_x_data_out_org354), .data_out_org355(_add_all_x_data_out_org355), .data_out_org356(_add_all_x_data_out_org356), .data_out_org357(_add_all_x_data_out_org357), .data_out_org358(_add_all_x_data_out_org358), .data_out_org359(_add_all_x_data_out_org359), .data_out_org360(_add_all_x_data_out_org360), .data_out_org361(_add_all_x_data_out_org361), .data_out_org362(_add_all_x_data_out_org362), .data_out_org363(_add_all_x_data_out_org363), .data_out_org364(_add_all_x_data_out_org364), .data_out_org365(_add_all_x_data_out_org365), .data_out_org366(_add_all_x_data_out_org366), .data_out_org367(_add_all_x_data_out_org367), .data_out_org368(_add_all_x_data_out_org368), .data_out_org369(_add_all_x_data_out_org369), .data_out_org370(_add_all_x_data_out_org370), .data_out_org371(_add_all_x_data_out_org371), .data_out_org372(_add_all_x_data_out_org372), .data_out_org373(_add_all_x_data_out_org373), .data_out_org374(_add_all_x_data_out_org374), .data_out_org375(_add_all_x_data_out_org375), .data_out_org376(_add_all_x_data_out_org376), .data_out_org377(_add_all_x_data_out_org377), .data_out_org378(_add_all_x_data_out_org378), .data_out_org379(_add_all_x_data_out_org379), .data_out_org380(_add_all_x_data_out_org380), .data_out_org381(_add_all_x_data_out_org381), .data_out_org382(_add_all_x_data_out_org382), .data_out_org385(_add_all_x_data_out_org385), .data_out_org386(_add_all_x_data_out_org386), .data_out_org387(_add_all_x_data_out_org387), .data_out_org388(_add_all_x_data_out_org388), .data_out_org389(_add_all_x_data_out_org389), .data_out_org390(_add_all_x_data_out_org390), .data_out_org391(_add_all_x_data_out_org391), .data_out_org392(_add_all_x_data_out_org392), .data_out_org393(_add_all_x_data_out_org393), .data_out_org394(_add_all_x_data_out_org394), .data_out_org395(_add_all_x_data_out_org395), .data_out_org396(_add_all_x_data_out_org396), .data_out_org397(_add_all_x_data_out_org397), .data_out_org398(_add_all_x_data_out_org398), .data_out_org399(_add_all_x_data_out_org399), .data_out_org400(_add_all_x_data_out_org400), .data_out_org401(_add_all_x_data_out_org401), .data_out_org402(_add_all_x_data_out_org402), .data_out_org403(_add_all_x_data_out_org403), .data_out_org404(_add_all_x_data_out_org404), .data_out_org405(_add_all_x_data_out_org405), .data_out_org406(_add_all_x_data_out_org406), .data_out_org407(_add_all_x_data_out_org407), .data_out_org408(_add_all_x_data_out_org408), .data_out_org409(_add_all_x_data_out_org409), .data_out_org410(_add_all_x_data_out_org410), .data_out_org411(_add_all_x_data_out_org411), .data_out_org412(_add_all_x_data_out_org412), .data_out_org413(_add_all_x_data_out_org413), .data_out_org414(_add_all_x_data_out_org414), .data_out_org417(_add_all_x_data_out_org417), .data_out_org418(_add_all_x_data_out_org418), .data_out_org419(_add_all_x_data_out_org419), .data_out_org420(_add_all_x_data_out_org420), .data_out_org421(_add_all_x_data_out_org421), .data_out_org422(_add_all_x_data_out_org422), .data_out_org423(_add_all_x_data_out_org423), .data_out_org424(_add_all_x_data_out_org424), .data_out_org425(_add_all_x_data_out_org425), .data_out_org426(_add_all_x_data_out_org426), .data_out_org427(_add_all_x_data_out_org427), .data_out_org428(_add_all_x_data_out_org428), .data_out_org429(_add_all_x_data_out_org429), .data_out_org430(_add_all_x_data_out_org430), .data_out_org431(_add_all_x_data_out_org431), .data_out_org432(_add_all_x_data_out_org432), .data_out_org433(_add_all_x_data_out_org433), .data_out_org434(_add_all_x_data_out_org434), .data_out_org435(_add_all_x_data_out_org435), .data_out_org436(_add_all_x_data_out_org436), .data_out_org437(_add_all_x_data_out_org437), .data_out_org438(_add_all_x_data_out_org438), .data_out_org439(_add_all_x_data_out_org439), .data_out_org440(_add_all_x_data_out_org440), .data_out_org441(_add_all_x_data_out_org441), .data_out_org442(_add_all_x_data_out_org442), .data_out_org443(_add_all_x_data_out_org443), .data_out_org444(_add_all_x_data_out_org444), .data_out_org445(_add_all_x_data_out_org445), .data_out_org446(_add_all_x_data_out_org446), .data_out_org449(_add_all_x_data_out_org449), .data_out_org450(_add_all_x_data_out_org450), .data_out_org451(_add_all_x_data_out_org451), .data_out_org452(_add_all_x_data_out_org452), .data_out_org453(_add_all_x_data_out_org453), .data_out_org454(_add_all_x_data_out_org454), .data_out_org455(_add_all_x_data_out_org455), .data_out_org456(_add_all_x_data_out_org456), .data_out_org457(_add_all_x_data_out_org457), .data_out_org458(_add_all_x_data_out_org458), .data_out_org459(_add_all_x_data_out_org459), .data_out_org460(_add_all_x_data_out_org460), .data_out_org461(_add_all_x_data_out_org461), .data_out_org462(_add_all_x_data_out_org462), .data_out_org463(_add_all_x_data_out_org463), .data_out_org464(_add_all_x_data_out_org464), .data_out_org465(_add_all_x_data_out_org465), .data_out_org466(_add_all_x_data_out_org466), .data_out_org467(_add_all_x_data_out_org467), .data_out_org468(_add_all_x_data_out_org468), .data_out_org469(_add_all_x_data_out_org469), .data_out_org470(_add_all_x_data_out_org470), .data_out_org471(_add_all_x_data_out_org471), .data_out_org472(_add_all_x_data_out_org472), .data_out_org473(_add_all_x_data_out_org473), .data_out_org474(_add_all_x_data_out_org474), .data_out_org475(_add_all_x_data_out_org475), .data_out_org476(_add_all_x_data_out_org476), .data_out_org477(_add_all_x_data_out_org477), .data_out_org478(_add_all_x_data_out_org478), .data_in33(_add_all_x_data_in33), .data_in34(_add_all_x_data_in34), .data_in35(_add_all_x_data_in35), .data_in36(_add_all_x_data_in36), .data_in37(_add_all_x_data_in37), .data_in38(_add_all_x_data_in38), .data_in39(_add_all_x_data_in39), .data_in40(_add_all_x_data_in40), .data_in41(_add_all_x_data_in41), .data_in42(_add_all_x_data_in42), .data_in43(_add_all_x_data_in43), .data_in44(_add_all_x_data_in44), .data_in45(_add_all_x_data_in45), .data_in46(_add_all_x_data_in46), .data_in47(_add_all_x_data_in47), .data_in48(_add_all_x_data_in48), .data_in49(_add_all_x_data_in49), .data_in50(_add_all_x_data_in50), .data_in51(_add_all_x_data_in51), .data_in52(_add_all_x_data_in52), .data_in53(_add_all_x_data_in53), .data_in54(_add_all_x_data_in54), .data_in55(_add_all_x_data_in55), .data_in56(_add_all_x_data_in56), .data_in57(_add_all_x_data_in57), .data_in58(_add_all_x_data_in58), .data_in59(_add_all_x_data_in59), .data_in60(_add_all_x_data_in60), .data_in61(_add_all_x_data_in61), .data_in62(_add_all_x_data_in62), .data_in65(_add_all_x_data_in65), .data_in66(_add_all_x_data_in66), .data_in67(_add_all_x_data_in67), .data_in68(_add_all_x_data_in68), .data_in69(_add_all_x_data_in69), .data_in70(_add_all_x_data_in70), .data_in71(_add_all_x_data_in71), .data_in72(_add_all_x_data_in72), .data_in73(_add_all_x_data_in73), .data_in74(_add_all_x_data_in74), .data_in75(_add_all_x_data_in75), .data_in76(_add_all_x_data_in76), .data_in77(_add_all_x_data_in77), .data_in78(_add_all_x_data_in78), .data_in79(_add_all_x_data_in79), .data_in80(_add_all_x_data_in80), .data_in81(_add_all_x_data_in81), .data_in82(_add_all_x_data_in82), .data_in83(_add_all_x_data_in83), .data_in84(_add_all_x_data_in84), .data_in85(_add_all_x_data_in85), .data_in86(_add_all_x_data_in86), .data_in87(_add_all_x_data_in87), .data_in88(_add_all_x_data_in88), .data_in89(_add_all_x_data_in89), .data_in90(_add_all_x_data_in90), .data_in91(_add_all_x_data_in91), .data_in92(_add_all_x_data_in92), .data_in93(_add_all_x_data_in93), .data_in94(_add_all_x_data_in94), .data_in97(_add_all_x_data_in97), .data_in98(_add_all_x_data_in98), .data_in99(_add_all_x_data_in99), .data_in100(_add_all_x_data_in100), .data_in101(_add_all_x_data_in101), .data_in102(_add_all_x_data_in102), .data_in103(_add_all_x_data_in103), .data_in104(_add_all_x_data_in104), .data_in105(_add_all_x_data_in105), .data_in106(_add_all_x_data_in106), .data_in107(_add_all_x_data_in107), .data_in108(_add_all_x_data_in108), .data_in109(_add_all_x_data_in109), .data_in110(_add_all_x_data_in110), .data_in111(_add_all_x_data_in111), .data_in112(_add_all_x_data_in112), .data_in113(_add_all_x_data_in113), .data_in114(_add_all_x_data_in114), .data_in115(_add_all_x_data_in115), .data_in116(_add_all_x_data_in116), .data_in117(_add_all_x_data_in117), .data_in118(_add_all_x_data_in118), .data_in119(_add_all_x_data_in119), .data_in120(_add_all_x_data_in120), .data_in121(_add_all_x_data_in121), .data_in122(_add_all_x_data_in122), .data_in123(_add_all_x_data_in123), .data_in124(_add_all_x_data_in124), .data_in125(_add_all_x_data_in125), .data_in126(_add_all_x_data_in126), .data_in129(_add_all_x_data_in129), .data_in130(_add_all_x_data_in130), .data_in131(_add_all_x_data_in131), .data_in132(_add_all_x_data_in132), .data_in133(_add_all_x_data_in133), .data_in134(_add_all_x_data_in134), .data_in135(_add_all_x_data_in135), .data_in136(_add_all_x_data_in136), .data_in137(_add_all_x_data_in137), .data_in138(_add_all_x_data_in138), .data_in139(_add_all_x_data_in139), .data_in140(_add_all_x_data_in140), .data_in141(_add_all_x_data_in141), .data_in142(_add_all_x_data_in142), .data_in143(_add_all_x_data_in143), .data_in144(_add_all_x_data_in144), .data_in145(_add_all_x_data_in145), .data_in146(_add_all_x_data_in146), .data_in147(_add_all_x_data_in147), .data_in148(_add_all_x_data_in148), .data_in149(_add_all_x_data_in149), .data_in150(_add_all_x_data_in150), .data_in151(_add_all_x_data_in151), .data_in152(_add_all_x_data_in152), .data_in153(_add_all_x_data_in153), .data_in154(_add_all_x_data_in154), .data_in155(_add_all_x_data_in155), .data_in156(_add_all_x_data_in156), .data_in157(_add_all_x_data_in157), .data_in158(_add_all_x_data_in158), .data_in161(_add_all_x_data_in161), .data_in162(_add_all_x_data_in162), .data_in163(_add_all_x_data_in163), .data_in164(_add_all_x_data_in164), .data_in165(_add_all_x_data_in165), .data_in166(_add_all_x_data_in166), .data_in167(_add_all_x_data_in167), .data_in168(_add_all_x_data_in168), .data_in169(_add_all_x_data_in169), .data_in170(_add_all_x_data_in170), .data_in171(_add_all_x_data_in171), .data_in172(_add_all_x_data_in172), .data_in173(_add_all_x_data_in173), .data_in174(_add_all_x_data_in174), .data_in175(_add_all_x_data_in175), .data_in176(_add_all_x_data_in176), .data_in177(_add_all_x_data_in177), .data_in178(_add_all_x_data_in178), .data_in179(_add_all_x_data_in179), .data_in180(_add_all_x_data_in180), .data_in181(_add_all_x_data_in181), .data_in182(_add_all_x_data_in182), .data_in183(_add_all_x_data_in183), .data_in184(_add_all_x_data_in184), .data_in185(_add_all_x_data_in185), .data_in186(_add_all_x_data_in186), .data_in187(_add_all_x_data_in187), .data_in188(_add_all_x_data_in188), .data_in189(_add_all_x_data_in189), .data_in190(_add_all_x_data_in190), .data_in193(_add_all_x_data_in193), .data_in194(_add_all_x_data_in194), .data_in195(_add_all_x_data_in195), .data_in196(_add_all_x_data_in196), .data_in197(_add_all_x_data_in197), .data_in198(_add_all_x_data_in198), .data_in199(_add_all_x_data_in199), .data_in200(_add_all_x_data_in200), .data_in201(_add_all_x_data_in201), .data_in202(_add_all_x_data_in202), .data_in203(_add_all_x_data_in203), .data_in204(_add_all_x_data_in204), .data_in205(_add_all_x_data_in205), .data_in206(_add_all_x_data_in206), .data_in207(_add_all_x_data_in207), .data_in208(_add_all_x_data_in208), .data_in209(_add_all_x_data_in209), .data_in210(_add_all_x_data_in210), .data_in211(_add_all_x_data_in211), .data_in212(_add_all_x_data_in212), .data_in213(_add_all_x_data_in213), .data_in214(_add_all_x_data_in214), .data_in215(_add_all_x_data_in215), .data_in216(_add_all_x_data_in216), .data_in217(_add_all_x_data_in217), .data_in218(_add_all_x_data_in218), .data_in219(_add_all_x_data_in219), .data_in220(_add_all_x_data_in220), .data_in221(_add_all_x_data_in221), .data_in222(_add_all_x_data_in222), .data_in225(_add_all_x_data_in225), .data_in226(_add_all_x_data_in226), .data_in227(_add_all_x_data_in227), .data_in228(_add_all_x_data_in228), .data_in229(_add_all_x_data_in229), .data_in230(_add_all_x_data_in230), .data_in231(_add_all_x_data_in231), .data_in232(_add_all_x_data_in232), .data_in233(_add_all_x_data_in233), .data_in234(_add_all_x_data_in234), .data_in235(_add_all_x_data_in235), .data_in236(_add_all_x_data_in236), .data_in237(_add_all_x_data_in237), .data_in238(_add_all_x_data_in238), .data_in239(_add_all_x_data_in239), .data_in240(_add_all_x_data_in240), .data_in241(_add_all_x_data_in241), .data_in242(_add_all_x_data_in242), .data_in243(_add_all_x_data_in243), .data_in244(_add_all_x_data_in244), .data_in245(_add_all_x_data_in245), .data_in246(_add_all_x_data_in246), .data_in247(_add_all_x_data_in247), .data_in248(_add_all_x_data_in248), .data_in249(_add_all_x_data_in249), .data_in250(_add_all_x_data_in250), .data_in251(_add_all_x_data_in251), .data_in252(_add_all_x_data_in252), .data_in253(_add_all_x_data_in253), .data_in254(_add_all_x_data_in254), .data_in257(_add_all_x_data_in257), .data_in258(_add_all_x_data_in258), .data_in259(_add_all_x_data_in259), .data_in260(_add_all_x_data_in260), .data_in261(_add_all_x_data_in261), .data_in262(_add_all_x_data_in262), .data_in263(_add_all_x_data_in263), .data_in264(_add_all_x_data_in264), .data_in265(_add_all_x_data_in265), .data_in266(_add_all_x_data_in266), .data_in267(_add_all_x_data_in267), .data_in268(_add_all_x_data_in268), .data_in269(_add_all_x_data_in269), .data_in270(_add_all_x_data_in270), .data_in271(_add_all_x_data_in271), .data_in272(_add_all_x_data_in272), .data_in273(_add_all_x_data_in273), .data_in274(_add_all_x_data_in274), .data_in275(_add_all_x_data_in275), .data_in276(_add_all_x_data_in276), .data_in277(_add_all_x_data_in277), .data_in278(_add_all_x_data_in278), .data_in279(_add_all_x_data_in279), .data_in280(_add_all_x_data_in280), .data_in281(_add_all_x_data_in281), .data_in282(_add_all_x_data_in282), .data_in283(_add_all_x_data_in283), .data_in284(_add_all_x_data_in284), .data_in285(_add_all_x_data_in285), .data_in286(_add_all_x_data_in286), .data_in289(_add_all_x_data_in289), .data_in290(_add_all_x_data_in290), .data_in291(_add_all_x_data_in291), .data_in292(_add_all_x_data_in292), .data_in293(_add_all_x_data_in293), .data_in294(_add_all_x_data_in294), .data_in295(_add_all_x_data_in295), .data_in296(_add_all_x_data_in296), .data_in297(_add_all_x_data_in297), .data_in298(_add_all_x_data_in298), .data_in299(_add_all_x_data_in299), .data_in300(_add_all_x_data_in300), .data_in301(_add_all_x_data_in301), .data_in302(_add_all_x_data_in302), .data_in303(_add_all_x_data_in303), .data_in304(_add_all_x_data_in304), .data_in305(_add_all_x_data_in305), .data_in306(_add_all_x_data_in306), .data_in307(_add_all_x_data_in307), .data_in308(_add_all_x_data_in308), .data_in309(_add_all_x_data_in309), .data_in310(_add_all_x_data_in310), .data_in311(_add_all_x_data_in311), .data_in312(_add_all_x_data_in312), .data_in313(_add_all_x_data_in313), .data_in314(_add_all_x_data_in314), .data_in315(_add_all_x_data_in315), .data_in316(_add_all_x_data_in316), .data_in317(_add_all_x_data_in317), .data_in318(_add_all_x_data_in318), .data_in321(_add_all_x_data_in321), .data_in322(_add_all_x_data_in322), .data_in323(_add_all_x_data_in323), .data_in324(_add_all_x_data_in324), .data_in325(_add_all_x_data_in325), .data_in326(_add_all_x_data_in326), .data_in327(_add_all_x_data_in327), .data_in328(_add_all_x_data_in328), .data_in329(_add_all_x_data_in329), .data_in330(_add_all_x_data_in330), .data_in331(_add_all_x_data_in331), .data_in332(_add_all_x_data_in332), .data_in333(_add_all_x_data_in333), .data_in334(_add_all_x_data_in334), .data_in335(_add_all_x_data_in335), .data_in336(_add_all_x_data_in336), .data_in337(_add_all_x_data_in337), .data_in338(_add_all_x_data_in338), .data_in339(_add_all_x_data_in339), .data_in340(_add_all_x_data_in340), .data_in341(_add_all_x_data_in341), .data_in342(_add_all_x_data_in342), .data_in343(_add_all_x_data_in343), .data_in344(_add_all_x_data_in344), .data_in345(_add_all_x_data_in345), .data_in346(_add_all_x_data_in346), .data_in347(_add_all_x_data_in347), .data_in348(_add_all_x_data_in348), .data_in349(_add_all_x_data_in349), .data_in350(_add_all_x_data_in350), .data_in353(_add_all_x_data_in353), .data_in354(_add_all_x_data_in354), .data_in355(_add_all_x_data_in355), .data_in356(_add_all_x_data_in356), .data_in357(_add_all_x_data_in357), .data_in358(_add_all_x_data_in358), .data_in359(_add_all_x_data_in359), .data_in360(_add_all_x_data_in360), .data_in361(_add_all_x_data_in361), .data_in362(_add_all_x_data_in362), .data_in363(_add_all_x_data_in363), .data_in364(_add_all_x_data_in364), .data_in365(_add_all_x_data_in365), .data_in366(_add_all_x_data_in366), .data_in367(_add_all_x_data_in367), .data_in368(_add_all_x_data_in368), .data_in369(_add_all_x_data_in369), .data_in370(_add_all_x_data_in370), .data_in371(_add_all_x_data_in371), .data_in372(_add_all_x_data_in372), .data_in373(_add_all_x_data_in373), .data_in374(_add_all_x_data_in374), .data_in375(_add_all_x_data_in375), .data_in376(_add_all_x_data_in376), .data_in377(_add_all_x_data_in377), .data_in378(_add_all_x_data_in378), .data_in379(_add_all_x_data_in379), .data_in380(_add_all_x_data_in380), .data_in381(_add_all_x_data_in381), .data_in382(_add_all_x_data_in382), .data_in385(_add_all_x_data_in385), .data_in386(_add_all_x_data_in386), .data_in387(_add_all_x_data_in387), .data_in388(_add_all_x_data_in388), .data_in389(_add_all_x_data_in389), .data_in390(_add_all_x_data_in390), .data_in391(_add_all_x_data_in391), .data_in392(_add_all_x_data_in392), .data_in393(_add_all_x_data_in393), .data_in394(_add_all_x_data_in394), .data_in395(_add_all_x_data_in395), .data_in396(_add_all_x_data_in396), .data_in397(_add_all_x_data_in397), .data_in398(_add_all_x_data_in398), .data_in399(_add_all_x_data_in399), .data_in400(_add_all_x_data_in400), .data_in401(_add_all_x_data_in401), .data_in402(_add_all_x_data_in402), .data_in403(_add_all_x_data_in403), .data_in404(_add_all_x_data_in404), .data_in405(_add_all_x_data_in405), .data_in406(_add_all_x_data_in406), .data_in407(_add_all_x_data_in407), .data_in408(_add_all_x_data_in408), .data_in409(_add_all_x_data_in409), .data_in410(_add_all_x_data_in410), .data_in411(_add_all_x_data_in411), .data_in412(_add_all_x_data_in412), .data_in413(_add_all_x_data_in413), .data_in414(_add_all_x_data_in414), .data_in417(_add_all_x_data_in417), .data_in418(_add_all_x_data_in418), .data_in419(_add_all_x_data_in419), .data_in420(_add_all_x_data_in420), .data_in421(_add_all_x_data_in421), .data_in422(_add_all_x_data_in422), .data_in423(_add_all_x_data_in423), .data_in424(_add_all_x_data_in424), .data_in425(_add_all_x_data_in425), .data_in426(_add_all_x_data_in426), .data_in427(_add_all_x_data_in427), .data_in428(_add_all_x_data_in428), .data_in429(_add_all_x_data_in429), .data_in430(_add_all_x_data_in430), .data_in431(_add_all_x_data_in431), .data_in432(_add_all_x_data_in432), .data_in433(_add_all_x_data_in433), .data_in434(_add_all_x_data_in434), .data_in435(_add_all_x_data_in435), .data_in436(_add_all_x_data_in436), .data_in437(_add_all_x_data_in437), .data_in438(_add_all_x_data_in438), .data_in439(_add_all_x_data_in439), .data_in440(_add_all_x_data_in440), .data_in441(_add_all_x_data_in441), .data_in442(_add_all_x_data_in442), .data_in443(_add_all_x_data_in443), .data_in444(_add_all_x_data_in444), .data_in445(_add_all_x_data_in445), .data_in446(_add_all_x_data_in446), .data_in449(_add_all_x_data_in449), .data_in450(_add_all_x_data_in450), .data_in451(_add_all_x_data_in451), .data_in452(_add_all_x_data_in452), .data_in453(_add_all_x_data_in453), .data_in454(_add_all_x_data_in454), .data_in455(_add_all_x_data_in455), .data_in456(_add_all_x_data_in456), .data_in457(_add_all_x_data_in457), .data_in458(_add_all_x_data_in458), .data_in459(_add_all_x_data_in459), .data_in460(_add_all_x_data_in460), .data_in461(_add_all_x_data_in461), .data_in462(_add_all_x_data_in462), .data_in463(_add_all_x_data_in463), .data_in464(_add_all_x_data_in464), .data_in465(_add_all_x_data_in465), .data_in466(_add_all_x_data_in466), .data_in467(_add_all_x_data_in467), .data_in468(_add_all_x_data_in468), .data_in469(_add_all_x_data_in469), .data_in470(_add_all_x_data_in470), .data_in471(_add_all_x_data_in471), .data_in472(_add_all_x_data_in472), .data_in473(_add_all_x_data_in473), .data_in474(_add_all_x_data_in474), .data_in475(_add_all_x_data_in475), .data_in476(_add_all_x_data_in476), .data_in477(_add_all_x_data_in477), .data_in478(_add_all_x_data_in478), .sig(_add_all_x_sig), .start(_add_all_x_start), .goal(_add_all_x_goal), .dig_w(_add_all_x_dig_w));

   assign  dig_exit = (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_add_all_x_dig_t0|_add_all_x_dig_t1)|_add_all_x_dig_t2)|_add_all_x_dig_t3)|_add_all_x_dig_t4)|_add_all_x_dig_t5)|_add_all_x_dig_t6)|_add_all_x_dig_t7)|_add_all_x_dig_t8)|_add_all_x_dig_t9)|_add_all_x_dig_t10)|_add_all_x_dig_t11)|_add_all_x_dig_t12)|_add_all_x_dig_t13)|_add_all_x_dig_t14)|_add_all_x_dig_t15)|_add_all_x_dig_t16)|_add_all_x_dig_t17)|_add_all_x_dig_t18)|_add_all_x_dig_t19)|_add_all_x_dig_t20)|_add_all_x_dig_t21)|_add_all_x_dig_t22)|_add_all_x_dig_t23)|_add_all_x_dig_t24)|_add_all_x_dig_t25)|_add_all_x_dig_t26)|_add_all_x_dig_t27)|_add_all_x_dig_t28)|_add_all_x_dig_t29)|_add_all_x_dig_t30)|_add_all_x_dig_t31)|_add_all_x_dig_t32)|_add_all_x_dig_t33)|_add_all_x_dig_t34)|_add_all_x_dig_t35)|_add_all_x_dig_t36)|_add_all_x_dig_t37)|_add_all_x_dig_t38)|_add_all_x_dig_t39)|_add_all_x_dig_t40)|_add_all_x_dig_t41)|_add_all_x_dig_t42)|_add_all_x_dig_t43)|_add_all_x_dig_t44)|_add_all_x_dig_t45)|_add_all_x_dig_t46)|_add_all_x_dig_t47)|_add_all_x_dig_t48)|_add_all_x_dig_t49)|_add_all_x_dig_t50)|_add_all_x_dig_t51)|_add_all_x_dig_t52)|_add_all_x_dig_t53)|_add_all_x_dig_t54)|_add_all_x_dig_t55)|_add_all_x_dig_t56)|_add_all_x_dig_t57)|_add_all_x_dig_t58)|_add_all_x_dig_t59)|_add_all_x_dig_t60)|_add_all_x_dig_t61)|_add_all_x_dig_t62)|_add_all_x_dig_t63)|_add_all_x_dig_t64)|_add_all_x_dig_t65)|_add_all_x_dig_t66)|_add_all_x_dig_t67)|_add_all_x_dig_t68)|_add_all_x_dig_t69)|_add_all_x_dig_t70)|_add_all_x_dig_t71)|_add_all_x_dig_t72)|_add_all_x_dig_t73)|_add_all_x_dig_t74)|_add_all_x_dig_t75)|_add_all_x_dig_t76)|_add_all_x_dig_t77)|_add_all_x_dig_t78)|_add_all_x_dig_t79)|_add_all_x_dig_t80)|_add_all_x_dig_t81)|_add_all_x_dig_t82)|_add_all_x_dig_t83)|_add_all_x_dig_t84)|_add_all_x_dig_t85)|_add_all_x_dig_t86)|_add_all_x_dig_t87)|_add_all_x_dig_t88)|_add_all_x_dig_t89)|_add_all_x_dig_t90)|_add_all_x_dig_t91)|_add_all_x_dig_t92)|_add_all_x_dig_t93)|_add_all_x_dig_t94)|_add_all_x_dig_t95)|_add_all_x_dig_t96)|_add_all_x_dig_t97)|_add_all_x_dig_t98)|_add_all_x_dig_t99)|_add_all_x_dig_t100)|_add_all_x_dig_t101)|_add_all_x_dig_t102)|_add_all_x_dig_t103)|_add_all_x_dig_t104)|_add_all_x_dig_t105)|_add_all_x_dig_t106)|_add_all_x_dig_t107)|_add_all_x_dig_t108)|_add_all_x_dig_t109)|_add_all_x_dig_t110)|_add_all_x_dig_t111)|_add_all_x_dig_t112)|_add_all_x_dig_t113)|_add_all_x_dig_t114)|_add_all_x_dig_t115)|_add_all_x_dig_t116)|_add_all_x_dig_t117)|_add_all_x_dig_t118)|_add_all_x_dig_t119)|_add_all_x_dig_t120)|_add_all_x_dig_t121)|_add_all_x_dig_t122)|_add_all_x_dig_t123)|_add_all_x_dig_t124)|_add_all_x_dig_t125)|_add_all_x_dig_t126)|_add_all_x_dig_t127)|_add_all_x_dig_t128)|_add_all_x_dig_t129)|_add_all_x_dig_t130)|_add_all_x_dig_t131)|_add_all_x_dig_t132)|_add_all_x_dig_t133)|_add_all_x_dig_t134)|_add_all_x_dig_t135)|_add_all_x_dig_t136)|_add_all_x_dig_t137)|_add_all_x_dig_t138)|_add_all_x_dig_t139)|_add_all_x_dig_t140)|_add_all_x_dig_t141)|_add_all_x_dig_t142)|_add_all_x_dig_t143)|_add_all_x_dig_t144)|_add_all_x_dig_t145)|_add_all_x_dig_t146)|_add_all_x_dig_t147)|_add_all_x_dig_t148)|_add_all_x_dig_t149)|_add_all_x_dig_t150)|_add_all_x_dig_t151)|_add_all_x_dig_t152)|_add_all_x_dig_t153)|_add_all_x_dig_t154)|_add_all_x_dig_t155)|_add_all_x_dig_t156)|_add_all_x_dig_t157)|_add_all_x_dig_t158)|_add_all_x_dig_t159)|_add_all_x_dig_t160)|_add_all_x_dig_t161)|_add_all_x_dig_t162)|_add_all_x_dig_t163)|_add_all_x_dig_t164)|_add_all_x_dig_t165)|_add_all_x_dig_t166)|_add_all_x_dig_t167)|_add_all_x_dig_t168)|_add_all_x_dig_t169)|_add_all_x_dig_t170)|_add_all_x_dig_t171)|_add_all_x_dig_t172)|_add_all_x_dig_t173)|_add_all_x_dig_t174)|_add_all_x_dig_t175)|_add_all_x_dig_t176)|_add_all_x_dig_t177)|_add_all_x_dig_t178)|_add_all_x_dig_t179)|_add_all_x_dig_t180)|_add_all_x_dig_t181)|_add_all_x_dig_t182)|_add_all_x_dig_t183)|_add_all_x_dig_t184)|_add_all_x_dig_t185)|_add_all_x_dig_t186)|_add_all_x_dig_t187)|_add_all_x_dig_t188)|_add_all_x_dig_t189)|_add_all_x_dig_t190)|_add_all_x_dig_t191)|_add_all_x_dig_t192)|_add_all_x_dig_t193)|_add_all_x_dig_t194)|_add_all_x_dig_t195)|_add_all_x_dig_t196)|_add_all_x_dig_t197)|_add_all_x_dig_t198)|_add_all_x_dig_t199)|_add_all_x_dig_t200)|_add_all_x_dig_t201)|_add_all_x_dig_t202)|_add_all_x_dig_t203)|_add_all_x_dig_t204)|_add_all_x_dig_t205)|_add_all_x_dig_t206)|_add_all_x_dig_t207)|_add_all_x_dig_t208)|_add_all_x_dig_t209);
   assign  even_w1 = ((_reg_2)?1'b0:1'b0)|
    (((_net_1279|_net_9))?1'b1:1'b0);
   assign  start_wire = ((_net_1278)?start:10'b0)|
    (((_reg_2|_net_8))?start_reg:10'b0);
   assign  goal_wire = ((_net_1277)?goal:10'b0)|
    (((_reg_2|_net_7))?goal_reg:10'b0);
   assign  wall_w = ((_net_1276)?1'b0:1'b0)|
    (((_reg_2|_net_6))?dig_exit:1'b0);
   assign  data_wire33 = ((_net_2539)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1269))?_add_all_x_data_out33:10'b0);
   assign  data_wire34 = ((_net_2538)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1268))?_add_all_x_data_out34:10'b0);
   assign  data_wire35 = ((_net_2537)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1267))?_add_all_x_data_out35:10'b0);
   assign  data_wire36 = ((_net_2536)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1266))?_add_all_x_data_out36:10'b0);
   assign  data_wire37 = ((_net_2535)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1265))?_add_all_x_data_out37:10'b0);
   assign  data_wire38 = ((_net_2534)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1264))?_add_all_x_data_out38:10'b0);
   assign  data_wire39 = ((_net_2533)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1263))?_add_all_x_data_out39:10'b0);
   assign  data_wire40 = ((_net_2532)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1262))?_add_all_x_data_out40:10'b0);
   assign  data_wire41 = ((_net_2531)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1261))?_add_all_x_data_out41:10'b0);
   assign  data_wire42 = ((_net_2530)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1260))?_add_all_x_data_out42:10'b0);
   assign  data_wire43 = ((_net_2529)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1259))?_add_all_x_data_out43:10'b0);
   assign  data_wire44 = ((_net_2528)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1258))?_add_all_x_data_out44:10'b0);
   assign  data_wire45 = ((_net_2527)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1257))?_add_all_x_data_out45:10'b0);
   assign  data_wire46 = ((_net_2526)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1256))?_add_all_x_data_out46:10'b0);
   assign  data_wire47 = ((_net_2525)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1255))?_add_all_x_data_out47:10'b0);
   assign  data_wire48 = ((_net_2524)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1254))?_add_all_x_data_out48:10'b0);
   assign  data_wire49 = ((_net_2523)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1253))?_add_all_x_data_out49:10'b0);
   assign  data_wire50 = ((_net_2522)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1252))?_add_all_x_data_out50:10'b0);
   assign  data_wire51 = ((_net_2521)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1251))?_add_all_x_data_out51:10'b0);
   assign  data_wire52 = ((_net_2520)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1250))?_add_all_x_data_out52:10'b0);
   assign  data_wire53 = ((_net_2519)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1249))?_add_all_x_data_out53:10'b0);
   assign  data_wire54 = ((_net_2518)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1248))?_add_all_x_data_out54:10'b0);
   assign  data_wire55 = ((_net_2517)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1247))?_add_all_x_data_out55:10'b0);
   assign  data_wire56 = ((_net_2516)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1246))?_add_all_x_data_out56:10'b0);
   assign  data_wire57 = ((_net_2515)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1245))?_add_all_x_data_out57:10'b0);
   assign  data_wire58 = ((_net_2514)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1244))?_add_all_x_data_out58:10'b0);
   assign  data_wire59 = ((_net_2513)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1243))?_add_all_x_data_out59:10'b0);
   assign  data_wire60 = ((_net_2512)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1242))?_add_all_x_data_out60:10'b0);
   assign  data_wire61 = ((_net_2511)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1241))?_add_all_x_data_out61:10'b0);
   assign  data_wire62 = ((_net_2510)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1240))?_add_all_x_data_out62:10'b0);
   assign  data_wire65 = ((_net_2509)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1239))?_add_all_x_data_out65:10'b0);
   assign  data_wire66 = ((_net_2508)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1238))?_add_all_x_data_out66:10'b0);
   assign  data_wire67 = ((_net_2507)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1237))?_add_all_x_data_out67:10'b0);
   assign  data_wire68 = ((_net_2506)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1236))?_add_all_x_data_out68:10'b0);
   assign  data_wire69 = ((_net_2505)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1235))?_add_all_x_data_out69:10'b0);
   assign  data_wire70 = ((_net_2504)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1234))?_add_all_x_data_out70:10'b0);
   assign  data_wire71 = ((_net_2503)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1233))?_add_all_x_data_out71:10'b0);
   assign  data_wire72 = ((_net_2502)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1232))?_add_all_x_data_out72:10'b0);
   assign  data_wire73 = ((_net_2501)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1231))?_add_all_x_data_out73:10'b0);
   assign  data_wire74 = ((_net_2500)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1230))?_add_all_x_data_out74:10'b0);
   assign  data_wire75 = ((_net_2499)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1229))?_add_all_x_data_out75:10'b0);
   assign  data_wire76 = ((_net_2498)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1228))?_add_all_x_data_out76:10'b0);
   assign  data_wire77 = ((_net_2497)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1227))?_add_all_x_data_out77:10'b0);
   assign  data_wire78 = ((_net_2496)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1226))?_add_all_x_data_out78:10'b0);
   assign  data_wire79 = ((_net_2495)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1225))?_add_all_x_data_out79:10'b0);
   assign  data_wire80 = ((_net_2494)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1224))?_add_all_x_data_out80:10'b0);
   assign  data_wire81 = ((_net_2493)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1223))?_add_all_x_data_out81:10'b0);
   assign  data_wire82 = ((_net_2492)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1222))?_add_all_x_data_out82:10'b0);
   assign  data_wire83 = ((_net_2491)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1221))?_add_all_x_data_out83:10'b0);
   assign  data_wire84 = ((_net_2490)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1220))?_add_all_x_data_out84:10'b0);
   assign  data_wire85 = ((_net_2489)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1219))?_add_all_x_data_out85:10'b0);
   assign  data_wire86 = ((_net_2488)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1218))?_add_all_x_data_out86:10'b0);
   assign  data_wire87 = ((_net_2487)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1217))?_add_all_x_data_out87:10'b0);
   assign  data_wire88 = ((_net_2486)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1216))?_add_all_x_data_out88:10'b0);
   assign  data_wire89 = ((_net_2485)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1215))?_add_all_x_data_out89:10'b0);
   assign  data_wire90 = ((_net_2484)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1214))?_add_all_x_data_out90:10'b0);
   assign  data_wire91 = ((_net_2483)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1213))?_add_all_x_data_out91:10'b0);
   assign  data_wire92 = ((_net_2482)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1212))?_add_all_x_data_out92:10'b0);
   assign  data_wire93 = ((_net_2481)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1211))?_add_all_x_data_out93:10'b0);
   assign  data_wire94 = ((_net_2480)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1210))?_add_all_x_data_out94:10'b0);
   assign  data_wire97 = ((_net_2479)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1209))?_add_all_x_data_out97:10'b0);
   assign  data_wire98 = ((_net_2478)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1208))?_add_all_x_data_out98:10'b0);
   assign  data_wire99 = ((_net_2477)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1207))?_add_all_x_data_out99:10'b0);
   assign  data_wire100 = ((_net_2476)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1206))?_add_all_x_data_out100:10'b0);
   assign  data_wire101 = ((_net_2475)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1205))?_add_all_x_data_out101:10'b0);
   assign  data_wire102 = ((_net_2474)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1204))?_add_all_x_data_out102:10'b0);
   assign  data_wire103 = ((_net_2473)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1203))?_add_all_x_data_out103:10'b0);
   assign  data_wire104 = ((_net_2472)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1202))?_add_all_x_data_out104:10'b0);
   assign  data_wire105 = ((_net_2471)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1201))?_add_all_x_data_out105:10'b0);
   assign  data_wire106 = ((_net_2470)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1200))?_add_all_x_data_out106:10'b0);
   assign  data_wire107 = ((_net_2469)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1199))?_add_all_x_data_out107:10'b0);
   assign  data_wire108 = ((_net_2468)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1198))?_add_all_x_data_out108:10'b0);
   assign  data_wire109 = ((_net_2467)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1197))?_add_all_x_data_out109:10'b0);
   assign  data_wire110 = ((_net_2466)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1196))?_add_all_x_data_out110:10'b0);
   assign  data_wire111 = ((_net_2465)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1195))?_add_all_x_data_out111:10'b0);
   assign  data_wire112 = ((_net_2464)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1194))?_add_all_x_data_out112:10'b0);
   assign  data_wire113 = ((_net_2463)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1193))?_add_all_x_data_out113:10'b0);
   assign  data_wire114 = ((_net_2462)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1192))?_add_all_x_data_out114:10'b0);
   assign  data_wire115 = ((_net_2461)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1191))?_add_all_x_data_out115:10'b0);
   assign  data_wire116 = ((_net_2460)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1190))?_add_all_x_data_out116:10'b0);
   assign  data_wire117 = ((_net_2459)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1189))?_add_all_x_data_out117:10'b0);
   assign  data_wire118 = ((_net_2458)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1188))?_add_all_x_data_out118:10'b0);
   assign  data_wire119 = ((_net_2457)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1187))?_add_all_x_data_out119:10'b0);
   assign  data_wire120 = ((_net_2456)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1186))?_add_all_x_data_out120:10'b0);
   assign  data_wire121 = ((_net_2455)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1185))?_add_all_x_data_out121:10'b0);
   assign  data_wire122 = ((_net_2454)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1184))?_add_all_x_data_out122:10'b0);
   assign  data_wire123 = ((_net_2453)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1183))?_add_all_x_data_out123:10'b0);
   assign  data_wire124 = ((_net_2452)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1182))?_add_all_x_data_out124:10'b0);
   assign  data_wire125 = ((_net_2451)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1181))?_add_all_x_data_out125:10'b0);
   assign  data_wire126 = ((_net_2450)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1180))?_add_all_x_data_out126:10'b0);
   assign  data_wire129 = ((_net_2449)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1179))?_add_all_x_data_out129:10'b0);
   assign  data_wire130 = ((_net_2448)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1178))?_add_all_x_data_out130:10'b0);
   assign  data_wire131 = ((_net_2447)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1177))?_add_all_x_data_out131:10'b0);
   assign  data_wire132 = ((_net_2446)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1176))?_add_all_x_data_out132:10'b0);
   assign  data_wire133 = ((_net_2445)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1175))?_add_all_x_data_out133:10'b0);
   assign  data_wire134 = ((_net_2444)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1174))?_add_all_x_data_out134:10'b0);
   assign  data_wire135 = ((_net_2443)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1173))?_add_all_x_data_out135:10'b0);
   assign  data_wire136 = ((_net_2442)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1172))?_add_all_x_data_out136:10'b0);
   assign  data_wire137 = ((_net_2441)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1171))?_add_all_x_data_out137:10'b0);
   assign  data_wire138 = ((_net_2440)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1170))?_add_all_x_data_out138:10'b0);
   assign  data_wire139 = ((_net_2439)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1169))?_add_all_x_data_out139:10'b0);
   assign  data_wire140 = ((_net_2438)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1168))?_add_all_x_data_out140:10'b0);
   assign  data_wire141 = ((_net_2437)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1167))?_add_all_x_data_out141:10'b0);
   assign  data_wire142 = ((_net_2436)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1166))?_add_all_x_data_out142:10'b0);
   assign  data_wire143 = ((_net_2435)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1165))?_add_all_x_data_out143:10'b0);
   assign  data_wire144 = ((_net_2434)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1164))?_add_all_x_data_out144:10'b0);
   assign  data_wire145 = ((_net_2433)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1163))?_add_all_x_data_out145:10'b0);
   assign  data_wire146 = ((_net_2432)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1162))?_add_all_x_data_out146:10'b0);
   assign  data_wire147 = ((_net_2431)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1161))?_add_all_x_data_out147:10'b0);
   assign  data_wire148 = ((_net_2430)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1160))?_add_all_x_data_out148:10'b0);
   assign  data_wire149 = ((_net_2429)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1159))?_add_all_x_data_out149:10'b0);
   assign  data_wire150 = ((_net_2428)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1158))?_add_all_x_data_out150:10'b0);
   assign  data_wire151 = ((_net_2427)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1157))?_add_all_x_data_out151:10'b0);
   assign  data_wire152 = ((_net_2426)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1156))?_add_all_x_data_out152:10'b0);
   assign  data_wire153 = ((_net_2425)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1155))?_add_all_x_data_out153:10'b0);
   assign  data_wire154 = ((_net_2424)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1154))?_add_all_x_data_out154:10'b0);
   assign  data_wire155 = ((_net_2423)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1153))?_add_all_x_data_out155:10'b0);
   assign  data_wire156 = ((_net_2422)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1152))?_add_all_x_data_out156:10'b0);
   assign  data_wire157 = ((_net_2421)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1151))?_add_all_x_data_out157:10'b0);
   assign  data_wire158 = ((_net_2420)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1150))?_add_all_x_data_out158:10'b0);
   assign  data_wire161 = ((_net_2419)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1149))?_add_all_x_data_out161:10'b0);
   assign  data_wire162 = ((_net_2418)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1148))?_add_all_x_data_out162:10'b0);
   assign  data_wire163 = ((_net_2417)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1147))?_add_all_x_data_out163:10'b0);
   assign  data_wire164 = ((_net_2416)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1146))?_add_all_x_data_out164:10'b0);
   assign  data_wire165 = ((_net_2415)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1145))?_add_all_x_data_out165:10'b0);
   assign  data_wire166 = ((_net_2414)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1144))?_add_all_x_data_out166:10'b0);
   assign  data_wire167 = ((_net_2413)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1143))?_add_all_x_data_out167:10'b0);
   assign  data_wire168 = ((_net_2412)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1142))?_add_all_x_data_out168:10'b0);
   assign  data_wire169 = ((_net_2411)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1141))?_add_all_x_data_out169:10'b0);
   assign  data_wire170 = ((_net_2410)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1140))?_add_all_x_data_out170:10'b0);
   assign  data_wire171 = ((_net_2409)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1139))?_add_all_x_data_out171:10'b0);
   assign  data_wire172 = ((_net_2408)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1138))?_add_all_x_data_out172:10'b0);
   assign  data_wire173 = ((_net_2407)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1137))?_add_all_x_data_out173:10'b0);
   assign  data_wire174 = ((_net_2406)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1136))?_add_all_x_data_out174:10'b0);
   assign  data_wire175 = ((_net_2405)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1135))?_add_all_x_data_out175:10'b0);
   assign  data_wire176 = ((_net_2404)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1134))?_add_all_x_data_out176:10'b0);
   assign  data_wire177 = ((_net_2403)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1133))?_add_all_x_data_out177:10'b0);
   assign  data_wire178 = ((_net_2402)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1132))?_add_all_x_data_out178:10'b0);
   assign  data_wire179 = ((_net_2401)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1131))?_add_all_x_data_out179:10'b0);
   assign  data_wire180 = ((_net_2400)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1130))?_add_all_x_data_out180:10'b0);
   assign  data_wire181 = ((_net_2399)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1129))?_add_all_x_data_out181:10'b0);
   assign  data_wire182 = ((_net_2398)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1128))?_add_all_x_data_out182:10'b0);
   assign  data_wire183 = ((_net_2397)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1127))?_add_all_x_data_out183:10'b0);
   assign  data_wire184 = ((_net_2396)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1126))?_add_all_x_data_out184:10'b0);
   assign  data_wire185 = ((_net_2395)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1125))?_add_all_x_data_out185:10'b0);
   assign  data_wire186 = ((_net_2394)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1124))?_add_all_x_data_out186:10'b0);
   assign  data_wire187 = ((_net_2393)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1123))?_add_all_x_data_out187:10'b0);
   assign  data_wire188 = ((_net_2392)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1122))?_add_all_x_data_out188:10'b0);
   assign  data_wire189 = ((_net_2391)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1121))?_add_all_x_data_out189:10'b0);
   assign  data_wire190 = ((_net_2390)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1120))?_add_all_x_data_out190:10'b0);
   assign  data_wire193 = ((_net_2389)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1119))?_add_all_x_data_out193:10'b0);
   assign  data_wire194 = ((_net_2388)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1118))?_add_all_x_data_out194:10'b0);
   assign  data_wire195 = ((_net_2387)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1117))?_add_all_x_data_out195:10'b0);
   assign  data_wire196 = ((_net_2386)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1116))?_add_all_x_data_out196:10'b0);
   assign  data_wire197 = ((_net_2385)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1115))?_add_all_x_data_out197:10'b0);
   assign  data_wire198 = ((_net_2384)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1114))?_add_all_x_data_out198:10'b0);
   assign  data_wire199 = ((_net_2383)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1113))?_add_all_x_data_out199:10'b0);
   assign  data_wire200 = ((_net_2382)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1112))?_add_all_x_data_out200:10'b0);
   assign  data_wire201 = ((_net_2381)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1111))?_add_all_x_data_out201:10'b0);
   assign  data_wire202 = ((_net_2380)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1110))?_add_all_x_data_out202:10'b0);
   assign  data_wire203 = ((_net_2379)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1109))?_add_all_x_data_out203:10'b0);
   assign  data_wire204 = ((_net_2378)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1108))?_add_all_x_data_out204:10'b0);
   assign  data_wire205 = ((_net_2377)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1107))?_add_all_x_data_out205:10'b0);
   assign  data_wire206 = ((_net_2376)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1106))?_add_all_x_data_out206:10'b0);
   assign  data_wire207 = ((_net_2375)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1105))?_add_all_x_data_out207:10'b0);
   assign  data_wire208 = ((_net_2374)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1104))?_add_all_x_data_out208:10'b0);
   assign  data_wire209 = ((_net_2373)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1103))?_add_all_x_data_out209:10'b0);
   assign  data_wire210 = ((_net_2372)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1102))?_add_all_x_data_out210:10'b0);
   assign  data_wire211 = ((_net_2371)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1101))?_add_all_x_data_out211:10'b0);
   assign  data_wire212 = ((_net_2370)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1100))?_add_all_x_data_out212:10'b0);
   assign  data_wire213 = ((_net_2369)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1099))?_add_all_x_data_out213:10'b0);
   assign  data_wire214 = ((_net_2368)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1098))?_add_all_x_data_out214:10'b0);
   assign  data_wire215 = ((_net_2367)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1097))?_add_all_x_data_out215:10'b0);
   assign  data_wire216 = ((_net_2366)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1096))?_add_all_x_data_out216:10'b0);
   assign  data_wire217 = ((_net_2365)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1095))?_add_all_x_data_out217:10'b0);
   assign  data_wire218 = ((_net_2364)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1094))?_add_all_x_data_out218:10'b0);
   assign  data_wire219 = ((_net_2363)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1093))?_add_all_x_data_out219:10'b0);
   assign  data_wire220 = ((_net_2362)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1092))?_add_all_x_data_out220:10'b0);
   assign  data_wire221 = ((_net_2361)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1091))?_add_all_x_data_out221:10'b0);
   assign  data_wire222 = ((_net_2360)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1090))?_add_all_x_data_out222:10'b0);
   assign  data_wire225 = ((_net_2359)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1089))?_add_all_x_data_out225:10'b0);
   assign  data_wire226 = ((_net_2358)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1088))?_add_all_x_data_out226:10'b0);
   assign  data_wire227 = ((_net_2357)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1087))?_add_all_x_data_out227:10'b0);
   assign  data_wire228 = ((_net_2356)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1086))?_add_all_x_data_out228:10'b0);
   assign  data_wire229 = ((_net_2355)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1085))?_add_all_x_data_out229:10'b0);
   assign  data_wire230 = ((_net_2354)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1084))?_add_all_x_data_out230:10'b0);
   assign  data_wire231 = ((_net_2353)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1083))?_add_all_x_data_out231:10'b0);
   assign  data_wire232 = ((_net_2352)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1082))?_add_all_x_data_out232:10'b0);
   assign  data_wire233 = ((_net_2351)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1081))?_add_all_x_data_out233:10'b0);
   assign  data_wire234 = ((_net_2350)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1080))?_add_all_x_data_out234:10'b0);
   assign  data_wire235 = ((_net_2349)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1079))?_add_all_x_data_out235:10'b0);
   assign  data_wire236 = ((_net_2348)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1078))?_add_all_x_data_out236:10'b0);
   assign  data_wire237 = ((_net_2347)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1077))?_add_all_x_data_out237:10'b0);
   assign  data_wire238 = ((_net_2346)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1076))?_add_all_x_data_out238:10'b0);
   assign  data_wire239 = ((_net_2345)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1075))?_add_all_x_data_out239:10'b0);
   assign  data_wire240 = ((_net_2344)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1074))?_add_all_x_data_out240:10'b0);
   assign  data_wire241 = ((_net_2343)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1073))?_add_all_x_data_out241:10'b0);
   assign  data_wire242 = ((_net_2342)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1072))?_add_all_x_data_out242:10'b0);
   assign  data_wire243 = ((_net_2341)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1071))?_add_all_x_data_out243:10'b0);
   assign  data_wire244 = ((_net_2340)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1070))?_add_all_x_data_out244:10'b0);
   assign  data_wire245 = ((_net_2339)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1069))?_add_all_x_data_out245:10'b0);
   assign  data_wire246 = ((_net_2338)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1068))?_add_all_x_data_out246:10'b0);
   assign  data_wire247 = ((_net_2337)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1067))?_add_all_x_data_out247:10'b0);
   assign  data_wire248 = ((_net_2336)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1066))?_add_all_x_data_out248:10'b0);
   assign  data_wire249 = ((_net_2335)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1065))?_add_all_x_data_out249:10'b0);
   assign  data_wire250 = ((_net_2334)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1064))?_add_all_x_data_out250:10'b0);
   assign  data_wire251 = ((_net_2333)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1063))?_add_all_x_data_out251:10'b0);
   assign  data_wire252 = ((_net_2332)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1062))?_add_all_x_data_out252:10'b0);
   assign  data_wire253 = ((_net_2331)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1061))?_add_all_x_data_out253:10'b0);
   assign  data_wire254 = ((_net_2330)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1060))?_add_all_x_data_out254:10'b0);
   assign  data_wire257 = ((_net_2329)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1059))?_add_all_x_data_out257:10'b0);
   assign  data_wire258 = ((_net_2328)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1058))?_add_all_x_data_out258:10'b0);
   assign  data_wire259 = ((_net_2327)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1057))?_add_all_x_data_out259:10'b0);
   assign  data_wire260 = ((_net_2326)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1056))?_add_all_x_data_out260:10'b0);
   assign  data_wire261 = ((_net_2325)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1055))?_add_all_x_data_out261:10'b0);
   assign  data_wire262 = ((_net_2324)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1054))?_add_all_x_data_out262:10'b0);
   assign  data_wire263 = ((_net_2323)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1053))?_add_all_x_data_out263:10'b0);
   assign  data_wire264 = ((_net_2322)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1052))?_add_all_x_data_out264:10'b0);
   assign  data_wire265 = ((_net_2321)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1051))?_add_all_x_data_out265:10'b0);
   assign  data_wire266 = ((_net_2320)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1050))?_add_all_x_data_out266:10'b0);
   assign  data_wire267 = ((_net_2319)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1049))?_add_all_x_data_out267:10'b0);
   assign  data_wire268 = ((_net_2318)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1048))?_add_all_x_data_out268:10'b0);
   assign  data_wire269 = ((_net_2317)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1047))?_add_all_x_data_out269:10'b0);
   assign  data_wire270 = ((_net_2316)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1046))?_add_all_x_data_out270:10'b0);
   assign  data_wire271 = ((_net_2315)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1045))?_add_all_x_data_out271:10'b0);
   assign  data_wire272 = ((_net_2314)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1044))?_add_all_x_data_out272:10'b0);
   assign  data_wire273 = ((_net_2313)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1043))?_add_all_x_data_out273:10'b0);
   assign  data_wire274 = ((_net_2312)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1042))?_add_all_x_data_out274:10'b0);
   assign  data_wire275 = ((_net_2311)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1041))?_add_all_x_data_out275:10'b0);
   assign  data_wire276 = ((_net_2310)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1040))?_add_all_x_data_out276:10'b0);
   assign  data_wire277 = ((_net_2309)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1039))?_add_all_x_data_out277:10'b0);
   assign  data_wire278 = ((_net_2308)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1038))?_add_all_x_data_out278:10'b0);
   assign  data_wire279 = ((_net_2307)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1037))?_add_all_x_data_out279:10'b0);
   assign  data_wire280 = ((_net_2306)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1036))?_add_all_x_data_out280:10'b0);
   assign  data_wire281 = ((_net_2305)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1035))?_add_all_x_data_out281:10'b0);
   assign  data_wire282 = ((_net_2304)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1034))?_add_all_x_data_out282:10'b0);
   assign  data_wire283 = ((_net_2303)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1033))?_add_all_x_data_out283:10'b0);
   assign  data_wire284 = ((_net_2302)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1032))?_add_all_x_data_out284:10'b0);
   assign  data_wire285 = ((_net_2301)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1031))?_add_all_x_data_out285:10'b0);
   assign  data_wire286 = ((_net_2300)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1030))?_add_all_x_data_out286:10'b0);
   assign  data_wire289 = ((_net_2299)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1029))?_add_all_x_data_out289:10'b0);
   assign  data_wire290 = ((_net_2298)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1028))?_add_all_x_data_out290:10'b0);
   assign  data_wire291 = ((_net_2297)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1027))?_add_all_x_data_out291:10'b0);
   assign  data_wire292 = ((_net_2296)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1026))?_add_all_x_data_out292:10'b0);
   assign  data_wire293 = ((_net_2295)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1025))?_add_all_x_data_out293:10'b0);
   assign  data_wire294 = ((_net_2294)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1024))?_add_all_x_data_out294:10'b0);
   assign  data_wire295 = ((_net_2293)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1023))?_add_all_x_data_out295:10'b0);
   assign  data_wire296 = ((_net_2292)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1022))?_add_all_x_data_out296:10'b0);
   assign  data_wire297 = ((_net_2291)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1021))?_add_all_x_data_out297:10'b0);
   assign  data_wire298 = ((_net_2290)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1020))?_add_all_x_data_out298:10'b0);
   assign  data_wire299 = ((_net_2289)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1019))?_add_all_x_data_out299:10'b0);
   assign  data_wire300 = ((_net_2288)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1018))?_add_all_x_data_out300:10'b0);
   assign  data_wire301 = ((_net_2287)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1017))?_add_all_x_data_out301:10'b0);
   assign  data_wire302 = ((_net_2286)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1016))?_add_all_x_data_out302:10'b0);
   assign  data_wire303 = ((_net_2285)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1015))?_add_all_x_data_out303:10'b0);
   assign  data_wire304 = ((_net_2284)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1014))?_add_all_x_data_out304:10'b0);
   assign  data_wire305 = ((_net_2283)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1013))?_add_all_x_data_out305:10'b0);
   assign  data_wire306 = ((_net_2282)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1012))?_add_all_x_data_out306:10'b0);
   assign  data_wire307 = ((_net_2281)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1011))?_add_all_x_data_out307:10'b0);
   assign  data_wire308 = ((_net_2280)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1010))?_add_all_x_data_out308:10'b0);
   assign  data_wire309 = ((_net_2279)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1009))?_add_all_x_data_out309:10'b0);
   assign  data_wire310 = ((_net_2278)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1008))?_add_all_x_data_out310:10'b0);
   assign  data_wire311 = ((_net_2277)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1007))?_add_all_x_data_out311:10'b0);
   assign  data_wire312 = ((_net_2276)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1006))?_add_all_x_data_out312:10'b0);
   assign  data_wire313 = ((_net_2275)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1005))?_add_all_x_data_out313:10'b0);
   assign  data_wire314 = ((_net_2274)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1004))?_add_all_x_data_out314:10'b0);
   assign  data_wire315 = ((_net_2273)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1003))?_add_all_x_data_out315:10'b0);
   assign  data_wire316 = ((_net_2272)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1002))?_add_all_x_data_out316:10'b0);
   assign  data_wire317 = ((_net_2271)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1001))?_add_all_x_data_out317:10'b0);
   assign  data_wire318 = ((_net_2270)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_1000))?_add_all_x_data_out318:10'b0);
   assign  data_wire321 = ((_net_2269)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_999))?_add_all_x_data_out321:10'b0);
   assign  data_wire322 = ((_net_2268)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_998))?_add_all_x_data_out322:10'b0);
   assign  data_wire323 = ((_net_2267)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_997))?_add_all_x_data_out323:10'b0);
   assign  data_wire324 = ((_net_2266)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_996))?_add_all_x_data_out324:10'b0);
   assign  data_wire325 = ((_net_2265)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_995))?_add_all_x_data_out325:10'b0);
   assign  data_wire326 = ((_net_2264)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_994))?_add_all_x_data_out326:10'b0);
   assign  data_wire327 = ((_net_2263)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_993))?_add_all_x_data_out327:10'b0);
   assign  data_wire328 = ((_net_2262)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_992))?_add_all_x_data_out328:10'b0);
   assign  data_wire329 = ((_net_2261)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_991))?_add_all_x_data_out329:10'b0);
   assign  data_wire330 = ((_net_2260)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_990))?_add_all_x_data_out330:10'b0);
   assign  data_wire331 = ((_net_2259)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_989))?_add_all_x_data_out331:10'b0);
   assign  data_wire332 = ((_net_2258)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_988))?_add_all_x_data_out332:10'b0);
   assign  data_wire333 = ((_net_2257)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_987))?_add_all_x_data_out333:10'b0);
   assign  data_wire334 = ((_net_2256)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_986))?_add_all_x_data_out334:10'b0);
   assign  data_wire335 = ((_net_2255)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_985))?_add_all_x_data_out335:10'b0);
   assign  data_wire336 = ((_net_2254)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_984))?_add_all_x_data_out336:10'b0);
   assign  data_wire337 = ((_net_2253)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_983))?_add_all_x_data_out337:10'b0);
   assign  data_wire338 = ((_net_2252)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_982))?_add_all_x_data_out338:10'b0);
   assign  data_wire339 = ((_net_2251)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_981))?_add_all_x_data_out339:10'b0);
   assign  data_wire340 = ((_net_2250)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_980))?_add_all_x_data_out340:10'b0);
   assign  data_wire341 = ((_net_2249)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_979))?_add_all_x_data_out341:10'b0);
   assign  data_wire342 = ((_net_2248)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_978))?_add_all_x_data_out342:10'b0);
   assign  data_wire343 = ((_net_2247)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_977))?_add_all_x_data_out343:10'b0);
   assign  data_wire344 = ((_net_2246)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_976))?_add_all_x_data_out344:10'b0);
   assign  data_wire345 = ((_net_2245)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_975))?_add_all_x_data_out345:10'b0);
   assign  data_wire346 = ((_net_2244)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_974))?_add_all_x_data_out346:10'b0);
   assign  data_wire347 = ((_net_2243)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_973))?_add_all_x_data_out347:10'b0);
   assign  data_wire348 = ((_net_2242)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_972))?_add_all_x_data_out348:10'b0);
   assign  data_wire349 = ((_net_2241)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_971))?_add_all_x_data_out349:10'b0);
   assign  data_wire350 = ((_net_2240)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_970))?_add_all_x_data_out350:10'b0);
   assign  data_wire353 = ((_net_2239)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_969))?_add_all_x_data_out353:10'b0);
   assign  data_wire354 = ((_net_2238)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_968))?_add_all_x_data_out354:10'b0);
   assign  data_wire355 = ((_net_2237)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_967))?_add_all_x_data_out355:10'b0);
   assign  data_wire356 = ((_net_2236)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_966))?_add_all_x_data_out356:10'b0);
   assign  data_wire357 = ((_net_2235)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_965))?_add_all_x_data_out357:10'b0);
   assign  data_wire358 = ((_net_2234)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_964))?_add_all_x_data_out358:10'b0);
   assign  data_wire359 = ((_net_2233)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_963))?_add_all_x_data_out359:10'b0);
   assign  data_wire360 = ((_net_2232)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_962))?_add_all_x_data_out360:10'b0);
   assign  data_wire361 = ((_net_2231)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_961))?_add_all_x_data_out361:10'b0);
   assign  data_wire362 = ((_net_2230)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_960))?_add_all_x_data_out362:10'b0);
   assign  data_wire363 = ((_net_2229)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_959))?_add_all_x_data_out363:10'b0);
   assign  data_wire364 = ((_net_2228)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_958))?_add_all_x_data_out364:10'b0);
   assign  data_wire365 = ((_net_2227)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_957))?_add_all_x_data_out365:10'b0);
   assign  data_wire366 = ((_net_2226)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_956))?_add_all_x_data_out366:10'b0);
   assign  data_wire367 = ((_net_2225)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_955))?_add_all_x_data_out367:10'b0);
   assign  data_wire368 = ((_net_2224)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_954))?_add_all_x_data_out368:10'b0);
   assign  data_wire369 = ((_net_2223)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_953))?_add_all_x_data_out369:10'b0);
   assign  data_wire370 = ((_net_2222)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_952))?_add_all_x_data_out370:10'b0);
   assign  data_wire371 = ((_net_2221)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_951))?_add_all_x_data_out371:10'b0);
   assign  data_wire372 = ((_net_2220)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_950))?_add_all_x_data_out372:10'b0);
   assign  data_wire373 = ((_net_2219)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_949))?_add_all_x_data_out373:10'b0);
   assign  data_wire374 = ((_net_2218)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_948))?_add_all_x_data_out374:10'b0);
   assign  data_wire375 = ((_net_2217)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_947))?_add_all_x_data_out375:10'b0);
   assign  data_wire376 = ((_net_2216)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_946))?_add_all_x_data_out376:10'b0);
   assign  data_wire377 = ((_net_2215)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_945))?_add_all_x_data_out377:10'b0);
   assign  data_wire378 = ((_net_2214)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_944))?_add_all_x_data_out378:10'b0);
   assign  data_wire379 = ((_net_2213)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_943))?_add_all_x_data_out379:10'b0);
   assign  data_wire380 = ((_net_2212)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_942))?_add_all_x_data_out380:10'b0);
   assign  data_wire381 = ((_net_2211)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_941))?_add_all_x_data_out381:10'b0);
   assign  data_wire382 = ((_net_2210)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_940))?_add_all_x_data_out382:10'b0);
   assign  data_wire385 = ((_net_2209)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_939))?_add_all_x_data_out385:10'b0);
   assign  data_wire386 = ((_net_2208)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_938))?_add_all_x_data_out386:10'b0);
   assign  data_wire387 = ((_net_2207)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_937))?_add_all_x_data_out387:10'b0);
   assign  data_wire388 = ((_net_2206)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_936))?_add_all_x_data_out388:10'b0);
   assign  data_wire389 = ((_net_2205)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_935))?_add_all_x_data_out389:10'b0);
   assign  data_wire390 = ((_net_2204)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_934))?_add_all_x_data_out390:10'b0);
   assign  data_wire391 = ((_net_2203)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_933))?_add_all_x_data_out391:10'b0);
   assign  data_wire392 = ((_net_2202)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_932))?_add_all_x_data_out392:10'b0);
   assign  data_wire393 = ((_net_2201)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_931))?_add_all_x_data_out393:10'b0);
   assign  data_wire394 = ((_net_2200)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_930))?_add_all_x_data_out394:10'b0);
   assign  data_wire395 = ((_net_2199)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_929))?_add_all_x_data_out395:10'b0);
   assign  data_wire396 = ((_net_2198)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_928))?_add_all_x_data_out396:10'b0);
   assign  data_wire397 = ((_net_2197)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_927))?_add_all_x_data_out397:10'b0);
   assign  data_wire398 = ((_net_2196)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_926))?_add_all_x_data_out398:10'b0);
   assign  data_wire399 = ((_net_2195)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_925))?_add_all_x_data_out399:10'b0);
   assign  data_wire400 = ((_net_2194)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_924))?_add_all_x_data_out400:10'b0);
   assign  data_wire401 = ((_net_2193)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_923))?_add_all_x_data_out401:10'b0);
   assign  data_wire402 = ((_net_2192)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_922))?_add_all_x_data_out402:10'b0);
   assign  data_wire403 = ((_net_2191)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_921))?_add_all_x_data_out403:10'b0);
   assign  data_wire404 = ((_net_2190)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_920))?_add_all_x_data_out404:10'b0);
   assign  data_wire405 = ((_net_2189)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_919))?_add_all_x_data_out405:10'b0);
   assign  data_wire406 = ((_net_2188)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_918))?_add_all_x_data_out406:10'b0);
   assign  data_wire407 = ((_net_2187)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_917))?_add_all_x_data_out407:10'b0);
   assign  data_wire408 = ((_net_2186)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_916))?_add_all_x_data_out408:10'b0);
   assign  data_wire409 = ((_net_2185)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_915))?_add_all_x_data_out409:10'b0);
   assign  data_wire410 = ((_net_2184)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_914))?_add_all_x_data_out410:10'b0);
   assign  data_wire411 = ((_net_2183)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_913))?_add_all_x_data_out411:10'b0);
   assign  data_wire412 = ((_net_2182)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_912))?_add_all_x_data_out412:10'b0);
   assign  data_wire413 = ((_net_2181)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_911))?_add_all_x_data_out413:10'b0);
   assign  data_wire414 = ((_net_2180)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_910))?_add_all_x_data_out414:10'b0);
   assign  data_wire417 = ((_net_2179)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_909))?_add_all_x_data_out417:10'b0);
   assign  data_wire418 = ((_net_2178)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_908))?_add_all_x_data_out418:10'b0);
   assign  data_wire419 = ((_net_2177)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_907))?_add_all_x_data_out419:10'b0);
   assign  data_wire420 = ((_net_2176)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_906))?_add_all_x_data_out420:10'b0);
   assign  data_wire421 = ((_net_2175)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_905))?_add_all_x_data_out421:10'b0);
   assign  data_wire422 = ((_net_2174)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_904))?_add_all_x_data_out422:10'b0);
   assign  data_wire423 = ((_net_2173)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_903))?_add_all_x_data_out423:10'b0);
   assign  data_wire424 = ((_net_2172)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_902))?_add_all_x_data_out424:10'b0);
   assign  data_wire425 = ((_net_2171)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_901))?_add_all_x_data_out425:10'b0);
   assign  data_wire426 = ((_net_2170)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_900))?_add_all_x_data_out426:10'b0);
   assign  data_wire427 = ((_net_2169)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_899))?_add_all_x_data_out427:10'b0);
   assign  data_wire428 = ((_net_2168)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_898))?_add_all_x_data_out428:10'b0);
   assign  data_wire429 = ((_net_2167)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_897))?_add_all_x_data_out429:10'b0);
   assign  data_wire430 = ((_net_2166)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_896))?_add_all_x_data_out430:10'b0);
   assign  data_wire431 = ((_net_2165)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_895))?_add_all_x_data_out431:10'b0);
   assign  data_wire432 = ((_net_2164)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_894))?_add_all_x_data_out432:10'b0);
   assign  data_wire433 = ((_net_2163)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_893))?_add_all_x_data_out433:10'b0);
   assign  data_wire434 = ((_net_2162)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_892))?_add_all_x_data_out434:10'b0);
   assign  data_wire435 = ((_net_2161)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_891))?_add_all_x_data_out435:10'b0);
   assign  data_wire436 = ((_net_2160)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_890))?_add_all_x_data_out436:10'b0);
   assign  data_wire437 = ((_net_2159)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_889))?_add_all_x_data_out437:10'b0);
   assign  data_wire438 = ((_net_2158)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_888))?_add_all_x_data_out438:10'b0);
   assign  data_wire439 = ((_net_2157)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_887))?_add_all_x_data_out439:10'b0);
   assign  data_wire440 = ((_net_2156)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_886))?_add_all_x_data_out440:10'b0);
   assign  data_wire441 = ((_net_2155)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_885))?_add_all_x_data_out441:10'b0);
   assign  data_wire442 = ((_net_2154)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_884))?_add_all_x_data_out442:10'b0);
   assign  data_wire443 = ((_net_2153)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_883))?_add_all_x_data_out443:10'b0);
   assign  data_wire444 = ((_net_2152)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_882))?_add_all_x_data_out444:10'b0);
   assign  data_wire445 = ((_net_2151)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_881))?_add_all_x_data_out445:10'b0);
   assign  data_wire446 = ((_net_2150)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_880))?_add_all_x_data_out446:10'b0);
   assign  data_wire449 = ((_net_2149)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_879))?_add_all_x_data_out449:10'b0);
   assign  data_wire450 = ((_net_2148)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_878))?_add_all_x_data_out450:10'b0);
   assign  data_wire451 = ((_net_2147)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_877))?_add_all_x_data_out451:10'b0);
   assign  data_wire452 = ((_net_2146)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_876))?_add_all_x_data_out452:10'b0);
   assign  data_wire453 = ((_net_2145)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_875))?_add_all_x_data_out453:10'b0);
   assign  data_wire454 = ((_net_2144)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_874))?_add_all_x_data_out454:10'b0);
   assign  data_wire455 = ((_net_2143)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_873))?_add_all_x_data_out455:10'b0);
   assign  data_wire456 = ((_net_2142)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_872))?_add_all_x_data_out456:10'b0);
   assign  data_wire457 = ((_net_2141)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_871))?_add_all_x_data_out457:10'b0);
   assign  data_wire458 = ((_net_2140)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_870))?_add_all_x_data_out458:10'b0);
   assign  data_wire459 = ((_net_2139)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_869))?_add_all_x_data_out459:10'b0);
   assign  data_wire460 = ((_net_2138)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_868))?_add_all_x_data_out460:10'b0);
   assign  data_wire461 = ((_net_2137)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_867))?_add_all_x_data_out461:10'b0);
   assign  data_wire462 = ((_net_2136)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_866))?_add_all_x_data_out462:10'b0);
   assign  data_wire463 = ((_net_2135)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_865))?_add_all_x_data_out463:10'b0);
   assign  data_wire464 = ((_net_2134)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_864))?_add_all_x_data_out464:10'b0);
   assign  data_wire465 = ((_net_2133)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_863))?_add_all_x_data_out465:10'b0);
   assign  data_wire466 = ((_net_2132)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_862))?_add_all_x_data_out466:10'b0);
   assign  data_wire467 = ((_net_2131)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_861))?_add_all_x_data_out467:10'b0);
   assign  data_wire468 = ((_net_2130)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_860))?_add_all_x_data_out468:10'b0);
   assign  data_wire469 = ((_net_2129)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_859))?_add_all_x_data_out469:10'b0);
   assign  data_wire470 = ((_net_2128)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_858))?_add_all_x_data_out470:10'b0);
   assign  data_wire471 = ((_net_2127)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_857))?_add_all_x_data_out471:10'b0);
   assign  data_wire472 = ((_net_2126)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_856))?_add_all_x_data_out472:10'b0);
   assign  data_wire473 = ((_net_2125)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_855))?_add_all_x_data_out473:10'b0);
   assign  data_wire474 = ((_net_2124)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_854))?_add_all_x_data_out474:10'b0);
   assign  data_wire475 = ((_net_2123)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_853))?_add_all_x_data_out475:10'b0);
   assign  data_wire476 = ((_net_2122)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_852))?_add_all_x_data_out476:10'b0);
   assign  data_wire477 = ((_net_2121)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_851))?_add_all_x_data_out477:10'b0);
   assign  data_wire478 = ((_net_2120)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    (((_reg_2|_net_850))?_add_all_x_data_out478:10'b0);
   assign  data_out_org33 = ((_net_2119)?data_in33:10'b0)|
    (((_reg_2|_net_849))?_add_all_x_data_out_org33:10'b0);
   assign  data_out_org34 = ((_net_2118)?data_in34:10'b0)|
    (((_reg_2|_net_848))?_add_all_x_data_out_org34:10'b0);
   assign  data_out_org35 = ((_net_2117)?data_in35:10'b0)|
    (((_reg_2|_net_847))?_add_all_x_data_out_org35:10'b0);
   assign  data_out_org36 = ((_net_2116)?data_in36:10'b0)|
    (((_reg_2|_net_846))?_add_all_x_data_out_org36:10'b0);
   assign  data_out_org37 = ((_net_2115)?data_in37:10'b0)|
    (((_reg_2|_net_845))?_add_all_x_data_out_org37:10'b0);
   assign  data_out_org38 = ((_net_2114)?data_in38:10'b0)|
    (((_reg_2|_net_844))?_add_all_x_data_out_org38:10'b0);
   assign  data_out_org39 = ((_net_2113)?data_in39:10'b0)|
    (((_reg_2|_net_843))?_add_all_x_data_out_org39:10'b0);
   assign  data_out_org40 = ((_net_2112)?data_in40:10'b0)|
    (((_reg_2|_net_842))?_add_all_x_data_out_org40:10'b0);
   assign  data_out_org41 = ((_net_2111)?data_in41:10'b0)|
    (((_reg_2|_net_841))?_add_all_x_data_out_org41:10'b0);
   assign  data_out_org42 = ((_net_2110)?data_in42:10'b0)|
    (((_reg_2|_net_840))?_add_all_x_data_out_org42:10'b0);
   assign  data_out_org43 = ((_net_2109)?data_in43:10'b0)|
    (((_reg_2|_net_839))?_add_all_x_data_out_org43:10'b0);
   assign  data_out_org44 = ((_net_2108)?data_in44:10'b0)|
    (((_reg_2|_net_838))?_add_all_x_data_out_org44:10'b0);
   assign  data_out_org45 = ((_net_2107)?data_in45:10'b0)|
    (((_reg_2|_net_837))?_add_all_x_data_out_org45:10'b0);
   assign  data_out_org46 = ((_net_2106)?data_in46:10'b0)|
    (((_reg_2|_net_836))?_add_all_x_data_out_org46:10'b0);
   assign  data_out_org47 = ((_net_2105)?data_in47:10'b0)|
    (((_reg_2|_net_835))?_add_all_x_data_out_org47:10'b0);
   assign  data_out_org48 = ((_net_2104)?data_in48:10'b0)|
    (((_reg_2|_net_834))?_add_all_x_data_out_org48:10'b0);
   assign  data_out_org49 = ((_net_2103)?data_in49:10'b0)|
    (((_reg_2|_net_833))?_add_all_x_data_out_org49:10'b0);
   assign  data_out_org50 = ((_net_2102)?data_in50:10'b0)|
    (((_reg_2|_net_832))?_add_all_x_data_out_org50:10'b0);
   assign  data_out_org51 = ((_net_2101)?data_in51:10'b0)|
    (((_reg_2|_net_831))?_add_all_x_data_out_org51:10'b0);
   assign  data_out_org52 = ((_net_2100)?data_in52:10'b0)|
    (((_reg_2|_net_830))?_add_all_x_data_out_org52:10'b0);
   assign  data_out_org53 = ((_net_2099)?data_in53:10'b0)|
    (((_reg_2|_net_829))?_add_all_x_data_out_org53:10'b0);
   assign  data_out_org54 = ((_net_2098)?data_in54:10'b0)|
    (((_reg_2|_net_828))?_add_all_x_data_out_org54:10'b0);
   assign  data_out_org55 = ((_net_2097)?data_in55:10'b0)|
    (((_reg_2|_net_827))?_add_all_x_data_out_org55:10'b0);
   assign  data_out_org56 = ((_net_2096)?data_in56:10'b0)|
    (((_reg_2|_net_826))?_add_all_x_data_out_org56:10'b0);
   assign  data_out_org57 = ((_net_2095)?data_in57:10'b0)|
    (((_reg_2|_net_825))?_add_all_x_data_out_org57:10'b0);
   assign  data_out_org58 = ((_net_2094)?data_in58:10'b0)|
    (((_reg_2|_net_824))?_add_all_x_data_out_org58:10'b0);
   assign  data_out_org59 = ((_net_2093)?data_in59:10'b0)|
    (((_reg_2|_net_823))?_add_all_x_data_out_org59:10'b0);
   assign  data_out_org60 = ((_net_2092)?data_in60:10'b0)|
    (((_reg_2|_net_822))?_add_all_x_data_out_org60:10'b0);
   assign  data_out_org61 = ((_net_2091)?data_in61:10'b0)|
    (((_reg_2|_net_821))?_add_all_x_data_out_org61:10'b0);
   assign  data_out_org62 = ((_net_2090)?data_in62:10'b0)|
    (((_reg_2|_net_820))?_add_all_x_data_out_org62:10'b0);
   assign  data_out_org65 = ((_net_2089)?data_in65:10'b0)|
    (((_reg_2|_net_819))?_add_all_x_data_out_org65:10'b0);
   assign  data_out_org66 = ((_net_2088)?data_in66:10'b0)|
    (((_reg_2|_net_818))?_add_all_x_data_out_org66:10'b0);
   assign  data_out_org67 = ((_net_2087)?data_in67:10'b0)|
    (((_reg_2|_net_817))?_add_all_x_data_out_org67:10'b0);
   assign  data_out_org68 = ((_net_2086)?data_in68:10'b0)|
    (((_reg_2|_net_816))?_add_all_x_data_out_org68:10'b0);
   assign  data_out_org69 = ((_net_2085)?data_in69:10'b0)|
    (((_reg_2|_net_815))?_add_all_x_data_out_org69:10'b0);
   assign  data_out_org70 = ((_net_2084)?data_in70:10'b0)|
    (((_reg_2|_net_814))?_add_all_x_data_out_org70:10'b0);
   assign  data_out_org71 = ((_net_2083)?data_in71:10'b0)|
    (((_reg_2|_net_813))?_add_all_x_data_out_org71:10'b0);
   assign  data_out_org72 = ((_net_2082)?data_in72:10'b0)|
    (((_reg_2|_net_812))?_add_all_x_data_out_org72:10'b0);
   assign  data_out_org73 = ((_net_2081)?data_in73:10'b0)|
    (((_reg_2|_net_811))?_add_all_x_data_out_org73:10'b0);
   assign  data_out_org74 = ((_net_2080)?data_in74:10'b0)|
    (((_reg_2|_net_810))?_add_all_x_data_out_org74:10'b0);
   assign  data_out_org75 = ((_net_2079)?data_in75:10'b0)|
    (((_reg_2|_net_809))?_add_all_x_data_out_org75:10'b0);
   assign  data_out_org76 = ((_net_2078)?data_in76:10'b0)|
    (((_reg_2|_net_808))?_add_all_x_data_out_org76:10'b0);
   assign  data_out_org77 = ((_net_2077)?data_in77:10'b0)|
    (((_reg_2|_net_807))?_add_all_x_data_out_org77:10'b0);
   assign  data_out_org78 = ((_net_2076)?data_in78:10'b0)|
    (((_reg_2|_net_806))?_add_all_x_data_out_org78:10'b0);
   assign  data_out_org79 = ((_net_2075)?data_in79:10'b0)|
    (((_reg_2|_net_805))?_add_all_x_data_out_org79:10'b0);
   assign  data_out_org80 = ((_net_2074)?data_in80:10'b0)|
    (((_reg_2|_net_804))?_add_all_x_data_out_org80:10'b0);
   assign  data_out_org81 = ((_net_2073)?data_in81:10'b0)|
    (((_reg_2|_net_803))?_add_all_x_data_out_org81:10'b0);
   assign  data_out_org82 = ((_net_2072)?data_in82:10'b0)|
    (((_reg_2|_net_802))?_add_all_x_data_out_org82:10'b0);
   assign  data_out_org83 = ((_net_2071)?data_in83:10'b0)|
    (((_reg_2|_net_801))?_add_all_x_data_out_org83:10'b0);
   assign  data_out_org84 = ((_net_2070)?data_in84:10'b0)|
    (((_reg_2|_net_800))?_add_all_x_data_out_org84:10'b0);
   assign  data_out_org85 = ((_net_2069)?data_in85:10'b0)|
    (((_reg_2|_net_799))?_add_all_x_data_out_org85:10'b0);
   assign  data_out_org86 = ((_net_2068)?data_in86:10'b0)|
    (((_reg_2|_net_798))?_add_all_x_data_out_org86:10'b0);
   assign  data_out_org87 = ((_net_2067)?data_in87:10'b0)|
    (((_reg_2|_net_797))?_add_all_x_data_out_org87:10'b0);
   assign  data_out_org88 = ((_net_2066)?data_in88:10'b0)|
    (((_reg_2|_net_796))?_add_all_x_data_out_org88:10'b0);
   assign  data_out_org89 = ((_net_2065)?data_in89:10'b0)|
    (((_reg_2|_net_795))?_add_all_x_data_out_org89:10'b0);
   assign  data_out_org90 = ((_net_2064)?data_in90:10'b0)|
    (((_reg_2|_net_794))?_add_all_x_data_out_org90:10'b0);
   assign  data_out_org91 = ((_net_2063)?data_in91:10'b0)|
    (((_reg_2|_net_793))?_add_all_x_data_out_org91:10'b0);
   assign  data_out_org92 = ((_net_2062)?data_in92:10'b0)|
    (((_reg_2|_net_792))?_add_all_x_data_out_org92:10'b0);
   assign  data_out_org93 = ((_net_2061)?data_in93:10'b0)|
    (((_reg_2|_net_791))?_add_all_x_data_out_org93:10'b0);
   assign  data_out_org94 = ((_net_2060)?data_in94:10'b0)|
    (((_reg_2|_net_790))?_add_all_x_data_out_org94:10'b0);
   assign  data_out_org97 = ((_net_2059)?data_in97:10'b0)|
    (((_reg_2|_net_789))?_add_all_x_data_out_org97:10'b0);
   assign  data_out_org98 = ((_net_2058)?data_in98:10'b0)|
    (((_reg_2|_net_788))?_add_all_x_data_out_org98:10'b0);
   assign  data_out_org99 = ((_net_2057)?data_in99:10'b0)|
    (((_reg_2|_net_787))?_add_all_x_data_out_org99:10'b0);
   assign  data_out_org100 = ((_net_2056)?data_in100:10'b0)|
    (((_reg_2|_net_786))?_add_all_x_data_out_org100:10'b0);
   assign  data_out_org101 = ((_net_2055)?data_in101:10'b0)|
    (((_reg_2|_net_785))?_add_all_x_data_out_org101:10'b0);
   assign  data_out_org102 = ((_net_2054)?data_in102:10'b0)|
    (((_reg_2|_net_784))?_add_all_x_data_out_org102:10'b0);
   assign  data_out_org103 = ((_net_2053)?data_in103:10'b0)|
    (((_reg_2|_net_783))?_add_all_x_data_out_org103:10'b0);
   assign  data_out_org104 = ((_net_2052)?data_in104:10'b0)|
    (((_reg_2|_net_782))?_add_all_x_data_out_org104:10'b0);
   assign  data_out_org105 = ((_net_2051)?data_in105:10'b0)|
    (((_reg_2|_net_781))?_add_all_x_data_out_org105:10'b0);
   assign  data_out_org106 = ((_net_2050)?data_in106:10'b0)|
    (((_reg_2|_net_780))?_add_all_x_data_out_org106:10'b0);
   assign  data_out_org107 = ((_net_2049)?data_in107:10'b0)|
    (((_reg_2|_net_779))?_add_all_x_data_out_org107:10'b0);
   assign  data_out_org108 = ((_net_2048)?data_in108:10'b0)|
    (((_reg_2|_net_778))?_add_all_x_data_out_org108:10'b0);
   assign  data_out_org109 = ((_net_2047)?data_in109:10'b0)|
    (((_reg_2|_net_777))?_add_all_x_data_out_org109:10'b0);
   assign  data_out_org110 = ((_net_2046)?data_in110:10'b0)|
    (((_reg_2|_net_776))?_add_all_x_data_out_org110:10'b0);
   assign  data_out_org111 = ((_net_2045)?data_in111:10'b0)|
    (((_reg_2|_net_775))?_add_all_x_data_out_org111:10'b0);
   assign  data_out_org112 = ((_net_2044)?data_in112:10'b0)|
    (((_reg_2|_net_774))?_add_all_x_data_out_org112:10'b0);
   assign  data_out_org113 = ((_net_2043)?data_in113:10'b0)|
    (((_reg_2|_net_773))?_add_all_x_data_out_org113:10'b0);
   assign  data_out_org114 = ((_net_2042)?data_in114:10'b0)|
    (((_reg_2|_net_772))?_add_all_x_data_out_org114:10'b0);
   assign  data_out_org115 = ((_net_2041)?data_in115:10'b0)|
    (((_reg_2|_net_771))?_add_all_x_data_out_org115:10'b0);
   assign  data_out_org116 = ((_net_2040)?data_in116:10'b0)|
    (((_reg_2|_net_770))?_add_all_x_data_out_org116:10'b0);
   assign  data_out_org117 = ((_net_2039)?data_in117:10'b0)|
    (((_reg_2|_net_769))?_add_all_x_data_out_org117:10'b0);
   assign  data_out_org118 = ((_net_2038)?data_in118:10'b0)|
    (((_reg_2|_net_768))?_add_all_x_data_out_org118:10'b0);
   assign  data_out_org119 = ((_net_2037)?data_in119:10'b0)|
    (((_reg_2|_net_767))?_add_all_x_data_out_org119:10'b0);
   assign  data_out_org120 = ((_net_2036)?data_in120:10'b0)|
    (((_reg_2|_net_766))?_add_all_x_data_out_org120:10'b0);
   assign  data_out_org121 = ((_net_2035)?data_in121:10'b0)|
    (((_reg_2|_net_765))?_add_all_x_data_out_org121:10'b0);
   assign  data_out_org122 = ((_net_2034)?data_in122:10'b0)|
    (((_reg_2|_net_764))?_add_all_x_data_out_org122:10'b0);
   assign  data_out_org123 = ((_net_2033)?data_in123:10'b0)|
    (((_reg_2|_net_763))?_add_all_x_data_out_org123:10'b0);
   assign  data_out_org124 = ((_net_2032)?data_in124:10'b0)|
    (((_reg_2|_net_762))?_add_all_x_data_out_org124:10'b0);
   assign  data_out_org125 = ((_net_2031)?data_in125:10'b0)|
    (((_reg_2|_net_761))?_add_all_x_data_out_org125:10'b0);
   assign  data_out_org126 = ((_net_2030)?data_in126:10'b0)|
    (((_reg_2|_net_760))?_add_all_x_data_out_org126:10'b0);
   assign  data_out_org129 = ((_net_2029)?data_in129:10'b0)|
    (((_reg_2|_net_759))?_add_all_x_data_out_org129:10'b0);
   assign  data_out_org130 = ((_net_2028)?data_in130:10'b0)|
    (((_reg_2|_net_758))?_add_all_x_data_out_org130:10'b0);
   assign  data_out_org131 = ((_net_2027)?data_in131:10'b0)|
    (((_reg_2|_net_757))?_add_all_x_data_out_org131:10'b0);
   assign  data_out_org132 = ((_net_2026)?data_in132:10'b0)|
    (((_reg_2|_net_756))?_add_all_x_data_out_org132:10'b0);
   assign  data_out_org133 = ((_net_2025)?data_in133:10'b0)|
    (((_reg_2|_net_755))?_add_all_x_data_out_org133:10'b0);
   assign  data_out_org134 = ((_net_2024)?data_in134:10'b0)|
    (((_reg_2|_net_754))?_add_all_x_data_out_org134:10'b0);
   assign  data_out_org135 = ((_net_2023)?data_in135:10'b0)|
    (((_reg_2|_net_753))?_add_all_x_data_out_org135:10'b0);
   assign  data_out_org136 = ((_net_2022)?data_in136:10'b0)|
    (((_reg_2|_net_752))?_add_all_x_data_out_org136:10'b0);
   assign  data_out_org137 = ((_net_2021)?data_in137:10'b0)|
    (((_reg_2|_net_751))?_add_all_x_data_out_org137:10'b0);
   assign  data_out_org138 = ((_net_2020)?data_in138:10'b0)|
    (((_reg_2|_net_750))?_add_all_x_data_out_org138:10'b0);
   assign  data_out_org139 = ((_net_2019)?data_in139:10'b0)|
    (((_reg_2|_net_749))?_add_all_x_data_out_org139:10'b0);
   assign  data_out_org140 = ((_net_2018)?data_in140:10'b0)|
    (((_reg_2|_net_748))?_add_all_x_data_out_org140:10'b0);
   assign  data_out_org141 = ((_net_2017)?data_in141:10'b0)|
    (((_reg_2|_net_747))?_add_all_x_data_out_org141:10'b0);
   assign  data_out_org142 = ((_net_2016)?data_in142:10'b0)|
    (((_reg_2|_net_746))?_add_all_x_data_out_org142:10'b0);
   assign  data_out_org143 = ((_net_2015)?data_in143:10'b0)|
    (((_reg_2|_net_745))?_add_all_x_data_out_org143:10'b0);
   assign  data_out_org144 = ((_net_2014)?data_in144:10'b0)|
    (((_reg_2|_net_744))?_add_all_x_data_out_org144:10'b0);
   assign  data_out_org145 = ((_net_2013)?data_in145:10'b0)|
    (((_reg_2|_net_743))?_add_all_x_data_out_org145:10'b0);
   assign  data_out_org146 = ((_net_2012)?data_in146:10'b0)|
    (((_reg_2|_net_742))?_add_all_x_data_out_org146:10'b0);
   assign  data_out_org147 = ((_net_2011)?data_in147:10'b0)|
    (((_reg_2|_net_741))?_add_all_x_data_out_org147:10'b0);
   assign  data_out_org148 = ((_net_2010)?data_in148:10'b0)|
    (((_reg_2|_net_740))?_add_all_x_data_out_org148:10'b0);
   assign  data_out_org149 = ((_net_2009)?data_in149:10'b0)|
    (((_reg_2|_net_739))?_add_all_x_data_out_org149:10'b0);
   assign  data_out_org150 = ((_net_2008)?data_in150:10'b0)|
    (((_reg_2|_net_738))?_add_all_x_data_out_org150:10'b0);
   assign  data_out_org151 = ((_net_2007)?data_in151:10'b0)|
    (((_reg_2|_net_737))?_add_all_x_data_out_org151:10'b0);
   assign  data_out_org152 = ((_net_2006)?data_in152:10'b0)|
    (((_reg_2|_net_736))?_add_all_x_data_out_org152:10'b0);
   assign  data_out_org153 = ((_net_2005)?data_in153:10'b0)|
    (((_reg_2|_net_735))?_add_all_x_data_out_org153:10'b0);
   assign  data_out_org154 = ((_net_2004)?data_in154:10'b0)|
    (((_reg_2|_net_734))?_add_all_x_data_out_org154:10'b0);
   assign  data_out_org155 = ((_net_2003)?data_in155:10'b0)|
    (((_reg_2|_net_733))?_add_all_x_data_out_org155:10'b0);
   assign  data_out_org156 = ((_net_2002)?data_in156:10'b0)|
    (((_reg_2|_net_732))?_add_all_x_data_out_org156:10'b0);
   assign  data_out_org157 = ((_net_2001)?data_in157:10'b0)|
    (((_reg_2|_net_731))?_add_all_x_data_out_org157:10'b0);
   assign  data_out_org158 = ((_net_2000)?data_in158:10'b0)|
    (((_reg_2|_net_730))?_add_all_x_data_out_org158:10'b0);
   assign  data_out_org161 = ((_net_1999)?data_in161:10'b0)|
    (((_reg_2|_net_729))?_add_all_x_data_out_org161:10'b0);
   assign  data_out_org162 = ((_net_1998)?data_in162:10'b0)|
    (((_reg_2|_net_728))?_add_all_x_data_out_org162:10'b0);
   assign  data_out_org163 = ((_net_1997)?data_in163:10'b0)|
    (((_reg_2|_net_727))?_add_all_x_data_out_org163:10'b0);
   assign  data_out_org164 = ((_net_1996)?data_in164:10'b0)|
    (((_reg_2|_net_726))?_add_all_x_data_out_org164:10'b0);
   assign  data_out_org165 = ((_net_1995)?data_in165:10'b0)|
    (((_reg_2|_net_725))?_add_all_x_data_out_org165:10'b0);
   assign  data_out_org166 = ((_net_1994)?data_in166:10'b0)|
    (((_reg_2|_net_724))?_add_all_x_data_out_org166:10'b0);
   assign  data_out_org167 = ((_net_1993)?data_in167:10'b0)|
    (((_reg_2|_net_723))?_add_all_x_data_out_org167:10'b0);
   assign  data_out_org168 = ((_net_1992)?data_in168:10'b0)|
    (((_reg_2|_net_722))?_add_all_x_data_out_org168:10'b0);
   assign  data_out_org169 = ((_net_1991)?data_in169:10'b0)|
    (((_reg_2|_net_721))?_add_all_x_data_out_org169:10'b0);
   assign  data_out_org170 = ((_net_1990)?data_in170:10'b0)|
    (((_reg_2|_net_720))?_add_all_x_data_out_org170:10'b0);
   assign  data_out_org171 = ((_net_1989)?data_in171:10'b0)|
    (((_reg_2|_net_719))?_add_all_x_data_out_org171:10'b0);
   assign  data_out_org172 = ((_net_1988)?data_in172:10'b0)|
    (((_reg_2|_net_718))?_add_all_x_data_out_org172:10'b0);
   assign  data_out_org173 = ((_net_1987)?data_in173:10'b0)|
    (((_reg_2|_net_717))?_add_all_x_data_out_org173:10'b0);
   assign  data_out_org174 = ((_net_1986)?data_in174:10'b0)|
    (((_reg_2|_net_716))?_add_all_x_data_out_org174:10'b0);
   assign  data_out_org175 = ((_net_1985)?data_in175:10'b0)|
    (((_reg_2|_net_715))?_add_all_x_data_out_org175:10'b0);
   assign  data_out_org176 = ((_net_1984)?data_in176:10'b0)|
    (((_reg_2|_net_714))?_add_all_x_data_out_org176:10'b0);
   assign  data_out_org177 = ((_net_1983)?data_in177:10'b0)|
    (((_reg_2|_net_713))?_add_all_x_data_out_org177:10'b0);
   assign  data_out_org178 = ((_net_1982)?data_in178:10'b0)|
    (((_reg_2|_net_712))?_add_all_x_data_out_org178:10'b0);
   assign  data_out_org179 = ((_net_1981)?data_in179:10'b0)|
    (((_reg_2|_net_711))?_add_all_x_data_out_org179:10'b0);
   assign  data_out_org180 = ((_net_1980)?data_in180:10'b0)|
    (((_reg_2|_net_710))?_add_all_x_data_out_org180:10'b0);
   assign  data_out_org181 = ((_net_1979)?data_in181:10'b0)|
    (((_reg_2|_net_709))?_add_all_x_data_out_org181:10'b0);
   assign  data_out_org182 = ((_net_1978)?data_in182:10'b0)|
    (((_reg_2|_net_708))?_add_all_x_data_out_org182:10'b0);
   assign  data_out_org183 = ((_net_1977)?data_in183:10'b0)|
    (((_reg_2|_net_707))?_add_all_x_data_out_org183:10'b0);
   assign  data_out_org184 = ((_net_1976)?data_in184:10'b0)|
    (((_reg_2|_net_706))?_add_all_x_data_out_org184:10'b0);
   assign  data_out_org185 = ((_net_1975)?data_in185:10'b0)|
    (((_reg_2|_net_705))?_add_all_x_data_out_org185:10'b0);
   assign  data_out_org186 = ((_net_1974)?data_in186:10'b0)|
    (((_reg_2|_net_704))?_add_all_x_data_out_org186:10'b0);
   assign  data_out_org187 = ((_net_1973)?data_in187:10'b0)|
    (((_reg_2|_net_703))?_add_all_x_data_out_org187:10'b0);
   assign  data_out_org188 = ((_net_1972)?data_in188:10'b0)|
    (((_reg_2|_net_702))?_add_all_x_data_out_org188:10'b0);
   assign  data_out_org189 = ((_net_1971)?data_in189:10'b0)|
    (((_reg_2|_net_701))?_add_all_x_data_out_org189:10'b0);
   assign  data_out_org190 = ((_net_1970)?data_in190:10'b0)|
    (((_reg_2|_net_700))?_add_all_x_data_out_org190:10'b0);
   assign  data_out_org193 = ((_net_1969)?data_in193:10'b0)|
    (((_reg_2|_net_699))?_add_all_x_data_out_org193:10'b0);
   assign  data_out_org194 = ((_net_1968)?data_in194:10'b0)|
    (((_reg_2|_net_698))?_add_all_x_data_out_org194:10'b0);
   assign  data_out_org195 = ((_net_1967)?data_in195:10'b0)|
    (((_reg_2|_net_697))?_add_all_x_data_out_org195:10'b0);
   assign  data_out_org196 = ((_net_1966)?data_in196:10'b0)|
    (((_reg_2|_net_696))?_add_all_x_data_out_org196:10'b0);
   assign  data_out_org197 = ((_net_1965)?data_in197:10'b0)|
    (((_reg_2|_net_695))?_add_all_x_data_out_org197:10'b0);
   assign  data_out_org198 = ((_net_1964)?data_in198:10'b0)|
    (((_reg_2|_net_694))?_add_all_x_data_out_org198:10'b0);
   assign  data_out_org199 = ((_net_1963)?data_in199:10'b0)|
    (((_reg_2|_net_693))?_add_all_x_data_out_org199:10'b0);
   assign  data_out_org200 = ((_net_1962)?data_in200:10'b0)|
    (((_reg_2|_net_692))?_add_all_x_data_out_org200:10'b0);
   assign  data_out_org201 = ((_net_1961)?data_in201:10'b0)|
    (((_reg_2|_net_691))?_add_all_x_data_out_org201:10'b0);
   assign  data_out_org202 = ((_net_1960)?data_in202:10'b0)|
    (((_reg_2|_net_690))?_add_all_x_data_out_org202:10'b0);
   assign  data_out_org203 = ((_net_1959)?data_in203:10'b0)|
    (((_reg_2|_net_689))?_add_all_x_data_out_org203:10'b0);
   assign  data_out_org204 = ((_net_1958)?data_in204:10'b0)|
    (((_reg_2|_net_688))?_add_all_x_data_out_org204:10'b0);
   assign  data_out_org205 = ((_net_1957)?data_in205:10'b0)|
    (((_reg_2|_net_687))?_add_all_x_data_out_org205:10'b0);
   assign  data_out_org206 = ((_net_1956)?data_in206:10'b0)|
    (((_reg_2|_net_686))?_add_all_x_data_out_org206:10'b0);
   assign  data_out_org207 = ((_net_1955)?data_in207:10'b0)|
    (((_reg_2|_net_685))?_add_all_x_data_out_org207:10'b0);
   assign  data_out_org208 = ((_net_1954)?data_in208:10'b0)|
    (((_reg_2|_net_684))?_add_all_x_data_out_org208:10'b0);
   assign  data_out_org209 = ((_net_1953)?data_in209:10'b0)|
    (((_reg_2|_net_683))?_add_all_x_data_out_org209:10'b0);
   assign  data_out_org210 = ((_net_1952)?data_in210:10'b0)|
    (((_reg_2|_net_682))?_add_all_x_data_out_org210:10'b0);
   assign  data_out_org211 = ((_net_1951)?data_in211:10'b0)|
    (((_reg_2|_net_681))?_add_all_x_data_out_org211:10'b0);
   assign  data_out_org212 = ((_net_1950)?data_in212:10'b0)|
    (((_reg_2|_net_680))?_add_all_x_data_out_org212:10'b0);
   assign  data_out_org213 = ((_net_1949)?data_in213:10'b0)|
    (((_reg_2|_net_679))?_add_all_x_data_out_org213:10'b0);
   assign  data_out_org214 = ((_net_1948)?data_in214:10'b0)|
    (((_reg_2|_net_678))?_add_all_x_data_out_org214:10'b0);
   assign  data_out_org215 = ((_net_1947)?data_in215:10'b0)|
    (((_reg_2|_net_677))?_add_all_x_data_out_org215:10'b0);
   assign  data_out_org216 = ((_net_1946)?data_in216:10'b0)|
    (((_reg_2|_net_676))?_add_all_x_data_out_org216:10'b0);
   assign  data_out_org217 = ((_net_1945)?data_in217:10'b0)|
    (((_reg_2|_net_675))?_add_all_x_data_out_org217:10'b0);
   assign  data_out_org218 = ((_net_1944)?data_in218:10'b0)|
    (((_reg_2|_net_674))?_add_all_x_data_out_org218:10'b0);
   assign  data_out_org219 = ((_net_1943)?data_in219:10'b0)|
    (((_reg_2|_net_673))?_add_all_x_data_out_org219:10'b0);
   assign  data_out_org220 = ((_net_1942)?data_in220:10'b0)|
    (((_reg_2|_net_672))?_add_all_x_data_out_org220:10'b0);
   assign  data_out_org221 = ((_net_1941)?data_in221:10'b0)|
    (((_reg_2|_net_671))?_add_all_x_data_out_org221:10'b0);
   assign  data_out_org222 = ((_net_1940)?data_in222:10'b0)|
    (((_reg_2|_net_670))?_add_all_x_data_out_org222:10'b0);
   assign  data_out_org225 = ((_net_1939)?data_in225:10'b0)|
    (((_reg_2|_net_669))?_add_all_x_data_out_org225:10'b0);
   assign  data_out_org226 = ((_net_1938)?data_in226:10'b0)|
    (((_reg_2|_net_668))?_add_all_x_data_out_org226:10'b0);
   assign  data_out_org227 = ((_net_1937)?data_in227:10'b0)|
    (((_reg_2|_net_667))?_add_all_x_data_out_org227:10'b0);
   assign  data_out_org228 = ((_net_1936)?data_in228:10'b0)|
    (((_reg_2|_net_666))?_add_all_x_data_out_org228:10'b0);
   assign  data_out_org229 = ((_net_1935)?data_in229:10'b0)|
    (((_reg_2|_net_665))?_add_all_x_data_out_org229:10'b0);
   assign  data_out_org230 = ((_net_1934)?data_in230:10'b0)|
    (((_reg_2|_net_664))?_add_all_x_data_out_org230:10'b0);
   assign  data_out_org231 = ((_net_1933)?data_in231:10'b0)|
    (((_reg_2|_net_663))?_add_all_x_data_out_org231:10'b0);
   assign  data_out_org232 = ((_net_1932)?data_in232:10'b0)|
    (((_reg_2|_net_662))?_add_all_x_data_out_org232:10'b0);
   assign  data_out_org233 = ((_net_1931)?data_in233:10'b0)|
    (((_reg_2|_net_661))?_add_all_x_data_out_org233:10'b0);
   assign  data_out_org234 = ((_net_1930)?data_in234:10'b0)|
    (((_reg_2|_net_660))?_add_all_x_data_out_org234:10'b0);
   assign  data_out_org235 = ((_net_1929)?data_in235:10'b0)|
    (((_reg_2|_net_659))?_add_all_x_data_out_org235:10'b0);
   assign  data_out_org236 = ((_net_1928)?data_in236:10'b0)|
    (((_reg_2|_net_658))?_add_all_x_data_out_org236:10'b0);
   assign  data_out_org237 = ((_net_1927)?data_in237:10'b0)|
    (((_reg_2|_net_657))?_add_all_x_data_out_org237:10'b0);
   assign  data_out_org238 = ((_net_1926)?data_in238:10'b0)|
    (((_reg_2|_net_656))?_add_all_x_data_out_org238:10'b0);
   assign  data_out_org239 = ((_net_1925)?data_in239:10'b0)|
    (((_reg_2|_net_655))?_add_all_x_data_out_org239:10'b0);
   assign  data_out_org240 = ((_net_1924)?data_in240:10'b0)|
    (((_reg_2|_net_654))?_add_all_x_data_out_org240:10'b0);
   assign  data_out_org241 = ((_net_1923)?data_in241:10'b0)|
    (((_reg_2|_net_653))?_add_all_x_data_out_org241:10'b0);
   assign  data_out_org242 = ((_net_1922)?data_in242:10'b0)|
    (((_reg_2|_net_652))?_add_all_x_data_out_org242:10'b0);
   assign  data_out_org243 = ((_net_1921)?data_in243:10'b0)|
    (((_reg_2|_net_651))?_add_all_x_data_out_org243:10'b0);
   assign  data_out_org244 = ((_net_1920)?data_in244:10'b0)|
    (((_reg_2|_net_650))?_add_all_x_data_out_org244:10'b0);
   assign  data_out_org245 = ((_net_1919)?data_in245:10'b0)|
    (((_reg_2|_net_649))?_add_all_x_data_out_org245:10'b0);
   assign  data_out_org246 = ((_net_1918)?data_in246:10'b0)|
    (((_reg_2|_net_648))?_add_all_x_data_out_org246:10'b0);
   assign  data_out_org247 = ((_net_1917)?data_in247:10'b0)|
    (((_reg_2|_net_647))?_add_all_x_data_out_org247:10'b0);
   assign  data_out_org248 = ((_net_1916)?data_in248:10'b0)|
    (((_reg_2|_net_646))?_add_all_x_data_out_org248:10'b0);
   assign  data_out_org249 = ((_net_1915)?data_in249:10'b0)|
    (((_reg_2|_net_645))?_add_all_x_data_out_org249:10'b0);
   assign  data_out_org250 = ((_net_1914)?data_in250:10'b0)|
    (((_reg_2|_net_644))?_add_all_x_data_out_org250:10'b0);
   assign  data_out_org251 = ((_net_1913)?data_in251:10'b0)|
    (((_reg_2|_net_643))?_add_all_x_data_out_org251:10'b0);
   assign  data_out_org252 = ((_net_1912)?data_in252:10'b0)|
    (((_reg_2|_net_642))?_add_all_x_data_out_org252:10'b0);
   assign  data_out_org253 = ((_net_1911)?data_in253:10'b0)|
    (((_reg_2|_net_641))?_add_all_x_data_out_org253:10'b0);
   assign  data_out_org254 = ((_net_1910)?data_in254:10'b0)|
    (((_reg_2|_net_640))?_add_all_x_data_out_org254:10'b0);
   assign  data_out_org257 = ((_net_1909)?data_in257:10'b0)|
    (((_reg_2|_net_639))?_add_all_x_data_out_org257:10'b0);
   assign  data_out_org258 = ((_net_1908)?data_in258:10'b0)|
    (((_reg_2|_net_638))?_add_all_x_data_out_org258:10'b0);
   assign  data_out_org259 = ((_net_1907)?data_in259:10'b0)|
    (((_reg_2|_net_637))?_add_all_x_data_out_org259:10'b0);
   assign  data_out_org260 = ((_net_1906)?data_in260:10'b0)|
    (((_reg_2|_net_636))?_add_all_x_data_out_org260:10'b0);
   assign  data_out_org261 = ((_net_1905)?data_in261:10'b0)|
    (((_reg_2|_net_635))?_add_all_x_data_out_org261:10'b0);
   assign  data_out_org262 = ((_net_1904)?data_in262:10'b0)|
    (((_reg_2|_net_634))?_add_all_x_data_out_org262:10'b0);
   assign  data_out_org263 = ((_net_1903)?data_in263:10'b0)|
    (((_reg_2|_net_633))?_add_all_x_data_out_org263:10'b0);
   assign  data_out_org264 = ((_net_1902)?data_in264:10'b0)|
    (((_reg_2|_net_632))?_add_all_x_data_out_org264:10'b0);
   assign  data_out_org265 = ((_net_1901)?data_in265:10'b0)|
    (((_reg_2|_net_631))?_add_all_x_data_out_org265:10'b0);
   assign  data_out_org266 = ((_net_1900)?data_in266:10'b0)|
    (((_reg_2|_net_630))?_add_all_x_data_out_org266:10'b0);
   assign  data_out_org267 = ((_net_1899)?data_in267:10'b0)|
    (((_reg_2|_net_629))?_add_all_x_data_out_org267:10'b0);
   assign  data_out_org268 = ((_net_1898)?data_in268:10'b0)|
    (((_reg_2|_net_628))?_add_all_x_data_out_org268:10'b0);
   assign  data_out_org269 = ((_net_1897)?data_in269:10'b0)|
    (((_reg_2|_net_627))?_add_all_x_data_out_org269:10'b0);
   assign  data_out_org270 = ((_net_1896)?data_in270:10'b0)|
    (((_reg_2|_net_626))?_add_all_x_data_out_org270:10'b0);
   assign  data_out_org271 = ((_net_1895)?data_in271:10'b0)|
    (((_reg_2|_net_625))?_add_all_x_data_out_org271:10'b0);
   assign  data_out_org272 = ((_net_1894)?data_in272:10'b0)|
    (((_reg_2|_net_624))?_add_all_x_data_out_org272:10'b0);
   assign  data_out_org273 = ((_net_1893)?data_in273:10'b0)|
    (((_reg_2|_net_623))?_add_all_x_data_out_org273:10'b0);
   assign  data_out_org274 = ((_net_1892)?data_in274:10'b0)|
    (((_reg_2|_net_622))?_add_all_x_data_out_org274:10'b0);
   assign  data_out_org275 = ((_net_1891)?data_in275:10'b0)|
    (((_reg_2|_net_621))?_add_all_x_data_out_org275:10'b0);
   assign  data_out_org276 = ((_net_1890)?data_in276:10'b0)|
    (((_reg_2|_net_620))?_add_all_x_data_out_org276:10'b0);
   assign  data_out_org277 = ((_net_1889)?data_in277:10'b0)|
    (((_reg_2|_net_619))?_add_all_x_data_out_org277:10'b0);
   assign  data_out_org278 = ((_net_1888)?data_in278:10'b0)|
    (((_reg_2|_net_618))?_add_all_x_data_out_org278:10'b0);
   assign  data_out_org279 = ((_net_1887)?data_in279:10'b0)|
    (((_reg_2|_net_617))?_add_all_x_data_out_org279:10'b0);
   assign  data_out_org280 = ((_net_1886)?data_in280:10'b0)|
    (((_reg_2|_net_616))?_add_all_x_data_out_org280:10'b0);
   assign  data_out_org281 = ((_net_1885)?data_in281:10'b0)|
    (((_reg_2|_net_615))?_add_all_x_data_out_org281:10'b0);
   assign  data_out_org282 = ((_net_1884)?data_in282:10'b0)|
    (((_reg_2|_net_614))?_add_all_x_data_out_org282:10'b0);
   assign  data_out_org283 = ((_net_1883)?data_in283:10'b0)|
    (((_reg_2|_net_613))?_add_all_x_data_out_org283:10'b0);
   assign  data_out_org284 = ((_net_1882)?data_in284:10'b0)|
    (((_reg_2|_net_612))?_add_all_x_data_out_org284:10'b0);
   assign  data_out_org285 = ((_net_1881)?data_in285:10'b0)|
    (((_reg_2|_net_611))?_add_all_x_data_out_org285:10'b0);
   assign  data_out_org286 = ((_net_1880)?data_in286:10'b0)|
    (((_reg_2|_net_610))?_add_all_x_data_out_org286:10'b0);
   assign  data_out_org289 = ((_net_1879)?data_in289:10'b0)|
    (((_reg_2|_net_609))?_add_all_x_data_out_org289:10'b0);
   assign  data_out_org290 = ((_net_1878)?data_in290:10'b0)|
    (((_reg_2|_net_608))?_add_all_x_data_out_org290:10'b0);
   assign  data_out_org291 = ((_net_1877)?data_in291:10'b0)|
    (((_reg_2|_net_607))?_add_all_x_data_out_org291:10'b0);
   assign  data_out_org292 = ((_net_1876)?data_in292:10'b0)|
    (((_reg_2|_net_606))?_add_all_x_data_out_org292:10'b0);
   assign  data_out_org293 = ((_net_1875)?data_in293:10'b0)|
    (((_reg_2|_net_605))?_add_all_x_data_out_org293:10'b0);
   assign  data_out_org294 = ((_net_1874)?data_in294:10'b0)|
    (((_reg_2|_net_604))?_add_all_x_data_out_org294:10'b0);
   assign  data_out_org295 = ((_net_1873)?data_in295:10'b0)|
    (((_reg_2|_net_603))?_add_all_x_data_out_org295:10'b0);
   assign  data_out_org296 = ((_net_1872)?data_in296:10'b0)|
    (((_reg_2|_net_602))?_add_all_x_data_out_org296:10'b0);
   assign  data_out_org297 = ((_net_1871)?data_in297:10'b0)|
    (((_reg_2|_net_601))?_add_all_x_data_out_org297:10'b0);
   assign  data_out_org298 = ((_net_1870)?data_in298:10'b0)|
    (((_reg_2|_net_600))?_add_all_x_data_out_org298:10'b0);
   assign  data_out_org299 = ((_net_1869)?data_in299:10'b0)|
    (((_reg_2|_net_599))?_add_all_x_data_out_org299:10'b0);
   assign  data_out_org300 = ((_net_1868)?data_in300:10'b0)|
    (((_reg_2|_net_598))?_add_all_x_data_out_org300:10'b0);
   assign  data_out_org301 = ((_net_1867)?data_in301:10'b0)|
    (((_reg_2|_net_597))?_add_all_x_data_out_org301:10'b0);
   assign  data_out_org302 = ((_net_1866)?data_in302:10'b0)|
    (((_reg_2|_net_596))?_add_all_x_data_out_org302:10'b0);
   assign  data_out_org303 = ((_net_1865)?data_in303:10'b0)|
    (((_reg_2|_net_595))?_add_all_x_data_out_org303:10'b0);
   assign  data_out_org304 = ((_net_1864)?data_in304:10'b0)|
    (((_reg_2|_net_594))?_add_all_x_data_out_org304:10'b0);
   assign  data_out_org305 = ((_net_1863)?data_in305:10'b0)|
    (((_reg_2|_net_593))?_add_all_x_data_out_org305:10'b0);
   assign  data_out_org306 = ((_net_1862)?data_in306:10'b0)|
    (((_reg_2|_net_592))?_add_all_x_data_out_org306:10'b0);
   assign  data_out_org307 = ((_net_1861)?data_in307:10'b0)|
    (((_reg_2|_net_591))?_add_all_x_data_out_org307:10'b0);
   assign  data_out_org308 = ((_net_1860)?data_in308:10'b0)|
    (((_reg_2|_net_590))?_add_all_x_data_out_org308:10'b0);
   assign  data_out_org309 = ((_net_1859)?data_in309:10'b0)|
    (((_reg_2|_net_589))?_add_all_x_data_out_org309:10'b0);
   assign  data_out_org310 = ((_net_1858)?data_in310:10'b0)|
    (((_reg_2|_net_588))?_add_all_x_data_out_org310:10'b0);
   assign  data_out_org311 = ((_net_1857)?data_in311:10'b0)|
    (((_reg_2|_net_587))?_add_all_x_data_out_org311:10'b0);
   assign  data_out_org312 = ((_net_1856)?data_in312:10'b0)|
    (((_reg_2|_net_586))?_add_all_x_data_out_org312:10'b0);
   assign  data_out_org313 = ((_net_1855)?data_in313:10'b0)|
    (((_reg_2|_net_585))?_add_all_x_data_out_org313:10'b0);
   assign  data_out_org314 = ((_net_1854)?data_in314:10'b0)|
    (((_reg_2|_net_584))?_add_all_x_data_out_org314:10'b0);
   assign  data_out_org315 = ((_net_1853)?data_in315:10'b0)|
    (((_reg_2|_net_583))?_add_all_x_data_out_org315:10'b0);
   assign  data_out_org316 = ((_net_1852)?data_in316:10'b0)|
    (((_reg_2|_net_582))?_add_all_x_data_out_org316:10'b0);
   assign  data_out_org317 = ((_net_1851)?data_in317:10'b0)|
    (((_reg_2|_net_581))?_add_all_x_data_out_org317:10'b0);
   assign  data_out_org318 = ((_net_1850)?data_in318:10'b0)|
    (((_reg_2|_net_580))?_add_all_x_data_out_org318:10'b0);
   assign  data_out_org321 = ((_net_1849)?data_in321:10'b0)|
    (((_reg_2|_net_579))?_add_all_x_data_out_org321:10'b0);
   assign  data_out_org322 = ((_net_1848)?data_in322:10'b0)|
    (((_reg_2|_net_578))?_add_all_x_data_out_org322:10'b0);
   assign  data_out_org323 = ((_net_1847)?data_in323:10'b0)|
    (((_reg_2|_net_577))?_add_all_x_data_out_org323:10'b0);
   assign  data_out_org324 = ((_net_1846)?data_in324:10'b0)|
    (((_reg_2|_net_576))?_add_all_x_data_out_org324:10'b0);
   assign  data_out_org325 = ((_net_1845)?data_in325:10'b0)|
    (((_reg_2|_net_575))?_add_all_x_data_out_org325:10'b0);
   assign  data_out_org326 = ((_net_1844)?data_in326:10'b0)|
    (((_reg_2|_net_574))?_add_all_x_data_out_org326:10'b0);
   assign  data_out_org327 = ((_net_1843)?data_in327:10'b0)|
    (((_reg_2|_net_573))?_add_all_x_data_out_org327:10'b0);
   assign  data_out_org328 = ((_net_1842)?data_in328:10'b0)|
    (((_reg_2|_net_572))?_add_all_x_data_out_org328:10'b0);
   assign  data_out_org329 = ((_net_1841)?data_in329:10'b0)|
    (((_reg_2|_net_571))?_add_all_x_data_out_org329:10'b0);
   assign  data_out_org330 = ((_net_1840)?data_in330:10'b0)|
    (((_reg_2|_net_570))?_add_all_x_data_out_org330:10'b0);
   assign  data_out_org331 = ((_net_1839)?data_in331:10'b0)|
    (((_reg_2|_net_569))?_add_all_x_data_out_org331:10'b0);
   assign  data_out_org332 = ((_net_1838)?data_in332:10'b0)|
    (((_reg_2|_net_568))?_add_all_x_data_out_org332:10'b0);
   assign  data_out_org333 = ((_net_1837)?data_in333:10'b0)|
    (((_reg_2|_net_567))?_add_all_x_data_out_org333:10'b0);
   assign  data_out_org334 = ((_net_1836)?data_in334:10'b0)|
    (((_reg_2|_net_566))?_add_all_x_data_out_org334:10'b0);
   assign  data_out_org335 = ((_net_1835)?data_in335:10'b0)|
    (((_reg_2|_net_565))?_add_all_x_data_out_org335:10'b0);
   assign  data_out_org336 = ((_net_1834)?data_in336:10'b0)|
    (((_reg_2|_net_564))?_add_all_x_data_out_org336:10'b0);
   assign  data_out_org337 = ((_net_1833)?data_in337:10'b0)|
    (((_reg_2|_net_563))?_add_all_x_data_out_org337:10'b0);
   assign  data_out_org338 = ((_net_1832)?data_in338:10'b0)|
    (((_reg_2|_net_562))?_add_all_x_data_out_org338:10'b0);
   assign  data_out_org339 = ((_net_1831)?data_in339:10'b0)|
    (((_reg_2|_net_561))?_add_all_x_data_out_org339:10'b0);
   assign  data_out_org340 = ((_net_1830)?data_in340:10'b0)|
    (((_reg_2|_net_560))?_add_all_x_data_out_org340:10'b0);
   assign  data_out_org341 = ((_net_1829)?data_in341:10'b0)|
    (((_reg_2|_net_559))?_add_all_x_data_out_org341:10'b0);
   assign  data_out_org342 = ((_net_1828)?data_in342:10'b0)|
    (((_reg_2|_net_558))?_add_all_x_data_out_org342:10'b0);
   assign  data_out_org343 = ((_net_1827)?data_in343:10'b0)|
    (((_reg_2|_net_557))?_add_all_x_data_out_org343:10'b0);
   assign  data_out_org344 = ((_net_1826)?data_in344:10'b0)|
    (((_reg_2|_net_556))?_add_all_x_data_out_org344:10'b0);
   assign  data_out_org345 = ((_net_1825)?data_in345:10'b0)|
    (((_reg_2|_net_555))?_add_all_x_data_out_org345:10'b0);
   assign  data_out_org346 = ((_net_1824)?data_in346:10'b0)|
    (((_reg_2|_net_554))?_add_all_x_data_out_org346:10'b0);
   assign  data_out_org347 = ((_net_1823)?data_in347:10'b0)|
    (((_reg_2|_net_553))?_add_all_x_data_out_org347:10'b0);
   assign  data_out_org348 = ((_net_1822)?data_in348:10'b0)|
    (((_reg_2|_net_552))?_add_all_x_data_out_org348:10'b0);
   assign  data_out_org349 = ((_net_1821)?data_in349:10'b0)|
    (((_reg_2|_net_551))?_add_all_x_data_out_org349:10'b0);
   assign  data_out_org350 = ((_net_1820)?data_in350:10'b0)|
    (((_reg_2|_net_550))?_add_all_x_data_out_org350:10'b0);
   assign  data_out_org353 = ((_net_1819)?data_in353:10'b0)|
    (((_reg_2|_net_549))?_add_all_x_data_out_org353:10'b0);
   assign  data_out_org354 = ((_net_1818)?data_in354:10'b0)|
    (((_reg_2|_net_548))?_add_all_x_data_out_org354:10'b0);
   assign  data_out_org355 = ((_net_1817)?data_in355:10'b0)|
    (((_reg_2|_net_547))?_add_all_x_data_out_org355:10'b0);
   assign  data_out_org356 = ((_net_1816)?data_in356:10'b0)|
    (((_reg_2|_net_546))?_add_all_x_data_out_org356:10'b0);
   assign  data_out_org357 = ((_net_1815)?data_in357:10'b0)|
    (((_reg_2|_net_545))?_add_all_x_data_out_org357:10'b0);
   assign  data_out_org358 = ((_net_1814)?data_in358:10'b0)|
    (((_reg_2|_net_544))?_add_all_x_data_out_org358:10'b0);
   assign  data_out_org359 = ((_net_1813)?data_in359:10'b0)|
    (((_reg_2|_net_543))?_add_all_x_data_out_org359:10'b0);
   assign  data_out_org360 = ((_net_1812)?data_in360:10'b0)|
    (((_reg_2|_net_542))?_add_all_x_data_out_org360:10'b0);
   assign  data_out_org361 = ((_net_1811)?data_in361:10'b0)|
    (((_reg_2|_net_541))?_add_all_x_data_out_org361:10'b0);
   assign  data_out_org362 = ((_net_1810)?data_in362:10'b0)|
    (((_reg_2|_net_540))?_add_all_x_data_out_org362:10'b0);
   assign  data_out_org363 = ((_net_1809)?data_in363:10'b0)|
    (((_reg_2|_net_539))?_add_all_x_data_out_org363:10'b0);
   assign  data_out_org364 = ((_net_1808)?data_in364:10'b0)|
    (((_reg_2|_net_538))?_add_all_x_data_out_org364:10'b0);
   assign  data_out_org365 = ((_net_1807)?data_in365:10'b0)|
    (((_reg_2|_net_537))?_add_all_x_data_out_org365:10'b0);
   assign  data_out_org366 = ((_net_1806)?data_in366:10'b0)|
    (((_reg_2|_net_536))?_add_all_x_data_out_org366:10'b0);
   assign  data_out_org367 = ((_net_1805)?data_in367:10'b0)|
    (((_reg_2|_net_535))?_add_all_x_data_out_org367:10'b0);
   assign  data_out_org368 = ((_net_1804)?data_in368:10'b0)|
    (((_reg_2|_net_534))?_add_all_x_data_out_org368:10'b0);
   assign  data_out_org369 = ((_net_1803)?data_in369:10'b0)|
    (((_reg_2|_net_533))?_add_all_x_data_out_org369:10'b0);
   assign  data_out_org370 = ((_net_1802)?data_in370:10'b0)|
    (((_reg_2|_net_532))?_add_all_x_data_out_org370:10'b0);
   assign  data_out_org371 = ((_net_1801)?data_in371:10'b0)|
    (((_reg_2|_net_531))?_add_all_x_data_out_org371:10'b0);
   assign  data_out_org372 = ((_net_1800)?data_in372:10'b0)|
    (((_reg_2|_net_530))?_add_all_x_data_out_org372:10'b0);
   assign  data_out_org373 = ((_net_1799)?data_in373:10'b0)|
    (((_reg_2|_net_529))?_add_all_x_data_out_org373:10'b0);
   assign  data_out_org374 = ((_net_1798)?data_in374:10'b0)|
    (((_reg_2|_net_528))?_add_all_x_data_out_org374:10'b0);
   assign  data_out_org375 = ((_net_1797)?data_in375:10'b0)|
    (((_reg_2|_net_527))?_add_all_x_data_out_org375:10'b0);
   assign  data_out_org376 = ((_net_1796)?data_in376:10'b0)|
    (((_reg_2|_net_526))?_add_all_x_data_out_org376:10'b0);
   assign  data_out_org377 = ((_net_1795)?data_in377:10'b0)|
    (((_reg_2|_net_525))?_add_all_x_data_out_org377:10'b0);
   assign  data_out_org378 = ((_net_1794)?data_in378:10'b0)|
    (((_reg_2|_net_524))?_add_all_x_data_out_org378:10'b0);
   assign  data_out_org379 = ((_net_1793)?data_in379:10'b0)|
    (((_reg_2|_net_523))?_add_all_x_data_out_org379:10'b0);
   assign  data_out_org380 = ((_net_1792)?data_in380:10'b0)|
    (((_reg_2|_net_522))?_add_all_x_data_out_org380:10'b0);
   assign  data_out_org381 = ((_net_1791)?data_in381:10'b0)|
    (((_reg_2|_net_521))?_add_all_x_data_out_org381:10'b0);
   assign  data_out_org382 = ((_net_1790)?data_in382:10'b0)|
    (((_reg_2|_net_520))?_add_all_x_data_out_org382:10'b0);
   assign  data_out_org385 = ((_net_1789)?data_in385:10'b0)|
    (((_reg_2|_net_519))?_add_all_x_data_out_org385:10'b0);
   assign  data_out_org386 = ((_net_1788)?data_in386:10'b0)|
    (((_reg_2|_net_518))?_add_all_x_data_out_org386:10'b0);
   assign  data_out_org387 = ((_net_1787)?data_in387:10'b0)|
    (((_reg_2|_net_517))?_add_all_x_data_out_org387:10'b0);
   assign  data_out_org388 = ((_net_1786)?data_in388:10'b0)|
    (((_reg_2|_net_516))?_add_all_x_data_out_org388:10'b0);
   assign  data_out_org389 = ((_net_1785)?data_in389:10'b0)|
    (((_reg_2|_net_515))?_add_all_x_data_out_org389:10'b0);
   assign  data_out_org390 = ((_net_1784)?data_in390:10'b0)|
    (((_reg_2|_net_514))?_add_all_x_data_out_org390:10'b0);
   assign  data_out_org391 = ((_net_1783)?data_in391:10'b0)|
    (((_reg_2|_net_513))?_add_all_x_data_out_org391:10'b0);
   assign  data_out_org392 = ((_net_1782)?data_in392:10'b0)|
    (((_reg_2|_net_512))?_add_all_x_data_out_org392:10'b0);
   assign  data_out_org393 = ((_net_1781)?data_in393:10'b0)|
    (((_reg_2|_net_511))?_add_all_x_data_out_org393:10'b0);
   assign  data_out_org394 = ((_net_1780)?data_in394:10'b0)|
    (((_reg_2|_net_510))?_add_all_x_data_out_org394:10'b0);
   assign  data_out_org395 = ((_net_1779)?data_in395:10'b0)|
    (((_reg_2|_net_509))?_add_all_x_data_out_org395:10'b0);
   assign  data_out_org396 = ((_net_1778)?data_in396:10'b0)|
    (((_reg_2|_net_508))?_add_all_x_data_out_org396:10'b0);
   assign  data_out_org397 = ((_net_1777)?data_in397:10'b0)|
    (((_reg_2|_net_507))?_add_all_x_data_out_org397:10'b0);
   assign  data_out_org398 = ((_net_1776)?data_in398:10'b0)|
    (((_reg_2|_net_506))?_add_all_x_data_out_org398:10'b0);
   assign  data_out_org399 = ((_net_1775)?data_in399:10'b0)|
    (((_reg_2|_net_505))?_add_all_x_data_out_org399:10'b0);
   assign  data_out_org400 = ((_net_1774)?data_in400:10'b0)|
    (((_reg_2|_net_504))?_add_all_x_data_out_org400:10'b0);
   assign  data_out_org401 = ((_net_1773)?data_in401:10'b0)|
    (((_reg_2|_net_503))?_add_all_x_data_out_org401:10'b0);
   assign  data_out_org402 = ((_net_1772)?data_in402:10'b0)|
    (((_reg_2|_net_502))?_add_all_x_data_out_org402:10'b0);
   assign  data_out_org403 = ((_net_1771)?data_in403:10'b0)|
    (((_reg_2|_net_501))?_add_all_x_data_out_org403:10'b0);
   assign  data_out_org404 = ((_net_1770)?data_in404:10'b0)|
    (((_reg_2|_net_500))?_add_all_x_data_out_org404:10'b0);
   assign  data_out_org405 = ((_net_1769)?data_in405:10'b0)|
    (((_reg_2|_net_499))?_add_all_x_data_out_org405:10'b0);
   assign  data_out_org406 = ((_net_1768)?data_in406:10'b0)|
    (((_reg_2|_net_498))?_add_all_x_data_out_org406:10'b0);
   assign  data_out_org407 = ((_net_1767)?data_in407:10'b0)|
    (((_reg_2|_net_497))?_add_all_x_data_out_org407:10'b0);
   assign  data_out_org408 = ((_net_1766)?data_in408:10'b0)|
    (((_reg_2|_net_496))?_add_all_x_data_out_org408:10'b0);
   assign  data_out_org409 = ((_net_1765)?data_in409:10'b0)|
    (((_reg_2|_net_495))?_add_all_x_data_out_org409:10'b0);
   assign  data_out_org410 = ((_net_1764)?data_in410:10'b0)|
    (((_reg_2|_net_494))?_add_all_x_data_out_org410:10'b0);
   assign  data_out_org411 = ((_net_1763)?data_in411:10'b0)|
    (((_reg_2|_net_493))?_add_all_x_data_out_org411:10'b0);
   assign  data_out_org412 = ((_net_1762)?data_in412:10'b0)|
    (((_reg_2|_net_492))?_add_all_x_data_out_org412:10'b0);
   assign  data_out_org413 = ((_net_1761)?data_in413:10'b0)|
    (((_reg_2|_net_491))?_add_all_x_data_out_org413:10'b0);
   assign  data_out_org414 = ((_net_1760)?data_in414:10'b0)|
    (((_reg_2|_net_490))?_add_all_x_data_out_org414:10'b0);
   assign  data_out_org417 = ((_net_1759)?data_in417:10'b0)|
    (((_reg_2|_net_489))?_add_all_x_data_out_org417:10'b0);
   assign  data_out_org418 = ((_net_1758)?data_in418:10'b0)|
    (((_reg_2|_net_488))?_add_all_x_data_out_org418:10'b0);
   assign  data_out_org419 = ((_net_1757)?data_in419:10'b0)|
    (((_reg_2|_net_487))?_add_all_x_data_out_org419:10'b0);
   assign  data_out_org420 = ((_net_1756)?data_in420:10'b0)|
    (((_reg_2|_net_486))?_add_all_x_data_out_org420:10'b0);
   assign  data_out_org421 = ((_net_1755)?data_in421:10'b0)|
    (((_reg_2|_net_485))?_add_all_x_data_out_org421:10'b0);
   assign  data_out_org422 = ((_net_1754)?data_in422:10'b0)|
    (((_reg_2|_net_484))?_add_all_x_data_out_org422:10'b0);
   assign  data_out_org423 = ((_net_1753)?data_in423:10'b0)|
    (((_reg_2|_net_483))?_add_all_x_data_out_org423:10'b0);
   assign  data_out_org424 = ((_net_1752)?data_in424:10'b0)|
    (((_reg_2|_net_482))?_add_all_x_data_out_org424:10'b0);
   assign  data_out_org425 = ((_net_1751)?data_in425:10'b0)|
    (((_reg_2|_net_481))?_add_all_x_data_out_org425:10'b0);
   assign  data_out_org426 = ((_net_1750)?data_in426:10'b0)|
    (((_reg_2|_net_480))?_add_all_x_data_out_org426:10'b0);
   assign  data_out_org427 = ((_net_1749)?data_in427:10'b0)|
    (((_reg_2|_net_479))?_add_all_x_data_out_org427:10'b0);
   assign  data_out_org428 = ((_net_1748)?data_in428:10'b0)|
    (((_reg_2|_net_478))?_add_all_x_data_out_org428:10'b0);
   assign  data_out_org429 = ((_net_1747)?data_in429:10'b0)|
    (((_reg_2|_net_477))?_add_all_x_data_out_org429:10'b0);
   assign  data_out_org430 = ((_net_1746)?data_in430:10'b0)|
    (((_reg_2|_net_476))?_add_all_x_data_out_org430:10'b0);
   assign  data_out_org431 = ((_net_1745)?data_in431:10'b0)|
    (((_reg_2|_net_475))?_add_all_x_data_out_org431:10'b0);
   assign  data_out_org432 = ((_net_1744)?data_in432:10'b0)|
    (((_reg_2|_net_474))?_add_all_x_data_out_org432:10'b0);
   assign  data_out_org433 = ((_net_1743)?data_in433:10'b0)|
    (((_reg_2|_net_473))?_add_all_x_data_out_org433:10'b0);
   assign  data_out_org434 = ((_net_1742)?data_in434:10'b0)|
    (((_reg_2|_net_472))?_add_all_x_data_out_org434:10'b0);
   assign  data_out_org435 = ((_net_1741)?data_in435:10'b0)|
    (((_reg_2|_net_471))?_add_all_x_data_out_org435:10'b0);
   assign  data_out_org436 = ((_net_1740)?data_in436:10'b0)|
    (((_reg_2|_net_470))?_add_all_x_data_out_org436:10'b0);
   assign  data_out_org437 = ((_net_1739)?data_in437:10'b0)|
    (((_reg_2|_net_469))?_add_all_x_data_out_org437:10'b0);
   assign  data_out_org438 = ((_net_1738)?data_in438:10'b0)|
    (((_reg_2|_net_468))?_add_all_x_data_out_org438:10'b0);
   assign  data_out_org439 = ((_net_1737)?data_in439:10'b0)|
    (((_reg_2|_net_467))?_add_all_x_data_out_org439:10'b0);
   assign  data_out_org440 = ((_net_1736)?data_in440:10'b0)|
    (((_reg_2|_net_466))?_add_all_x_data_out_org440:10'b0);
   assign  data_out_org441 = ((_net_1735)?data_in441:10'b0)|
    (((_reg_2|_net_465))?_add_all_x_data_out_org441:10'b0);
   assign  data_out_org442 = ((_net_1734)?data_in442:10'b0)|
    (((_reg_2|_net_464))?_add_all_x_data_out_org442:10'b0);
   assign  data_out_org443 = ((_net_1733)?data_in443:10'b0)|
    (((_reg_2|_net_463))?_add_all_x_data_out_org443:10'b0);
   assign  data_out_org444 = ((_net_1732)?data_in444:10'b0)|
    (((_reg_2|_net_462))?_add_all_x_data_out_org444:10'b0);
   assign  data_out_org445 = ((_net_1731)?data_in445:10'b0)|
    (((_reg_2|_net_461))?_add_all_x_data_out_org445:10'b0);
   assign  data_out_org446 = ((_net_1730)?data_in446:10'b0)|
    (((_reg_2|_net_460))?_add_all_x_data_out_org446:10'b0);
   assign  data_out_org449 = ((_net_1729)?data_in449:10'b0)|
    (((_reg_2|_net_459))?_add_all_x_data_out_org449:10'b0);
   assign  data_out_org450 = ((_net_1728)?data_in450:10'b0)|
    (((_reg_2|_net_458))?_add_all_x_data_out_org450:10'b0);
   assign  data_out_org451 = ((_net_1727)?data_in451:10'b0)|
    (((_reg_2|_net_457))?_add_all_x_data_out_org451:10'b0);
   assign  data_out_org452 = ((_net_1726)?data_in452:10'b0)|
    (((_reg_2|_net_456))?_add_all_x_data_out_org452:10'b0);
   assign  data_out_org453 = ((_net_1725)?data_in453:10'b0)|
    (((_reg_2|_net_455))?_add_all_x_data_out_org453:10'b0);
   assign  data_out_org454 = ((_net_1724)?data_in454:10'b0)|
    (((_reg_2|_net_454))?_add_all_x_data_out_org454:10'b0);
   assign  data_out_org455 = ((_net_1723)?data_in455:10'b0)|
    (((_reg_2|_net_453))?_add_all_x_data_out_org455:10'b0);
   assign  data_out_org456 = ((_net_1722)?data_in456:10'b0)|
    (((_reg_2|_net_452))?_add_all_x_data_out_org456:10'b0);
   assign  data_out_org457 = ((_net_1721)?data_in457:10'b0)|
    (((_reg_2|_net_451))?_add_all_x_data_out_org457:10'b0);
   assign  data_out_org458 = ((_net_1720)?data_in458:10'b0)|
    (((_reg_2|_net_450))?_add_all_x_data_out_org458:10'b0);
   assign  data_out_org459 = ((_net_1719)?data_in459:10'b0)|
    (((_reg_2|_net_449))?_add_all_x_data_out_org459:10'b0);
   assign  data_out_org460 = ((_net_1718)?data_in460:10'b0)|
    (((_reg_2|_net_448))?_add_all_x_data_out_org460:10'b0);
   assign  data_out_org461 = ((_net_1717)?data_in461:10'b0)|
    (((_reg_2|_net_447))?_add_all_x_data_out_org461:10'b0);
   assign  data_out_org462 = ((_net_1716)?data_in462:10'b0)|
    (((_reg_2|_net_446))?_add_all_x_data_out_org462:10'b0);
   assign  data_out_org463 = ((_net_1715)?data_in463:10'b0)|
    (((_reg_2|_net_445))?_add_all_x_data_out_org463:10'b0);
   assign  data_out_org464 = ((_net_1714)?data_in464:10'b0)|
    (((_reg_2|_net_444))?_add_all_x_data_out_org464:10'b0);
   assign  data_out_org465 = ((_net_1713)?data_in465:10'b0)|
    (((_reg_2|_net_443))?_add_all_x_data_out_org465:10'b0);
   assign  data_out_org466 = ((_net_1712)?data_in466:10'b0)|
    (((_reg_2|_net_442))?_add_all_x_data_out_org466:10'b0);
   assign  data_out_org467 = ((_net_1711)?data_in467:10'b0)|
    (((_reg_2|_net_441))?_add_all_x_data_out_org467:10'b0);
   assign  data_out_org468 = ((_net_1710)?data_in468:10'b0)|
    (((_reg_2|_net_440))?_add_all_x_data_out_org468:10'b0);
   assign  data_out_org469 = ((_net_1709)?data_in469:10'b0)|
    (((_reg_2|_net_439))?_add_all_x_data_out_org469:10'b0);
   assign  data_out_org470 = ((_net_1708)?data_in470:10'b0)|
    (((_reg_2|_net_438))?_add_all_x_data_out_org470:10'b0);
   assign  data_out_org471 = ((_net_1707)?data_in471:10'b0)|
    (((_reg_2|_net_437))?_add_all_x_data_out_org471:10'b0);
   assign  data_out_org472 = ((_net_1706)?data_in472:10'b0)|
    (((_reg_2|_net_436))?_add_all_x_data_out_org472:10'b0);
   assign  data_out_org473 = ((_net_1705)?data_in473:10'b0)|
    (((_reg_2|_net_435))?_add_all_x_data_out_org473:10'b0);
   assign  data_out_org474 = ((_net_1704)?data_in474:10'b0)|
    (((_reg_2|_net_434))?_add_all_x_data_out_org474:10'b0);
   assign  data_out_org475 = ((_net_1703)?data_in475:10'b0)|
    (((_reg_2|_net_433))?_add_all_x_data_out_org475:10'b0);
   assign  data_out_org476 = ((_net_1702)?data_in476:10'b0)|
    (((_reg_2|_net_432))?_add_all_x_data_out_org476:10'b0);
   assign  data_out_org477 = ((_net_1701)?data_in477:10'b0)|
    (((_reg_2|_net_431))?_add_all_x_data_out_org477:10'b0);
   assign  data_out_org478 = ((_net_1700)?data_in478:10'b0)|
    (((_reg_2|_net_430))?_add_all_x_data_out_org478:10'b0);
   assign  sg33 = ((_net_1699)?2'b00:2'b0)|
    (((_reg_2|_net_429))?_add_all_x_sg_out33:2'b0);
   assign  sg34 = ((_net_1698)?2'b00:2'b0)|
    (((_reg_2|_net_428))?_add_all_x_sg_out34:2'b0);
   assign  sg35 = ((_net_1697)?2'b00:2'b0)|
    (((_reg_2|_net_427))?_add_all_x_sg_out35:2'b0);
   assign  sg36 = ((_net_1696)?2'b00:2'b0)|
    (((_reg_2|_net_426))?_add_all_x_sg_out36:2'b0);
   assign  sg37 = ((_net_1695)?2'b00:2'b0)|
    (((_reg_2|_net_425))?_add_all_x_sg_out37:2'b0);
   assign  sg38 = ((_net_1694)?2'b00:2'b0)|
    (((_reg_2|_net_424))?_add_all_x_sg_out38:2'b0);
   assign  sg39 = ((_net_1693)?2'b00:2'b0)|
    (((_reg_2|_net_423))?_add_all_x_sg_out39:2'b0);
   assign  sg40 = ((_net_1692)?2'b00:2'b0)|
    (((_reg_2|_net_422))?_add_all_x_sg_out40:2'b0);
   assign  sg41 = ((_net_1691)?2'b00:2'b0)|
    (((_reg_2|_net_421))?_add_all_x_sg_out41:2'b0);
   assign  sg42 = ((_net_1690)?2'b00:2'b0)|
    (((_reg_2|_net_420))?_add_all_x_sg_out42:2'b0);
   assign  sg43 = ((_net_1689)?2'b00:2'b0)|
    (((_reg_2|_net_419))?_add_all_x_sg_out43:2'b0);
   assign  sg44 = ((_net_1688)?2'b00:2'b0)|
    (((_reg_2|_net_418))?_add_all_x_sg_out44:2'b0);
   assign  sg45 = ((_net_1687)?2'b00:2'b0)|
    (((_reg_2|_net_417))?_add_all_x_sg_out45:2'b0);
   assign  sg46 = ((_net_1686)?2'b00:2'b0)|
    (((_reg_2|_net_416))?_add_all_x_sg_out46:2'b0);
   assign  sg47 = ((_net_1685)?2'b00:2'b0)|
    (((_reg_2|_net_415))?_add_all_x_sg_out47:2'b0);
   assign  sg48 = ((_net_1684)?2'b00:2'b0)|
    (((_reg_2|_net_414))?_add_all_x_sg_out48:2'b0);
   assign  sg49 = ((_net_1683)?2'b00:2'b0)|
    (((_reg_2|_net_413))?_add_all_x_sg_out49:2'b0);
   assign  sg50 = ((_net_1682)?2'b00:2'b0)|
    (((_reg_2|_net_412))?_add_all_x_sg_out50:2'b0);
   assign  sg51 = ((_net_1681)?2'b00:2'b0)|
    (((_reg_2|_net_411))?_add_all_x_sg_out51:2'b0);
   assign  sg52 = ((_net_1680)?2'b00:2'b0)|
    (((_reg_2|_net_410))?_add_all_x_sg_out52:2'b0);
   assign  sg53 = ((_net_1679)?2'b00:2'b0)|
    (((_reg_2|_net_409))?_add_all_x_sg_out53:2'b0);
   assign  sg54 = ((_net_1678)?2'b00:2'b0)|
    (((_reg_2|_net_408))?_add_all_x_sg_out54:2'b0);
   assign  sg55 = ((_net_1677)?2'b00:2'b0)|
    (((_reg_2|_net_407))?_add_all_x_sg_out55:2'b0);
   assign  sg56 = ((_net_1676)?2'b00:2'b0)|
    (((_reg_2|_net_406))?_add_all_x_sg_out56:2'b0);
   assign  sg57 = ((_net_1675)?2'b00:2'b0)|
    (((_reg_2|_net_405))?_add_all_x_sg_out57:2'b0);
   assign  sg58 = ((_net_1674)?2'b00:2'b0)|
    (((_reg_2|_net_404))?_add_all_x_sg_out58:2'b0);
   assign  sg59 = ((_net_1673)?2'b00:2'b0)|
    (((_reg_2|_net_403))?_add_all_x_sg_out59:2'b0);
   assign  sg60 = ((_net_1672)?2'b00:2'b0)|
    (((_reg_2|_net_402))?_add_all_x_sg_out60:2'b0);
   assign  sg61 = ((_net_1671)?2'b00:2'b0)|
    (((_reg_2|_net_401))?_add_all_x_sg_out61:2'b0);
   assign  sg62 = ((_net_1670)?2'b00:10'b0)|
    (((_reg_2|_net_400))?_add_all_x_sg_out62:10'b0);
   assign  sg65 = ((_net_1669)?2'b00:2'b0)|
    (((_reg_2|_net_399))?_add_all_x_sg_out65:2'b0);
   assign  sg66 = ((_net_1668)?2'b00:2'b0)|
    (((_reg_2|_net_398))?_add_all_x_sg_out66:2'b0);
   assign  sg67 = ((_net_1667)?2'b00:2'b0)|
    (((_reg_2|_net_397))?_add_all_x_sg_out67:2'b0);
   assign  sg68 = ((_net_1666)?2'b00:2'b0)|
    (((_reg_2|_net_396))?_add_all_x_sg_out68:2'b0);
   assign  sg69 = ((_net_1665)?2'b00:2'b0)|
    (((_reg_2|_net_395))?_add_all_x_sg_out69:2'b0);
   assign  sg70 = ((_net_1664)?2'b00:2'b0)|
    (((_reg_2|_net_394))?_add_all_x_sg_out70:2'b0);
   assign  sg71 = ((_net_1663)?2'b00:2'b0)|
    (((_reg_2|_net_393))?_add_all_x_sg_out71:2'b0);
   assign  sg72 = ((_net_1662)?2'b00:2'b0)|
    (((_reg_2|_net_392))?_add_all_x_sg_out72:2'b0);
   assign  sg73 = ((_net_1661)?2'b00:2'b0)|
    (((_reg_2|_net_391))?_add_all_x_sg_out73:2'b0);
   assign  sg74 = ((_net_1660)?2'b00:2'b0)|
    (((_reg_2|_net_390))?_add_all_x_sg_out74:2'b0);
   assign  sg75 = ((_net_1659)?2'b00:2'b0)|
    (((_reg_2|_net_389))?_add_all_x_sg_out75:2'b0);
   assign  sg76 = ((_net_1658)?2'b00:2'b0)|
    (((_reg_2|_net_388))?_add_all_x_sg_out76:2'b0);
   assign  sg77 = ((_net_1657)?2'b00:2'b0)|
    (((_reg_2|_net_387))?_add_all_x_sg_out77:2'b0);
   assign  sg78 = ((_net_1656)?2'b00:2'b0)|
    (((_reg_2|_net_386))?_add_all_x_sg_out78:2'b0);
   assign  sg79 = ((_net_1655)?2'b00:2'b0)|
    (((_reg_2|_net_385))?_add_all_x_sg_out79:2'b0);
   assign  sg80 = ((_net_1654)?2'b00:2'b0)|
    (((_reg_2|_net_384))?_add_all_x_sg_out80:2'b0);
   assign  sg81 = ((_net_1653)?2'b00:2'b0)|
    (((_reg_2|_net_383))?_add_all_x_sg_out81:2'b0);
   assign  sg82 = ((_net_1652)?2'b00:2'b0)|
    (((_reg_2|_net_382))?_add_all_x_sg_out82:2'b0);
   assign  sg83 = ((_net_1651)?2'b00:2'b0)|
    (((_reg_2|_net_381))?_add_all_x_sg_out83:2'b0);
   assign  sg84 = ((_net_1650)?2'b00:2'b0)|
    (((_reg_2|_net_380))?_add_all_x_sg_out84:2'b0);
   assign  sg85 = ((_net_1649)?2'b00:2'b0)|
    (((_reg_2|_net_379))?_add_all_x_sg_out85:2'b0);
   assign  sg86 = ((_net_1648)?2'b00:2'b0)|
    (((_reg_2|_net_378))?_add_all_x_sg_out86:2'b0);
   assign  sg87 = ((_net_1647)?2'b00:2'b0)|
    (((_reg_2|_net_377))?_add_all_x_sg_out87:2'b0);
   assign  sg88 = ((_net_1646)?2'b00:2'b0)|
    (((_reg_2|_net_376))?_add_all_x_sg_out88:2'b0);
   assign  sg89 = ((_net_1645)?2'b00:2'b0)|
    (((_reg_2|_net_375))?_add_all_x_sg_out89:2'b0);
   assign  sg90 = ((_net_1644)?2'b00:2'b0)|
    (((_reg_2|_net_374))?_add_all_x_sg_out90:2'b0);
   assign  sg91 = ((_net_1643)?2'b00:2'b0)|
    (((_reg_2|_net_373))?_add_all_x_sg_out91:2'b0);
   assign  sg92 = ((_net_1642)?2'b00:2'b0)|
    (((_reg_2|_net_372))?_add_all_x_sg_out92:2'b0);
   assign  sg93 = ((_net_1641)?2'b00:2'b0)|
    (((_reg_2|_net_371))?_add_all_x_sg_out93:2'b0);
   assign  sg94 = ((_net_1640)?2'b00:10'b0)|
    (((_reg_2|_net_370))?_add_all_x_sg_out94:10'b0);
   assign  sg97 = ((_net_1639)?2'b00:2'b0)|
    (((_reg_2|_net_369))?_add_all_x_sg_out97:2'b0);
   assign  sg98 = ((_net_1638)?2'b00:2'b0)|
    (((_reg_2|_net_368))?_add_all_x_sg_out98:2'b0);
   assign  sg99 = ((_net_1637)?2'b00:2'b0)|
    (((_reg_2|_net_367))?_add_all_x_sg_out99:2'b0);
   assign  sg100 = ((_net_1636)?2'b00:2'b0)|
    (((_reg_2|_net_366))?_add_all_x_sg_out100:2'b0);
   assign  sg101 = ((_net_1635)?2'b00:2'b0)|
    (((_reg_2|_net_365))?_add_all_x_sg_out101:2'b0);
   assign  sg102 = ((_net_1634)?2'b00:2'b0)|
    (((_reg_2|_net_364))?_add_all_x_sg_out102:2'b0);
   assign  sg103 = ((_net_1633)?2'b00:2'b0)|
    (((_reg_2|_net_363))?_add_all_x_sg_out103:2'b0);
   assign  sg104 = ((_net_1632)?2'b00:2'b0)|
    (((_reg_2|_net_362))?_add_all_x_sg_out104:2'b0);
   assign  sg105 = ((_net_1631)?2'b00:2'b0)|
    (((_reg_2|_net_361))?_add_all_x_sg_out105:2'b0);
   assign  sg106 = ((_net_1630)?2'b00:2'b0)|
    (((_reg_2|_net_360))?_add_all_x_sg_out106:2'b0);
   assign  sg107 = ((_net_1629)?2'b00:2'b0)|
    (((_reg_2|_net_359))?_add_all_x_sg_out107:2'b0);
   assign  sg108 = ((_net_1628)?2'b00:2'b0)|
    (((_reg_2|_net_358))?_add_all_x_sg_out108:2'b0);
   assign  sg109 = ((_net_1627)?2'b00:2'b0)|
    (((_reg_2|_net_357))?_add_all_x_sg_out109:2'b0);
   assign  sg110 = ((_net_1626)?2'b00:2'b0)|
    (((_reg_2|_net_356))?_add_all_x_sg_out110:2'b0);
   assign  sg111 = ((_net_1625)?2'b00:2'b0)|
    (((_reg_2|_net_355))?_add_all_x_sg_out111:2'b0);
   assign  sg112 = ((_net_1624)?2'b00:2'b0)|
    (((_reg_2|_net_354))?_add_all_x_sg_out112:2'b0);
   assign  sg113 = ((_net_1623)?2'b00:2'b0)|
    (((_reg_2|_net_353))?_add_all_x_sg_out113:2'b0);
   assign  sg114 = ((_net_1622)?2'b00:2'b0)|
    (((_reg_2|_net_352))?_add_all_x_sg_out114:2'b0);
   assign  sg115 = ((_net_1621)?2'b00:2'b0)|
    (((_reg_2|_net_351))?_add_all_x_sg_out115:2'b0);
   assign  sg116 = ((_net_1620)?2'b00:2'b0)|
    (((_reg_2|_net_350))?_add_all_x_sg_out116:2'b0);
   assign  sg117 = ((_net_1619)?2'b00:2'b0)|
    (((_reg_2|_net_349))?_add_all_x_sg_out117:2'b0);
   assign  sg118 = ((_net_1618)?2'b00:2'b0)|
    (((_reg_2|_net_348))?_add_all_x_sg_out118:2'b0);
   assign  sg119 = ((_net_1617)?2'b00:2'b0)|
    (((_reg_2|_net_347))?_add_all_x_sg_out119:2'b0);
   assign  sg120 = ((_net_1616)?2'b00:2'b0)|
    (((_reg_2|_net_346))?_add_all_x_sg_out120:2'b0);
   assign  sg121 = ((_net_1615)?2'b00:2'b0)|
    (((_reg_2|_net_345))?_add_all_x_sg_out121:2'b0);
   assign  sg122 = ((_net_1614)?2'b00:2'b0)|
    (((_reg_2|_net_344))?_add_all_x_sg_out122:2'b0);
   assign  sg123 = ((_net_1613)?2'b00:2'b0)|
    (((_reg_2|_net_343))?_add_all_x_sg_out123:2'b0);
   assign  sg124 = ((_net_1612)?2'b00:2'b0)|
    (((_reg_2|_net_342))?_add_all_x_sg_out124:2'b0);
   assign  sg125 = ((_net_1611)?2'b00:2'b0)|
    (((_reg_2|_net_341))?_add_all_x_sg_out125:2'b0);
   assign  sg126 = ((_net_1610)?2'b00:10'b0)|
    (((_reg_2|_net_340))?_add_all_x_sg_out126:10'b0);
   assign  sg129 = ((_net_1609)?2'b00:2'b0)|
    (((_reg_2|_net_339))?_add_all_x_sg_out129:2'b0);
   assign  sg130 = ((_net_1608)?2'b00:2'b0)|
    (((_reg_2|_net_338))?_add_all_x_sg_out130:2'b0);
   assign  sg131 = ((_net_1607)?2'b00:2'b0)|
    (((_reg_2|_net_337))?_add_all_x_sg_out131:2'b0);
   assign  sg132 = ((_net_1606)?2'b00:2'b0)|
    (((_reg_2|_net_336))?_add_all_x_sg_out132:2'b0);
   assign  sg133 = ((_net_1605)?2'b00:2'b0)|
    (((_reg_2|_net_335))?_add_all_x_sg_out133:2'b0);
   assign  sg134 = ((_net_1604)?2'b00:2'b0)|
    (((_reg_2|_net_334))?_add_all_x_sg_out134:2'b0);
   assign  sg135 = ((_net_1603)?2'b00:2'b0)|
    (((_reg_2|_net_333))?_add_all_x_sg_out135:2'b0);
   assign  sg136 = ((_net_1602)?2'b00:2'b0)|
    (((_reg_2|_net_332))?_add_all_x_sg_out136:2'b0);
   assign  sg137 = ((_net_1601)?2'b00:2'b0)|
    (((_reg_2|_net_331))?_add_all_x_sg_out137:2'b0);
   assign  sg138 = ((_net_1600)?2'b00:2'b0)|
    (((_reg_2|_net_330))?_add_all_x_sg_out138:2'b0);
   assign  sg139 = ((_net_1599)?2'b00:2'b0)|
    (((_reg_2|_net_329))?_add_all_x_sg_out139:2'b0);
   assign  sg140 = ((_net_1598)?2'b00:2'b0)|
    (((_reg_2|_net_328))?_add_all_x_sg_out140:2'b0);
   assign  sg141 = ((_net_1597)?2'b00:2'b0)|
    (((_reg_2|_net_327))?_add_all_x_sg_out141:2'b0);
   assign  sg142 = ((_net_1596)?2'b00:2'b0)|
    (((_reg_2|_net_326))?_add_all_x_sg_out142:2'b0);
   assign  sg143 = ((_net_1595)?2'b00:2'b0)|
    (((_reg_2|_net_325))?_add_all_x_sg_out143:2'b0);
   assign  sg144 = ((_net_1594)?2'b00:2'b0)|
    (((_reg_2|_net_324))?_add_all_x_sg_out144:2'b0);
   assign  sg145 = ((_net_1593)?2'b00:2'b0)|
    (((_reg_2|_net_323))?_add_all_x_sg_out145:2'b0);
   assign  sg146 = ((_net_1592)?2'b00:2'b0)|
    (((_reg_2|_net_322))?_add_all_x_sg_out146:2'b0);
   assign  sg147 = ((_net_1591)?2'b00:2'b0)|
    (((_reg_2|_net_321))?_add_all_x_sg_out147:2'b0);
   assign  sg148 = ((_net_1590)?2'b00:2'b0)|
    (((_reg_2|_net_320))?_add_all_x_sg_out148:2'b0);
   assign  sg149 = ((_net_1589)?2'b00:2'b0)|
    (((_reg_2|_net_319))?_add_all_x_sg_out149:2'b0);
   assign  sg150 = ((_net_1588)?2'b00:2'b0)|
    (((_reg_2|_net_318))?_add_all_x_sg_out150:2'b0);
   assign  sg151 = ((_net_1587)?2'b00:2'b0)|
    (((_reg_2|_net_317))?_add_all_x_sg_out151:2'b0);
   assign  sg152 = ((_net_1586)?2'b00:2'b0)|
    (((_reg_2|_net_316))?_add_all_x_sg_out152:2'b0);
   assign  sg153 = ((_net_1585)?2'b00:2'b0)|
    (((_reg_2|_net_315))?_add_all_x_sg_out153:2'b0);
   assign  sg154 = ((_net_1584)?2'b00:2'b0)|
    (((_reg_2|_net_314))?_add_all_x_sg_out154:2'b0);
   assign  sg155 = ((_net_1583)?2'b00:2'b0)|
    (((_reg_2|_net_313))?_add_all_x_sg_out155:2'b0);
   assign  sg156 = ((_net_1582)?2'b00:2'b0)|
    (((_reg_2|_net_312))?_add_all_x_sg_out156:2'b0);
   assign  sg157 = ((_net_1581)?2'b00:2'b0)|
    (((_reg_2|_net_311))?_add_all_x_sg_out157:2'b0);
   assign  sg158 = ((_net_1580)?2'b00:10'b0)|
    (((_reg_2|_net_310))?_add_all_x_sg_out158:10'b0);
   assign  sg161 = ((_net_1579)?2'b00:2'b0)|
    (((_reg_2|_net_309))?_add_all_x_sg_out161:2'b0);
   assign  sg162 = ((_net_1578)?2'b00:2'b0)|
    (((_reg_2|_net_308))?_add_all_x_sg_out162:2'b0);
   assign  sg163 = ((_net_1577)?2'b00:2'b0)|
    (((_reg_2|_net_307))?_add_all_x_sg_out163:2'b0);
   assign  sg164 = ((_net_1576)?2'b00:2'b0)|
    (((_reg_2|_net_306))?_add_all_x_sg_out164:2'b0);
   assign  sg165 = ((_net_1575)?2'b00:2'b0)|
    (((_reg_2|_net_305))?_add_all_x_sg_out165:2'b0);
   assign  sg166 = ((_net_1574)?2'b00:2'b0)|
    (((_reg_2|_net_304))?_add_all_x_sg_out166:2'b0);
   assign  sg167 = ((_net_1573)?2'b00:2'b0)|
    (((_reg_2|_net_303))?_add_all_x_sg_out167:2'b0);
   assign  sg168 = ((_net_1572)?2'b00:2'b0)|
    (((_reg_2|_net_302))?_add_all_x_sg_out168:2'b0);
   assign  sg169 = ((_net_1571)?2'b00:2'b0)|
    (((_reg_2|_net_301))?_add_all_x_sg_out169:2'b0);
   assign  sg170 = ((_net_1570)?2'b00:2'b0)|
    (((_reg_2|_net_300))?_add_all_x_sg_out170:2'b0);
   assign  sg171 = ((_net_1569)?2'b00:2'b0)|
    (((_reg_2|_net_299))?_add_all_x_sg_out171:2'b0);
   assign  sg172 = ((_net_1568)?2'b00:2'b0)|
    (((_reg_2|_net_298))?_add_all_x_sg_out172:2'b0);
   assign  sg173 = ((_net_1567)?2'b00:2'b0)|
    (((_reg_2|_net_297))?_add_all_x_sg_out173:2'b0);
   assign  sg174 = ((_net_1566)?2'b00:2'b0)|
    (((_reg_2|_net_296))?_add_all_x_sg_out174:2'b0);
   assign  sg175 = ((_net_1565)?2'b00:2'b0)|
    (((_reg_2|_net_295))?_add_all_x_sg_out175:2'b0);
   assign  sg176 = ((_net_1564)?2'b00:2'b0)|
    (((_reg_2|_net_294))?_add_all_x_sg_out176:2'b0);
   assign  sg177 = ((_net_1563)?2'b00:2'b0)|
    (((_reg_2|_net_293))?_add_all_x_sg_out177:2'b0);
   assign  sg178 = ((_net_1562)?2'b00:2'b0)|
    (((_reg_2|_net_292))?_add_all_x_sg_out178:2'b0);
   assign  sg179 = ((_net_1561)?2'b00:2'b0)|
    (((_reg_2|_net_291))?_add_all_x_sg_out179:2'b0);
   assign  sg180 = ((_net_1560)?2'b00:2'b0)|
    (((_reg_2|_net_290))?_add_all_x_sg_out180:2'b0);
   assign  sg181 = ((_net_1559)?2'b00:2'b0)|
    (((_reg_2|_net_289))?_add_all_x_sg_out181:2'b0);
   assign  sg182 = ((_net_1558)?2'b00:2'b0)|
    (((_reg_2|_net_288))?_add_all_x_sg_out182:2'b0);
   assign  sg183 = ((_net_1557)?2'b00:2'b0)|
    (((_reg_2|_net_287))?_add_all_x_sg_out183:2'b0);
   assign  sg184 = ((_net_1556)?2'b00:2'b0)|
    (((_reg_2|_net_286))?_add_all_x_sg_out184:2'b0);
   assign  sg185 = ((_net_1555)?2'b00:2'b0)|
    (((_reg_2|_net_285))?_add_all_x_sg_out185:2'b0);
   assign  sg186 = ((_net_1554)?2'b00:2'b0)|
    (((_reg_2|_net_284))?_add_all_x_sg_out186:2'b0);
   assign  sg187 = ((_net_1553)?2'b00:2'b0)|
    (((_reg_2|_net_283))?_add_all_x_sg_out187:2'b0);
   assign  sg188 = ((_net_1552)?2'b00:2'b0)|
    (((_reg_2|_net_282))?_add_all_x_sg_out188:2'b0);
   assign  sg189 = ((_net_1551)?2'b00:2'b0)|
    (((_reg_2|_net_281))?_add_all_x_sg_out189:2'b0);
   assign  sg190 = ((_net_1550)?2'b00:10'b0)|
    (((_reg_2|_net_280))?_add_all_x_sg_out190:10'b0);
   assign  sg193 = ((_net_1549)?2'b00:2'b0)|
    (((_reg_2|_net_279))?_add_all_x_sg_out193:2'b0);
   assign  sg194 = ((_net_1548)?2'b00:2'b0)|
    (((_reg_2|_net_278))?_add_all_x_sg_out194:2'b0);
   assign  sg195 = ((_net_1547)?2'b00:2'b0)|
    (((_reg_2|_net_277))?_add_all_x_sg_out195:2'b0);
   assign  sg196 = ((_net_1546)?2'b00:2'b0)|
    (((_reg_2|_net_276))?_add_all_x_sg_out196:2'b0);
   assign  sg197 = ((_net_1545)?2'b00:2'b0)|
    (((_reg_2|_net_275))?_add_all_x_sg_out197:2'b0);
   assign  sg198 = ((_net_1544)?2'b00:2'b0)|
    (((_reg_2|_net_274))?_add_all_x_sg_out198:2'b0);
   assign  sg199 = ((_net_1543)?2'b00:2'b0)|
    (((_reg_2|_net_273))?_add_all_x_sg_out199:2'b0);
   assign  sg200 = ((_net_1542)?2'b00:2'b0)|
    (((_reg_2|_net_272))?_add_all_x_sg_out200:2'b0);
   assign  sg201 = ((_net_1541)?2'b00:2'b0)|
    (((_reg_2|_net_271))?_add_all_x_sg_out201:2'b0);
   assign  sg202 = ((_net_1540)?2'b00:2'b0)|
    (((_reg_2|_net_270))?_add_all_x_sg_out202:2'b0);
   assign  sg203 = ((_net_1539)?2'b00:2'b0)|
    (((_reg_2|_net_269))?_add_all_x_sg_out203:2'b0);
   assign  sg204 = ((_net_1538)?2'b00:2'b0)|
    (((_reg_2|_net_268))?_add_all_x_sg_out204:2'b0);
   assign  sg205 = ((_net_1537)?2'b00:2'b0)|
    (((_reg_2|_net_267))?_add_all_x_sg_out205:2'b0);
   assign  sg206 = ((_net_1536)?2'b00:2'b0)|
    (((_reg_2|_net_266))?_add_all_x_sg_out206:2'b0);
   assign  sg207 = ((_net_1535)?2'b00:2'b0)|
    (((_reg_2|_net_265))?_add_all_x_sg_out207:2'b0);
   assign  sg208 = ((_net_1534)?2'b00:2'b0)|
    (((_reg_2|_net_264))?_add_all_x_sg_out208:2'b0);
   assign  sg209 = ((_net_1533)?2'b00:2'b0)|
    (((_reg_2|_net_263))?_add_all_x_sg_out209:2'b0);
   assign  sg210 = ((_net_1532)?2'b00:2'b0)|
    (((_reg_2|_net_262))?_add_all_x_sg_out210:2'b0);
   assign  sg211 = ((_net_1531)?2'b00:2'b0)|
    (((_reg_2|_net_261))?_add_all_x_sg_out211:2'b0);
   assign  sg212 = ((_net_1530)?2'b00:2'b0)|
    (((_reg_2|_net_260))?_add_all_x_sg_out212:2'b0);
   assign  sg213 = ((_net_1529)?2'b00:2'b0)|
    (((_reg_2|_net_259))?_add_all_x_sg_out213:2'b0);
   assign  sg214 = ((_net_1528)?2'b00:2'b0)|
    (((_reg_2|_net_258))?_add_all_x_sg_out214:2'b0);
   assign  sg215 = ((_net_1527)?2'b00:2'b0)|
    (((_reg_2|_net_257))?_add_all_x_sg_out215:2'b0);
   assign  sg216 = ((_net_1526)?2'b00:2'b0)|
    (((_reg_2|_net_256))?_add_all_x_sg_out216:2'b0);
   assign  sg217 = ((_net_1525)?2'b00:2'b0)|
    (((_reg_2|_net_255))?_add_all_x_sg_out217:2'b0);
   assign  sg218 = ((_net_1524)?2'b00:2'b0)|
    (((_reg_2|_net_254))?_add_all_x_sg_out218:2'b0);
   assign  sg219 = ((_net_1523)?2'b00:2'b0)|
    (((_reg_2|_net_253))?_add_all_x_sg_out219:2'b0);
   assign  sg220 = ((_net_1522)?2'b00:2'b0)|
    (((_reg_2|_net_252))?_add_all_x_sg_out220:2'b0);
   assign  sg221 = ((_net_1521)?2'b00:2'b0)|
    (((_reg_2|_net_251))?_add_all_x_sg_out221:2'b0);
   assign  sg222 = ((_net_1520)?2'b00:10'b0)|
    (((_reg_2|_net_250))?_add_all_x_sg_out222:10'b0);
   assign  sg225 = ((_net_1519)?2'b00:2'b0)|
    (((_reg_2|_net_249))?_add_all_x_sg_out225:2'b0);
   assign  sg226 = ((_net_1518)?2'b00:2'b0)|
    (((_reg_2|_net_248))?_add_all_x_sg_out226:2'b0);
   assign  sg227 = ((_net_1517)?2'b00:2'b0)|
    (((_reg_2|_net_247))?_add_all_x_sg_out227:2'b0);
   assign  sg228 = ((_net_1516)?2'b00:2'b0)|
    (((_reg_2|_net_246))?_add_all_x_sg_out228:2'b0);
   assign  sg229 = ((_net_1515)?2'b00:2'b0)|
    (((_reg_2|_net_245))?_add_all_x_sg_out229:2'b0);
   assign  sg230 = ((_net_1514)?2'b00:2'b0)|
    (((_reg_2|_net_244))?_add_all_x_sg_out230:2'b0);
   assign  sg231 = ((_net_1513)?2'b00:2'b0)|
    (((_reg_2|_net_243))?_add_all_x_sg_out231:2'b0);
   assign  sg232 = ((_net_1512)?2'b00:2'b0)|
    (((_reg_2|_net_242))?_add_all_x_sg_out232:2'b0);
   assign  sg233 = ((_net_1511)?2'b00:2'b0)|
    (((_reg_2|_net_241))?_add_all_x_sg_out233:2'b0);
   assign  sg234 = ((_net_1510)?2'b00:2'b0)|
    (((_reg_2|_net_240))?_add_all_x_sg_out234:2'b0);
   assign  sg235 = ((_net_1509)?2'b00:2'b0)|
    (((_reg_2|_net_239))?_add_all_x_sg_out235:2'b0);
   assign  sg236 = ((_net_1508)?2'b00:2'b0)|
    (((_reg_2|_net_238))?_add_all_x_sg_out236:2'b0);
   assign  sg237 = ((_net_1507)?2'b00:2'b0)|
    (((_reg_2|_net_237))?_add_all_x_sg_out237:2'b0);
   assign  sg238 = ((_net_1506)?2'b00:2'b0)|
    (((_reg_2|_net_236))?_add_all_x_sg_out238:2'b0);
   assign  sg239 = ((_net_1505)?2'b00:2'b0)|
    (((_reg_2|_net_235))?_add_all_x_sg_out239:2'b0);
   assign  sg240 = ((_net_1504)?2'b00:2'b0)|
    (((_reg_2|_net_234))?_add_all_x_sg_out240:2'b0);
   assign  sg241 = ((_net_1503)?2'b00:2'b0)|
    (((_reg_2|_net_233))?_add_all_x_sg_out241:2'b0);
   assign  sg242 = ((_net_1502)?2'b00:2'b0)|
    (((_reg_2|_net_232))?_add_all_x_sg_out242:2'b0);
   assign  sg243 = ((_net_1501)?2'b00:2'b0)|
    (((_reg_2|_net_231))?_add_all_x_sg_out243:2'b0);
   assign  sg244 = ((_net_1500)?2'b00:2'b0)|
    (((_reg_2|_net_230))?_add_all_x_sg_out244:2'b0);
   assign  sg245 = ((_net_1499)?2'b00:2'b0)|
    (((_reg_2|_net_229))?_add_all_x_sg_out245:2'b0);
   assign  sg246 = ((_net_1498)?2'b00:2'b0)|
    (((_reg_2|_net_228))?_add_all_x_sg_out246:2'b0);
   assign  sg247 = ((_net_1497)?2'b00:2'b0)|
    (((_reg_2|_net_227))?_add_all_x_sg_out247:2'b0);
   assign  sg248 = ((_net_1496)?2'b00:2'b0)|
    (((_reg_2|_net_226))?_add_all_x_sg_out248:2'b0);
   assign  sg249 = ((_net_1495)?2'b00:2'b0)|
    (((_reg_2|_net_225))?_add_all_x_sg_out249:2'b0);
   assign  sg250 = ((_net_1494)?2'b00:2'b0)|
    (((_reg_2|_net_224))?_add_all_x_sg_out250:2'b0);
   assign  sg251 = ((_net_1493)?2'b00:2'b0)|
    (((_reg_2|_net_223))?_add_all_x_sg_out251:2'b0);
   assign  sg252 = ((_net_1492)?2'b00:2'b0)|
    (((_reg_2|_net_222))?_add_all_x_sg_out252:2'b0);
   assign  sg253 = ((_net_1491)?2'b00:2'b0)|
    (((_reg_2|_net_221))?_add_all_x_sg_out253:2'b0);
   assign  sg254 = ((_net_1490)?2'b00:10'b0)|
    (((_reg_2|_net_220))?_add_all_x_sg_out254:10'b0);
   assign  sg257 = ((_net_1489)?2'b00:2'b0)|
    (((_reg_2|_net_219))?_add_all_x_sg_out257:2'b0);
   assign  sg258 = ((_net_1488)?2'b00:2'b0)|
    (((_reg_2|_net_218))?_add_all_x_sg_out258:2'b0);
   assign  sg259 = ((_net_1487)?2'b00:2'b0)|
    (((_reg_2|_net_217))?_add_all_x_sg_out259:2'b0);
   assign  sg260 = ((_net_1486)?2'b00:2'b0)|
    (((_reg_2|_net_216))?_add_all_x_sg_out260:2'b0);
   assign  sg261 = ((_net_1485)?2'b00:2'b0)|
    (((_reg_2|_net_215))?_add_all_x_sg_out261:2'b0);
   assign  sg262 = ((_net_1484)?2'b00:2'b0)|
    (((_reg_2|_net_214))?_add_all_x_sg_out262:2'b0);
   assign  sg263 = ((_net_1483)?2'b00:2'b0)|
    (((_reg_2|_net_213))?_add_all_x_sg_out263:2'b0);
   assign  sg264 = ((_net_1482)?2'b00:2'b0)|
    (((_reg_2|_net_212))?_add_all_x_sg_out264:2'b0);
   assign  sg265 = ((_net_1481)?2'b00:2'b0)|
    (((_reg_2|_net_211))?_add_all_x_sg_out265:2'b0);
   assign  sg266 = ((_net_1480)?2'b00:2'b0)|
    (((_reg_2|_net_210))?_add_all_x_sg_out266:2'b0);
   assign  sg267 = ((_net_1479)?2'b00:2'b0)|
    (((_reg_2|_net_209))?_add_all_x_sg_out267:2'b0);
   assign  sg268 = ((_net_1478)?2'b00:2'b0)|
    (((_reg_2|_net_208))?_add_all_x_sg_out268:2'b0);
   assign  sg269 = ((_net_1477)?2'b00:2'b0)|
    (((_reg_2|_net_207))?_add_all_x_sg_out269:2'b0);
   assign  sg270 = ((_net_1476)?2'b00:2'b0)|
    (((_reg_2|_net_206))?_add_all_x_sg_out270:2'b0);
   assign  sg271 = ((_net_1475)?2'b00:2'b0)|
    (((_reg_2|_net_205))?_add_all_x_sg_out271:2'b0);
   assign  sg272 = ((_net_1474)?2'b00:2'b0)|
    (((_reg_2|_net_204))?_add_all_x_sg_out272:2'b0);
   assign  sg273 = ((_net_1473)?2'b00:2'b0)|
    (((_reg_2|_net_203))?_add_all_x_sg_out273:2'b0);
   assign  sg274 = ((_net_1472)?2'b00:2'b0)|
    (((_reg_2|_net_202))?_add_all_x_sg_out274:2'b0);
   assign  sg275 = ((_net_1471)?2'b00:2'b0)|
    (((_reg_2|_net_201))?_add_all_x_sg_out275:2'b0);
   assign  sg276 = ((_net_1470)?2'b00:2'b0)|
    (((_reg_2|_net_200))?_add_all_x_sg_out276:2'b0);
   assign  sg277 = ((_net_1469)?2'b00:2'b0)|
    (((_reg_2|_net_199))?_add_all_x_sg_out277:2'b0);
   assign  sg278 = ((_net_1468)?2'b00:2'b0)|
    (((_reg_2|_net_198))?_add_all_x_sg_out278:2'b0);
   assign  sg279 = ((_net_1467)?2'b00:2'b0)|
    (((_reg_2|_net_197))?_add_all_x_sg_out279:2'b0);
   assign  sg280 = ((_net_1466)?2'b00:2'b0)|
    (((_reg_2|_net_196))?_add_all_x_sg_out280:2'b0);
   assign  sg281 = ((_net_1465)?2'b00:2'b0)|
    (((_reg_2|_net_195))?_add_all_x_sg_out281:2'b0);
   assign  sg282 = ((_net_1464)?2'b00:2'b0)|
    (((_reg_2|_net_194))?_add_all_x_sg_out282:2'b0);
   assign  sg283 = ((_net_1463)?2'b00:2'b0)|
    (((_reg_2|_net_193))?_add_all_x_sg_out283:2'b0);
   assign  sg284 = ((_net_1462)?2'b00:2'b0)|
    (((_reg_2|_net_192))?_add_all_x_sg_out284:2'b0);
   assign  sg285 = ((_net_1461)?2'b00:2'b0)|
    (((_reg_2|_net_191))?_add_all_x_sg_out285:2'b0);
   assign  sg286 = ((_net_1460)?2'b00:10'b0)|
    (((_reg_2|_net_190))?_add_all_x_sg_out286:10'b0);
   assign  sg289 = ((_net_1459)?2'b00:2'b0)|
    (((_reg_2|_net_189))?_add_all_x_sg_out289:2'b0);
   assign  sg290 = ((_net_1458)?2'b00:2'b0)|
    (((_reg_2|_net_188))?_add_all_x_sg_out290:2'b0);
   assign  sg291 = ((_net_1457)?2'b00:2'b0)|
    (((_reg_2|_net_187))?_add_all_x_sg_out291:2'b0);
   assign  sg292 = ((_net_1456)?2'b00:2'b0)|
    (((_reg_2|_net_186))?_add_all_x_sg_out292:2'b0);
   assign  sg293 = ((_net_1455)?2'b00:2'b0)|
    (((_reg_2|_net_185))?_add_all_x_sg_out293:2'b0);
   assign  sg294 = ((_net_1454)?2'b00:2'b0)|
    (((_reg_2|_net_184))?_add_all_x_sg_out294:2'b0);
   assign  sg295 = ((_net_1453)?2'b00:2'b0)|
    (((_reg_2|_net_183))?_add_all_x_sg_out295:2'b0);
   assign  sg296 = ((_net_1452)?2'b00:2'b0)|
    (((_reg_2|_net_182))?_add_all_x_sg_out296:2'b0);
   assign  sg297 = ((_net_1451)?2'b00:2'b0)|
    (((_reg_2|_net_181))?_add_all_x_sg_out297:2'b0);
   assign  sg298 = ((_net_1450)?2'b00:2'b0)|
    (((_reg_2|_net_180))?_add_all_x_sg_out298:2'b0);
   assign  sg299 = ((_net_1449)?2'b00:2'b0)|
    (((_reg_2|_net_179))?_add_all_x_sg_out299:2'b0);
   assign  sg300 = ((_net_1448)?2'b00:2'b0)|
    (((_reg_2|_net_178))?_add_all_x_sg_out300:2'b0);
   assign  sg301 = ((_net_1447)?2'b00:2'b0)|
    (((_reg_2|_net_177))?_add_all_x_sg_out301:2'b0);
   assign  sg302 = ((_net_1446)?2'b00:2'b0)|
    (((_reg_2|_net_176))?_add_all_x_sg_out302:2'b0);
   assign  sg303 = ((_net_1445)?2'b00:2'b0)|
    (((_reg_2|_net_175))?_add_all_x_sg_out303:2'b0);
   assign  sg304 = ((_net_1444)?2'b00:2'b0)|
    (((_reg_2|_net_174))?_add_all_x_sg_out304:2'b0);
   assign  sg305 = ((_net_1443)?2'b00:2'b0)|
    (((_reg_2|_net_173))?_add_all_x_sg_out305:2'b0);
   assign  sg306 = ((_net_1442)?2'b00:2'b0)|
    (((_reg_2|_net_172))?_add_all_x_sg_out306:2'b0);
   assign  sg307 = ((_net_1441)?2'b00:2'b0)|
    (((_reg_2|_net_171))?_add_all_x_sg_out307:2'b0);
   assign  sg308 = ((_net_1440)?2'b00:2'b0)|
    (((_reg_2|_net_170))?_add_all_x_sg_out308:2'b0);
   assign  sg309 = ((_net_1439)?2'b00:2'b0)|
    (((_reg_2|_net_169))?_add_all_x_sg_out309:2'b0);
   assign  sg310 = ((_net_1438)?2'b00:2'b0)|
    (((_reg_2|_net_168))?_add_all_x_sg_out310:2'b0);
   assign  sg311 = ((_net_1437)?2'b00:2'b0)|
    (((_reg_2|_net_167))?_add_all_x_sg_out311:2'b0);
   assign  sg312 = ((_net_1436)?2'b00:2'b0)|
    (((_reg_2|_net_166))?_add_all_x_sg_out312:2'b0);
   assign  sg313 = ((_net_1435)?2'b00:2'b0)|
    (((_reg_2|_net_165))?_add_all_x_sg_out313:2'b0);
   assign  sg314 = ((_net_1434)?2'b00:2'b0)|
    (((_reg_2|_net_164))?_add_all_x_sg_out314:2'b0);
   assign  sg315 = ((_net_1433)?2'b00:2'b0)|
    (((_reg_2|_net_163))?_add_all_x_sg_out315:2'b0);
   assign  sg316 = ((_net_1432)?2'b00:2'b0)|
    (((_reg_2|_net_162))?_add_all_x_sg_out316:2'b0);
   assign  sg317 = ((_net_1431)?2'b00:2'b0)|
    (((_reg_2|_net_161))?_add_all_x_sg_out317:2'b0);
   assign  sg318 = ((_net_1430)?2'b00:10'b0)|
    (((_reg_2|_net_160))?_add_all_x_sg_out318:10'b0);
   assign  sg321 = ((_net_1429)?2'b00:2'b0)|
    (((_reg_2|_net_159))?_add_all_x_sg_out321:2'b0);
   assign  sg322 = ((_net_1428)?2'b00:2'b0)|
    (((_reg_2|_net_158))?_add_all_x_sg_out322:2'b0);
   assign  sg323 = ((_net_1427)?2'b00:2'b0)|
    (((_reg_2|_net_157))?_add_all_x_sg_out323:2'b0);
   assign  sg324 = ((_net_1426)?2'b00:2'b0)|
    (((_reg_2|_net_156))?_add_all_x_sg_out324:2'b0);
   assign  sg325 = ((_net_1425)?2'b00:2'b0)|
    (((_reg_2|_net_155))?_add_all_x_sg_out325:2'b0);
   assign  sg326 = ((_net_1424)?2'b00:2'b0)|
    (((_reg_2|_net_154))?_add_all_x_sg_out326:2'b0);
   assign  sg327 = ((_net_1423)?2'b00:2'b0)|
    (((_reg_2|_net_153))?_add_all_x_sg_out327:2'b0);
   assign  sg328 = ((_net_1422)?2'b00:2'b0)|
    (((_reg_2|_net_152))?_add_all_x_sg_out328:2'b0);
   assign  sg329 = ((_net_1421)?2'b00:2'b0)|
    (((_reg_2|_net_151))?_add_all_x_sg_out329:2'b0);
   assign  sg330 = ((_net_1420)?2'b00:2'b0)|
    (((_reg_2|_net_150))?_add_all_x_sg_out330:2'b0);
   assign  sg331 = ((_net_1419)?2'b00:2'b0)|
    (((_reg_2|_net_149))?_add_all_x_sg_out331:2'b0);
   assign  sg332 = ((_net_1418)?2'b00:2'b0)|
    (((_reg_2|_net_148))?_add_all_x_sg_out332:2'b0);
   assign  sg333 = ((_net_1417)?2'b00:2'b0)|
    (((_reg_2|_net_147))?_add_all_x_sg_out333:2'b0);
   assign  sg334 = ((_net_1416)?2'b00:2'b0)|
    (((_reg_2|_net_146))?_add_all_x_sg_out334:2'b0);
   assign  sg335 = ((_net_1415)?2'b00:2'b0)|
    (((_reg_2|_net_145))?_add_all_x_sg_out335:2'b0);
   assign  sg336 = ((_net_1414)?2'b00:2'b0)|
    (((_reg_2|_net_144))?_add_all_x_sg_out336:2'b0);
   assign  sg337 = ((_net_1413)?2'b00:2'b0)|
    (((_reg_2|_net_143))?_add_all_x_sg_out337:2'b0);
   assign  sg338 = ((_net_1412)?2'b00:2'b0)|
    (((_reg_2|_net_142))?_add_all_x_sg_out338:2'b0);
   assign  sg339 = ((_net_1411)?2'b00:2'b0)|
    (((_reg_2|_net_141))?_add_all_x_sg_out339:2'b0);
   assign  sg340 = ((_net_1410)?2'b00:2'b0)|
    (((_reg_2|_net_140))?_add_all_x_sg_out340:2'b0);
   assign  sg341 = ((_net_1409)?2'b00:2'b0)|
    (((_reg_2|_net_139))?_add_all_x_sg_out341:2'b0);
   assign  sg342 = ((_net_1408)?2'b00:2'b0)|
    (((_reg_2|_net_138))?_add_all_x_sg_out342:2'b0);
   assign  sg343 = ((_net_1407)?2'b00:2'b0)|
    (((_reg_2|_net_137))?_add_all_x_sg_out343:2'b0);
   assign  sg344 = ((_net_1406)?2'b00:2'b0)|
    (((_reg_2|_net_136))?_add_all_x_sg_out344:2'b0);
   assign  sg345 = ((_net_1405)?2'b00:2'b0)|
    (((_reg_2|_net_135))?_add_all_x_sg_out345:2'b0);
   assign  sg346 = ((_net_1404)?2'b00:2'b0)|
    (((_reg_2|_net_134))?_add_all_x_sg_out346:2'b0);
   assign  sg347 = ((_net_1403)?2'b00:2'b0)|
    (((_reg_2|_net_133))?_add_all_x_sg_out347:2'b0);
   assign  sg348 = ((_net_1402)?2'b00:2'b0)|
    (((_reg_2|_net_132))?_add_all_x_sg_out348:2'b0);
   assign  sg349 = ((_net_1401)?2'b00:2'b0)|
    (((_reg_2|_net_131))?_add_all_x_sg_out349:2'b0);
   assign  sg350 = ((_net_1400)?2'b00:10'b0)|
    (((_reg_2|_net_130))?_add_all_x_sg_out350:10'b0);
   assign  sg353 = ((_net_1399)?2'b00:2'b0)|
    (((_reg_2|_net_129))?_add_all_x_sg_out353:2'b0);
   assign  sg354 = ((_net_1398)?2'b00:2'b0)|
    (((_reg_2|_net_128))?_add_all_x_sg_out354:2'b0);
   assign  sg355 = ((_net_1397)?2'b00:2'b0)|
    (((_reg_2|_net_127))?_add_all_x_sg_out355:2'b0);
   assign  sg356 = ((_net_1396)?2'b00:2'b0)|
    (((_reg_2|_net_126))?_add_all_x_sg_out356:2'b0);
   assign  sg357 = ((_net_1395)?2'b00:2'b0)|
    (((_reg_2|_net_125))?_add_all_x_sg_out357:2'b0);
   assign  sg358 = ((_net_1394)?2'b00:2'b0)|
    (((_reg_2|_net_124))?_add_all_x_sg_out358:2'b0);
   assign  sg359 = ((_net_1393)?2'b00:2'b0)|
    (((_reg_2|_net_123))?_add_all_x_sg_out359:2'b0);
   assign  sg360 = ((_net_1392)?2'b00:2'b0)|
    (((_reg_2|_net_122))?_add_all_x_sg_out360:2'b0);
   assign  sg361 = ((_net_1391)?2'b00:2'b0)|
    (((_reg_2|_net_121))?_add_all_x_sg_out361:2'b0);
   assign  sg362 = ((_net_1390)?2'b00:2'b0)|
    (((_reg_2|_net_120))?_add_all_x_sg_out362:2'b0);
   assign  sg363 = ((_net_1389)?2'b00:2'b0)|
    (((_reg_2|_net_119))?_add_all_x_sg_out363:2'b0);
   assign  sg364 = ((_net_1388)?2'b00:2'b0)|
    (((_reg_2|_net_118))?_add_all_x_sg_out364:2'b0);
   assign  sg365 = ((_net_1387)?2'b00:2'b0)|
    (((_reg_2|_net_117))?_add_all_x_sg_out365:2'b0);
   assign  sg366 = ((_net_1386)?2'b00:2'b0)|
    (((_reg_2|_net_116))?_add_all_x_sg_out366:2'b0);
   assign  sg367 = ((_net_1385)?2'b00:2'b0)|
    (((_reg_2|_net_115))?_add_all_x_sg_out367:2'b0);
   assign  sg368 = ((_net_1384)?2'b00:2'b0)|
    (((_reg_2|_net_114))?_add_all_x_sg_out368:2'b0);
   assign  sg369 = ((_net_1383)?2'b00:2'b0)|
    (((_reg_2|_net_113))?_add_all_x_sg_out369:2'b0);
   assign  sg370 = ((_net_1382)?2'b00:2'b0)|
    (((_reg_2|_net_112))?_add_all_x_sg_out370:2'b0);
   assign  sg371 = ((_net_1381)?2'b00:2'b0)|
    (((_reg_2|_net_111))?_add_all_x_sg_out371:2'b0);
   assign  sg372 = ((_net_1380)?2'b00:2'b0)|
    (((_reg_2|_net_110))?_add_all_x_sg_out372:2'b0);
   assign  sg373 = ((_net_1379)?2'b00:2'b0)|
    (((_reg_2|_net_109))?_add_all_x_sg_out373:2'b0);
   assign  sg374 = ((_net_1378)?2'b00:2'b0)|
    (((_reg_2|_net_108))?_add_all_x_sg_out374:2'b0);
   assign  sg375 = ((_net_1377)?2'b00:2'b0)|
    (((_reg_2|_net_107))?_add_all_x_sg_out375:2'b0);
   assign  sg376 = ((_net_1376)?2'b00:2'b0)|
    (((_reg_2|_net_106))?_add_all_x_sg_out376:2'b0);
   assign  sg377 = ((_net_1375)?2'b00:2'b0)|
    (((_reg_2|_net_105))?_add_all_x_sg_out377:2'b0);
   assign  sg378 = ((_net_1374)?2'b00:2'b0)|
    (((_reg_2|_net_104))?_add_all_x_sg_out378:2'b0);
   assign  sg379 = ((_net_1373)?2'b00:2'b0)|
    (((_reg_2|_net_103))?_add_all_x_sg_out379:2'b0);
   assign  sg380 = ((_net_1372)?2'b00:2'b0)|
    (((_reg_2|_net_102))?_add_all_x_sg_out380:2'b0);
   assign  sg381 = ((_net_1371)?2'b00:2'b0)|
    (((_reg_2|_net_101))?_add_all_x_sg_out381:2'b0);
   assign  sg382 = ((_net_1370)?2'b00:10'b0)|
    (((_reg_2|_net_100))?_add_all_x_sg_out382:10'b0);
   assign  sg385 = ((_net_1369)?2'b00:2'b0)|
    (((_reg_2|_net_99))?_add_all_x_sg_out385:2'b0);
   assign  sg386 = ((_net_1368)?2'b00:2'b0)|
    (((_reg_2|_net_98))?_add_all_x_sg_out386:2'b0);
   assign  sg387 = ((_net_1367)?2'b00:2'b0)|
    (((_reg_2|_net_97))?_add_all_x_sg_out387:2'b0);
   assign  sg388 = ((_net_1366)?2'b00:2'b0)|
    (((_reg_2|_net_96))?_add_all_x_sg_out388:2'b0);
   assign  sg389 = ((_net_1365)?2'b00:2'b0)|
    (((_reg_2|_net_95))?_add_all_x_sg_out389:2'b0);
   assign  sg390 = ((_net_1364)?2'b00:2'b0)|
    (((_reg_2|_net_94))?_add_all_x_sg_out390:2'b0);
   assign  sg391 = ((_net_1363)?2'b00:2'b0)|
    (((_reg_2|_net_93))?_add_all_x_sg_out391:2'b0);
   assign  sg392 = ((_net_1362)?2'b00:2'b0)|
    (((_reg_2|_net_92))?_add_all_x_sg_out392:2'b0);
   assign  sg393 = ((_net_1361)?2'b00:2'b0)|
    (((_reg_2|_net_91))?_add_all_x_sg_out393:2'b0);
   assign  sg394 = ((_net_1360)?2'b00:2'b0)|
    (((_reg_2|_net_90))?_add_all_x_sg_out394:2'b0);
   assign  sg395 = ((_net_1359)?2'b00:2'b0)|
    (((_reg_2|_net_89))?_add_all_x_sg_out395:2'b0);
   assign  sg396 = ((_net_1358)?2'b00:2'b0)|
    (((_reg_2|_net_88))?_add_all_x_sg_out396:2'b0);
   assign  sg397 = ((_net_1357)?2'b00:2'b0)|
    (((_reg_2|_net_87))?_add_all_x_sg_out397:2'b0);
   assign  sg398 = ((_net_1356)?2'b00:2'b0)|
    (((_reg_2|_net_86))?_add_all_x_sg_out398:2'b0);
   assign  sg399 = ((_net_1355)?2'b00:2'b0)|
    (((_reg_2|_net_85))?_add_all_x_sg_out399:2'b0);
   assign  sg400 = ((_net_1354)?2'b00:2'b0)|
    (((_reg_2|_net_84))?_add_all_x_sg_out400:2'b0);
   assign  sg401 = ((_net_1353)?2'b00:2'b0)|
    (((_reg_2|_net_83))?_add_all_x_sg_out401:2'b0);
   assign  sg402 = ((_net_1352)?2'b00:2'b0)|
    (((_reg_2|_net_82))?_add_all_x_sg_out402:2'b0);
   assign  sg403 = ((_net_1351)?2'b00:2'b0)|
    (((_reg_2|_net_81))?_add_all_x_sg_out403:2'b0);
   assign  sg404 = ((_net_1350)?2'b00:2'b0)|
    (((_reg_2|_net_80))?_add_all_x_sg_out404:2'b0);
   assign  sg405 = ((_net_1349)?2'b00:2'b0)|
    (((_reg_2|_net_79))?_add_all_x_sg_out405:2'b0);
   assign  sg406 = ((_net_1348)?2'b00:2'b0)|
    (((_reg_2|_net_78))?_add_all_x_sg_out406:2'b0);
   assign  sg407 = ((_net_1347)?2'b00:2'b0)|
    (((_reg_2|_net_77))?_add_all_x_sg_out407:2'b0);
   assign  sg408 = ((_net_1346)?2'b00:2'b0)|
    (((_reg_2|_net_76))?_add_all_x_sg_out408:2'b0);
   assign  sg409 = ((_net_1345)?2'b00:2'b0)|
    (((_reg_2|_net_75))?_add_all_x_sg_out409:2'b0);
   assign  sg410 = ((_net_1344)?2'b00:2'b0)|
    (((_reg_2|_net_74))?_add_all_x_sg_out410:2'b0);
   assign  sg411 = ((_net_1343)?2'b00:2'b0)|
    (((_reg_2|_net_73))?_add_all_x_sg_out411:2'b0);
   assign  sg412 = ((_net_1342)?2'b00:2'b0)|
    (((_reg_2|_net_72))?_add_all_x_sg_out412:2'b0);
   assign  sg413 = ((_net_1341)?2'b00:2'b0)|
    (((_reg_2|_net_71))?_add_all_x_sg_out413:2'b0);
   assign  sg414 = ((_net_1340)?2'b00:10'b0)|
    (((_reg_2|_net_70))?_add_all_x_sg_out414:10'b0);
   assign  sg417 = ((_net_1339)?2'b00:2'b0)|
    (((_reg_2|_net_69))?_add_all_x_sg_out417:2'b0);
   assign  sg418 = ((_net_1338)?2'b00:2'b0)|
    (((_reg_2|_net_68))?_add_all_x_sg_out418:2'b0);
   assign  sg419 = ((_net_1337)?2'b00:2'b0)|
    (((_reg_2|_net_67))?_add_all_x_sg_out419:2'b0);
   assign  sg420 = ((_net_1336)?2'b00:2'b0)|
    (((_reg_2|_net_66))?_add_all_x_sg_out420:2'b0);
   assign  sg421 = ((_net_1335)?2'b00:2'b0)|
    (((_reg_2|_net_65))?_add_all_x_sg_out421:2'b0);
   assign  sg422 = ((_net_1334)?2'b00:2'b0)|
    (((_reg_2|_net_64))?_add_all_x_sg_out422:2'b0);
   assign  sg423 = ((_net_1333)?2'b00:2'b0)|
    (((_reg_2|_net_63))?_add_all_x_sg_out423:2'b0);
   assign  sg424 = ((_net_1332)?2'b00:2'b0)|
    (((_reg_2|_net_62))?_add_all_x_sg_out424:2'b0);
   assign  sg425 = ((_net_1331)?2'b00:2'b0)|
    (((_reg_2|_net_61))?_add_all_x_sg_out425:2'b0);
   assign  sg426 = ((_net_1330)?2'b00:2'b0)|
    (((_reg_2|_net_60))?_add_all_x_sg_out426:2'b0);
   assign  sg427 = ((_net_1329)?2'b00:2'b0)|
    (((_reg_2|_net_59))?_add_all_x_sg_out427:2'b0);
   assign  sg428 = ((_net_1328)?2'b00:2'b0)|
    (((_reg_2|_net_58))?_add_all_x_sg_out428:2'b0);
   assign  sg429 = ((_net_1327)?2'b00:2'b0)|
    (((_reg_2|_net_57))?_add_all_x_sg_out429:2'b0);
   assign  sg430 = ((_net_1326)?2'b00:2'b0)|
    (((_reg_2|_net_56))?_add_all_x_sg_out430:2'b0);
   assign  sg431 = ((_net_1325)?2'b00:2'b0)|
    (((_reg_2|_net_55))?_add_all_x_sg_out431:2'b0);
   assign  sg432 = ((_net_1324)?2'b00:2'b0)|
    (((_reg_2|_net_54))?_add_all_x_sg_out432:2'b0);
   assign  sg433 = ((_net_1323)?2'b00:2'b0)|
    (((_reg_2|_net_53))?_add_all_x_sg_out433:2'b0);
   assign  sg434 = ((_net_1322)?2'b00:2'b0)|
    (((_reg_2|_net_52))?_add_all_x_sg_out434:2'b0);
   assign  sg435 = ((_net_1321)?2'b00:2'b0)|
    (((_reg_2|_net_51))?_add_all_x_sg_out435:2'b0);
   assign  sg436 = ((_net_1320)?2'b00:2'b0)|
    (((_reg_2|_net_50))?_add_all_x_sg_out436:2'b0);
   assign  sg437 = ((_net_1319)?2'b00:2'b0)|
    (((_reg_2|_net_49))?_add_all_x_sg_out437:2'b0);
   assign  sg438 = ((_net_1318)?2'b00:2'b0)|
    (((_reg_2|_net_48))?_add_all_x_sg_out438:2'b0);
   assign  sg439 = ((_net_1317)?2'b00:2'b0)|
    (((_reg_2|_net_47))?_add_all_x_sg_out439:2'b0);
   assign  sg440 = ((_net_1316)?2'b00:2'b0)|
    (((_reg_2|_net_46))?_add_all_x_sg_out440:2'b0);
   assign  sg441 = ((_net_1315)?2'b00:2'b0)|
    (((_reg_2|_net_45))?_add_all_x_sg_out441:2'b0);
   assign  sg442 = ((_net_1314)?2'b00:2'b0)|
    (((_reg_2|_net_44))?_add_all_x_sg_out442:2'b0);
   assign  sg443 = ((_net_1313)?2'b00:2'b0)|
    (((_reg_2|_net_43))?_add_all_x_sg_out443:2'b0);
   assign  sg444 = ((_net_1312)?2'b00:2'b0)|
    (((_reg_2|_net_42))?_add_all_x_sg_out444:2'b0);
   assign  sg445 = ((_net_1311)?2'b00:2'b0)|
    (((_reg_2|_net_41))?_add_all_x_sg_out445:2'b0);
   assign  sg446 = ((_net_1310)?2'b00:10'b0)|
    (((_reg_2|_net_40))?_add_all_x_sg_out446:10'b0);
   assign  sg449 = ((_net_1309)?2'b00:2'b0)|
    (((_reg_2|_net_39))?_add_all_x_sg_out449:2'b0);
   assign  sg450 = ((_net_1308)?2'b00:2'b0)|
    (((_reg_2|_net_38))?_add_all_x_sg_out450:2'b0);
   assign  sg451 = ((_net_1307)?2'b00:2'b0)|
    (((_reg_2|_net_37))?_add_all_x_sg_out451:2'b0);
   assign  sg452 = ((_net_1306)?2'b00:2'b0)|
    (((_reg_2|_net_36))?_add_all_x_sg_out452:2'b0);
   assign  sg453 = ((_net_1305)?2'b00:2'b0)|
    (((_reg_2|_net_35))?_add_all_x_sg_out453:2'b0);
   assign  sg454 = ((_net_1304)?2'b00:2'b0)|
    (((_reg_2|_net_34))?_add_all_x_sg_out454:2'b0);
   assign  sg455 = ((_net_1303)?2'b00:2'b0)|
    (((_reg_2|_net_33))?_add_all_x_sg_out455:2'b0);
   assign  sg456 = ((_net_1302)?2'b00:2'b0)|
    (((_reg_2|_net_32))?_add_all_x_sg_out456:2'b0);
   assign  sg457 = ((_net_1301)?2'b00:2'b0)|
    (((_reg_2|_net_31))?_add_all_x_sg_out457:2'b0);
   assign  sg458 = ((_net_1300)?2'b00:2'b0)|
    (((_reg_2|_net_30))?_add_all_x_sg_out458:2'b0);
   assign  sg459 = ((_net_1299)?2'b00:2'b0)|
    (((_reg_2|_net_29))?_add_all_x_sg_out459:2'b0);
   assign  sg460 = ((_net_1298)?2'b00:2'b0)|
    (((_reg_2|_net_28))?_add_all_x_sg_out460:2'b0);
   assign  sg461 = ((_net_1297)?2'b00:2'b0)|
    (((_reg_2|_net_27))?_add_all_x_sg_out461:2'b0);
   assign  sg462 = ((_net_1296)?2'b00:2'b0)|
    (((_reg_2|_net_26))?_add_all_x_sg_out462:2'b0);
   assign  sg463 = ((_net_1295)?2'b00:2'b0)|
    (((_reg_2|_net_25))?_add_all_x_sg_out463:2'b0);
   assign  sg464 = ((_net_1294)?2'b00:2'b0)|
    (((_reg_2|_net_24))?_add_all_x_sg_out464:2'b0);
   assign  sg465 = ((_net_1293)?2'b00:2'b0)|
    (((_reg_2|_net_23))?_add_all_x_sg_out465:2'b0);
   assign  sg466 = ((_net_1292)?2'b00:2'b0)|
    (((_reg_2|_net_22))?_add_all_x_sg_out466:2'b0);
   assign  sg467 = ((_net_1291)?2'b00:2'b0)|
    (((_reg_2|_net_21))?_add_all_x_sg_out467:2'b0);
   assign  sg468 = ((_net_1290)?2'b00:2'b0)|
    (((_reg_2|_net_20))?_add_all_x_sg_out468:2'b0);
   assign  sg469 = ((_net_1289)?2'b00:2'b0)|
    (((_reg_2|_net_19))?_add_all_x_sg_out469:2'b0);
   assign  sg470 = ((_net_1288)?2'b00:2'b0)|
    (((_reg_2|_net_18))?_add_all_x_sg_out470:2'b0);
   assign  sg471 = ((_net_1287)?2'b00:2'b0)|
    (((_reg_2|_net_17))?_add_all_x_sg_out471:2'b0);
   assign  sg472 = ((_net_1286)?2'b00:2'b0)|
    (((_reg_2|_net_16))?_add_all_x_sg_out472:2'b0);
   assign  sg473 = ((_net_1285)?2'b00:2'b0)|
    (((_reg_2|_net_15))?_add_all_x_sg_out473:2'b0);
   assign  sg474 = ((_net_1284)?2'b00:2'b0)|
    (((_reg_2|_net_14))?_add_all_x_sg_out474:2'b0);
   assign  sg475 = ((_net_1283)?2'b00:2'b0)|
    (((_reg_2|_net_13))?_add_all_x_sg_out475:2'b0);
   assign  sg476 = ((_net_1282)?2'b00:2'b0)|
    (((_reg_2|_net_12))?_add_all_x_sg_out476:2'b0);
   assign  sg477 = ((_net_1281)?2'b00:2'b0)|
    (((_reg_2|_net_11))?_add_all_x_sg_out477:2'b0);
   assign  sg478 = ((_net_1280)?2'b00:2'b0)|
    (((_reg_2|_net_10))?_add_all_x_sg_out478:2'b0);
   assign  kanwa_s = (_net_1275|(_reg_2|_net_5));
   assign  _add_all_x_sig = even_w1;
   assign  _add_all_x_start = start_wire;
   assign  _add_all_x_goal = goal_wire;
   assign  _add_all_x_dig_w = wall_w;
   assign  _add_all_x_data_in33 = data_wire33;
   assign  _add_all_x_data_in34 = data_wire34;
   assign  _add_all_x_data_in35 = data_wire35;
   assign  _add_all_x_data_in36 = data_wire36;
   assign  _add_all_x_data_in37 = data_wire37;
   assign  _add_all_x_data_in38 = data_wire38;
   assign  _add_all_x_data_in39 = data_wire39;
   assign  _add_all_x_data_in40 = data_wire40;
   assign  _add_all_x_data_in41 = data_wire41;
   assign  _add_all_x_data_in42 = data_wire42;
   assign  _add_all_x_data_in43 = data_wire43;
   assign  _add_all_x_data_in44 = data_wire44;
   assign  _add_all_x_data_in45 = data_wire45;
   assign  _add_all_x_data_in46 = data_wire46;
   assign  _add_all_x_data_in47 = data_wire47;
   assign  _add_all_x_data_in48 = data_wire48;
   assign  _add_all_x_data_in49 = data_wire49;
   assign  _add_all_x_data_in50 = data_wire50;
   assign  _add_all_x_data_in51 = data_wire51;
   assign  _add_all_x_data_in52 = data_wire52;
   assign  _add_all_x_data_in53 = data_wire53;
   assign  _add_all_x_data_in54 = data_wire54;
   assign  _add_all_x_data_in55 = data_wire55;
   assign  _add_all_x_data_in56 = data_wire56;
   assign  _add_all_x_data_in57 = data_wire57;
   assign  _add_all_x_data_in58 = data_wire58;
   assign  _add_all_x_data_in59 = data_wire59;
   assign  _add_all_x_data_in60 = data_wire60;
   assign  _add_all_x_data_in61 = data_wire61;
   assign  _add_all_x_data_in62 = data_wire62;
   assign  _add_all_x_data_in65 = data_wire65;
   assign  _add_all_x_data_in66 = data_wire66;
   assign  _add_all_x_data_in67 = data_wire67;
   assign  _add_all_x_data_in68 = data_wire68;
   assign  _add_all_x_data_in69 = data_wire69;
   assign  _add_all_x_data_in70 = data_wire70;
   assign  _add_all_x_data_in71 = data_wire71;
   assign  _add_all_x_data_in72 = data_wire72;
   assign  _add_all_x_data_in73 = data_wire73;
   assign  _add_all_x_data_in74 = data_wire74;
   assign  _add_all_x_data_in75 = data_wire75;
   assign  _add_all_x_data_in76 = data_wire76;
   assign  _add_all_x_data_in77 = data_wire77;
   assign  _add_all_x_data_in78 = data_wire78;
   assign  _add_all_x_data_in79 = data_wire79;
   assign  _add_all_x_data_in80 = data_wire80;
   assign  _add_all_x_data_in81 = data_wire81;
   assign  _add_all_x_data_in82 = data_wire82;
   assign  _add_all_x_data_in83 = data_wire83;
   assign  _add_all_x_data_in84 = data_wire84;
   assign  _add_all_x_data_in85 = data_wire85;
   assign  _add_all_x_data_in86 = data_wire86;
   assign  _add_all_x_data_in87 = data_wire87;
   assign  _add_all_x_data_in88 = data_wire88;
   assign  _add_all_x_data_in89 = data_wire89;
   assign  _add_all_x_data_in90 = data_wire90;
   assign  _add_all_x_data_in91 = data_wire91;
   assign  _add_all_x_data_in92 = data_wire92;
   assign  _add_all_x_data_in93 = data_wire93;
   assign  _add_all_x_data_in94 = data_wire94;
   assign  _add_all_x_data_in97 = data_wire97;
   assign  _add_all_x_data_in98 = data_wire98;
   assign  _add_all_x_data_in99 = data_wire99;
   assign  _add_all_x_data_in100 = data_wire100;
   assign  _add_all_x_data_in101 = data_wire101;
   assign  _add_all_x_data_in102 = data_wire102;
   assign  _add_all_x_data_in103 = data_wire103;
   assign  _add_all_x_data_in104 = data_wire104;
   assign  _add_all_x_data_in105 = data_wire105;
   assign  _add_all_x_data_in106 = data_wire106;
   assign  _add_all_x_data_in107 = data_wire107;
   assign  _add_all_x_data_in108 = data_wire108;
   assign  _add_all_x_data_in109 = data_wire109;
   assign  _add_all_x_data_in110 = data_wire110;
   assign  _add_all_x_data_in111 = data_wire111;
   assign  _add_all_x_data_in112 = data_wire112;
   assign  _add_all_x_data_in113 = data_wire113;
   assign  _add_all_x_data_in114 = data_wire114;
   assign  _add_all_x_data_in115 = data_wire115;
   assign  _add_all_x_data_in116 = data_wire116;
   assign  _add_all_x_data_in117 = data_wire117;
   assign  _add_all_x_data_in118 = data_wire118;
   assign  _add_all_x_data_in119 = data_wire119;
   assign  _add_all_x_data_in120 = data_wire120;
   assign  _add_all_x_data_in121 = data_wire121;
   assign  _add_all_x_data_in122 = data_wire122;
   assign  _add_all_x_data_in123 = data_wire123;
   assign  _add_all_x_data_in124 = data_wire124;
   assign  _add_all_x_data_in125 = data_wire125;
   assign  _add_all_x_data_in126 = data_wire126;
   assign  _add_all_x_data_in129 = data_wire129;
   assign  _add_all_x_data_in130 = data_wire130;
   assign  _add_all_x_data_in131 = data_wire131;
   assign  _add_all_x_data_in132 = data_wire132;
   assign  _add_all_x_data_in133 = data_wire133;
   assign  _add_all_x_data_in134 = data_wire134;
   assign  _add_all_x_data_in135 = data_wire135;
   assign  _add_all_x_data_in136 = data_wire136;
   assign  _add_all_x_data_in137 = data_wire137;
   assign  _add_all_x_data_in138 = data_wire138;
   assign  _add_all_x_data_in139 = data_wire139;
   assign  _add_all_x_data_in140 = data_wire140;
   assign  _add_all_x_data_in141 = data_wire141;
   assign  _add_all_x_data_in142 = data_wire142;
   assign  _add_all_x_data_in143 = data_wire143;
   assign  _add_all_x_data_in144 = data_wire144;
   assign  _add_all_x_data_in145 = data_wire145;
   assign  _add_all_x_data_in146 = data_wire146;
   assign  _add_all_x_data_in147 = data_wire147;
   assign  _add_all_x_data_in148 = data_wire148;
   assign  _add_all_x_data_in149 = data_wire149;
   assign  _add_all_x_data_in150 = data_wire150;
   assign  _add_all_x_data_in151 = data_wire151;
   assign  _add_all_x_data_in152 = data_wire152;
   assign  _add_all_x_data_in153 = data_wire153;
   assign  _add_all_x_data_in154 = data_wire154;
   assign  _add_all_x_data_in155 = data_wire155;
   assign  _add_all_x_data_in156 = data_wire156;
   assign  _add_all_x_data_in157 = data_wire157;
   assign  _add_all_x_data_in158 = data_wire158;
   assign  _add_all_x_data_in161 = data_wire161;
   assign  _add_all_x_data_in162 = data_wire162;
   assign  _add_all_x_data_in163 = data_wire163;
   assign  _add_all_x_data_in164 = data_wire164;
   assign  _add_all_x_data_in165 = data_wire165;
   assign  _add_all_x_data_in166 = data_wire166;
   assign  _add_all_x_data_in167 = data_wire167;
   assign  _add_all_x_data_in168 = data_wire168;
   assign  _add_all_x_data_in169 = data_wire169;
   assign  _add_all_x_data_in170 = data_wire170;
   assign  _add_all_x_data_in171 = data_wire171;
   assign  _add_all_x_data_in172 = data_wire172;
   assign  _add_all_x_data_in173 = data_wire173;
   assign  _add_all_x_data_in174 = data_wire174;
   assign  _add_all_x_data_in175 = data_wire175;
   assign  _add_all_x_data_in176 = data_wire176;
   assign  _add_all_x_data_in177 = data_wire177;
   assign  _add_all_x_data_in178 = data_wire178;
   assign  _add_all_x_data_in179 = data_wire179;
   assign  _add_all_x_data_in180 = data_wire180;
   assign  _add_all_x_data_in181 = data_wire181;
   assign  _add_all_x_data_in182 = data_wire182;
   assign  _add_all_x_data_in183 = data_wire183;
   assign  _add_all_x_data_in184 = data_wire184;
   assign  _add_all_x_data_in185 = data_wire185;
   assign  _add_all_x_data_in186 = data_wire186;
   assign  _add_all_x_data_in187 = data_wire187;
   assign  _add_all_x_data_in188 = data_wire188;
   assign  _add_all_x_data_in189 = data_wire189;
   assign  _add_all_x_data_in190 = data_wire190;
   assign  _add_all_x_data_in193 = data_wire193;
   assign  _add_all_x_data_in194 = data_wire194;
   assign  _add_all_x_data_in195 = data_wire195;
   assign  _add_all_x_data_in196 = data_wire196;
   assign  _add_all_x_data_in197 = data_wire197;
   assign  _add_all_x_data_in198 = data_wire198;
   assign  _add_all_x_data_in199 = data_wire199;
   assign  _add_all_x_data_in200 = data_wire200;
   assign  _add_all_x_data_in201 = data_wire201;
   assign  _add_all_x_data_in202 = data_wire202;
   assign  _add_all_x_data_in203 = data_wire203;
   assign  _add_all_x_data_in204 = data_wire204;
   assign  _add_all_x_data_in205 = data_wire205;
   assign  _add_all_x_data_in206 = data_wire206;
   assign  _add_all_x_data_in207 = data_wire207;
   assign  _add_all_x_data_in208 = data_wire208;
   assign  _add_all_x_data_in209 = data_wire209;
   assign  _add_all_x_data_in210 = data_wire210;
   assign  _add_all_x_data_in211 = data_wire211;
   assign  _add_all_x_data_in212 = data_wire212;
   assign  _add_all_x_data_in213 = data_wire213;
   assign  _add_all_x_data_in214 = data_wire214;
   assign  _add_all_x_data_in215 = data_wire215;
   assign  _add_all_x_data_in216 = data_wire216;
   assign  _add_all_x_data_in217 = data_wire217;
   assign  _add_all_x_data_in218 = data_wire218;
   assign  _add_all_x_data_in219 = data_wire219;
   assign  _add_all_x_data_in220 = data_wire220;
   assign  _add_all_x_data_in221 = data_wire221;
   assign  _add_all_x_data_in222 = data_wire222;
   assign  _add_all_x_data_in225 = data_wire225;
   assign  _add_all_x_data_in226 = data_wire226;
   assign  _add_all_x_data_in227 = data_wire227;
   assign  _add_all_x_data_in228 = data_wire228;
   assign  _add_all_x_data_in229 = data_wire229;
   assign  _add_all_x_data_in230 = data_wire230;
   assign  _add_all_x_data_in231 = data_wire231;
   assign  _add_all_x_data_in232 = data_wire232;
   assign  _add_all_x_data_in233 = data_wire233;
   assign  _add_all_x_data_in234 = data_wire234;
   assign  _add_all_x_data_in235 = data_wire235;
   assign  _add_all_x_data_in236 = data_wire236;
   assign  _add_all_x_data_in237 = data_wire237;
   assign  _add_all_x_data_in238 = data_wire238;
   assign  _add_all_x_data_in239 = data_wire239;
   assign  _add_all_x_data_in240 = data_wire240;
   assign  _add_all_x_data_in241 = data_wire241;
   assign  _add_all_x_data_in242 = data_wire242;
   assign  _add_all_x_data_in243 = data_wire243;
   assign  _add_all_x_data_in244 = data_wire244;
   assign  _add_all_x_data_in245 = data_wire245;
   assign  _add_all_x_data_in246 = data_wire246;
   assign  _add_all_x_data_in247 = data_wire247;
   assign  _add_all_x_data_in248 = data_wire248;
   assign  _add_all_x_data_in249 = data_wire249;
   assign  _add_all_x_data_in250 = data_wire250;
   assign  _add_all_x_data_in251 = data_wire251;
   assign  _add_all_x_data_in252 = data_wire252;
   assign  _add_all_x_data_in253 = data_wire253;
   assign  _add_all_x_data_in254 = data_wire254;
   assign  _add_all_x_data_in257 = data_wire257;
   assign  _add_all_x_data_in258 = data_wire258;
   assign  _add_all_x_data_in259 = data_wire259;
   assign  _add_all_x_data_in260 = data_wire260;
   assign  _add_all_x_data_in261 = data_wire261;
   assign  _add_all_x_data_in262 = data_wire262;
   assign  _add_all_x_data_in263 = data_wire263;
   assign  _add_all_x_data_in264 = data_wire264;
   assign  _add_all_x_data_in265 = data_wire265;
   assign  _add_all_x_data_in266 = data_wire266;
   assign  _add_all_x_data_in267 = data_wire267;
   assign  _add_all_x_data_in268 = data_wire268;
   assign  _add_all_x_data_in269 = data_wire269;
   assign  _add_all_x_data_in270 = data_wire270;
   assign  _add_all_x_data_in271 = data_wire271;
   assign  _add_all_x_data_in272 = data_wire272;
   assign  _add_all_x_data_in273 = data_wire273;
   assign  _add_all_x_data_in274 = data_wire274;
   assign  _add_all_x_data_in275 = data_wire275;
   assign  _add_all_x_data_in276 = data_wire276;
   assign  _add_all_x_data_in277 = data_wire277;
   assign  _add_all_x_data_in278 = data_wire278;
   assign  _add_all_x_data_in279 = data_wire279;
   assign  _add_all_x_data_in280 = data_wire280;
   assign  _add_all_x_data_in281 = data_wire281;
   assign  _add_all_x_data_in282 = data_wire282;
   assign  _add_all_x_data_in283 = data_wire283;
   assign  _add_all_x_data_in284 = data_wire284;
   assign  _add_all_x_data_in285 = data_wire285;
   assign  _add_all_x_data_in286 = data_wire286;
   assign  _add_all_x_data_in289 = data_wire289;
   assign  _add_all_x_data_in290 = data_wire290;
   assign  _add_all_x_data_in291 = data_wire291;
   assign  _add_all_x_data_in292 = data_wire292;
   assign  _add_all_x_data_in293 = data_wire293;
   assign  _add_all_x_data_in294 = data_wire294;
   assign  _add_all_x_data_in295 = data_wire295;
   assign  _add_all_x_data_in296 = data_wire296;
   assign  _add_all_x_data_in297 = data_wire297;
   assign  _add_all_x_data_in298 = data_wire298;
   assign  _add_all_x_data_in299 = data_wire299;
   assign  _add_all_x_data_in300 = data_wire300;
   assign  _add_all_x_data_in301 = data_wire301;
   assign  _add_all_x_data_in302 = data_wire302;
   assign  _add_all_x_data_in303 = data_wire303;
   assign  _add_all_x_data_in304 = data_wire304;
   assign  _add_all_x_data_in305 = data_wire305;
   assign  _add_all_x_data_in306 = data_wire306;
   assign  _add_all_x_data_in307 = data_wire307;
   assign  _add_all_x_data_in308 = data_wire308;
   assign  _add_all_x_data_in309 = data_wire309;
   assign  _add_all_x_data_in310 = data_wire310;
   assign  _add_all_x_data_in311 = data_wire311;
   assign  _add_all_x_data_in312 = data_wire312;
   assign  _add_all_x_data_in313 = data_wire313;
   assign  _add_all_x_data_in314 = data_wire314;
   assign  _add_all_x_data_in315 = data_wire315;
   assign  _add_all_x_data_in316 = data_wire316;
   assign  _add_all_x_data_in317 = data_wire317;
   assign  _add_all_x_data_in318 = data_wire318;
   assign  _add_all_x_data_in321 = data_wire321;
   assign  _add_all_x_data_in322 = data_wire322;
   assign  _add_all_x_data_in323 = data_wire323;
   assign  _add_all_x_data_in324 = data_wire324;
   assign  _add_all_x_data_in325 = data_wire325;
   assign  _add_all_x_data_in326 = data_wire326;
   assign  _add_all_x_data_in327 = data_wire327;
   assign  _add_all_x_data_in328 = data_wire328;
   assign  _add_all_x_data_in329 = data_wire329;
   assign  _add_all_x_data_in330 = data_wire330;
   assign  _add_all_x_data_in331 = data_wire331;
   assign  _add_all_x_data_in332 = data_wire332;
   assign  _add_all_x_data_in333 = data_wire333;
   assign  _add_all_x_data_in334 = data_wire334;
   assign  _add_all_x_data_in335 = data_wire335;
   assign  _add_all_x_data_in336 = data_wire336;
   assign  _add_all_x_data_in337 = data_wire337;
   assign  _add_all_x_data_in338 = data_wire338;
   assign  _add_all_x_data_in339 = data_wire339;
   assign  _add_all_x_data_in340 = data_wire340;
   assign  _add_all_x_data_in341 = data_wire341;
   assign  _add_all_x_data_in342 = data_wire342;
   assign  _add_all_x_data_in343 = data_wire343;
   assign  _add_all_x_data_in344 = data_wire344;
   assign  _add_all_x_data_in345 = data_wire345;
   assign  _add_all_x_data_in346 = data_wire346;
   assign  _add_all_x_data_in347 = data_wire347;
   assign  _add_all_x_data_in348 = data_wire348;
   assign  _add_all_x_data_in349 = data_wire349;
   assign  _add_all_x_data_in350 = data_wire350;
   assign  _add_all_x_data_in353 = data_wire353;
   assign  _add_all_x_data_in354 = data_wire354;
   assign  _add_all_x_data_in355 = data_wire355;
   assign  _add_all_x_data_in356 = data_wire356;
   assign  _add_all_x_data_in357 = data_wire357;
   assign  _add_all_x_data_in358 = data_wire358;
   assign  _add_all_x_data_in359 = data_wire359;
   assign  _add_all_x_data_in360 = data_wire360;
   assign  _add_all_x_data_in361 = data_wire361;
   assign  _add_all_x_data_in362 = data_wire362;
   assign  _add_all_x_data_in363 = data_wire363;
   assign  _add_all_x_data_in364 = data_wire364;
   assign  _add_all_x_data_in365 = data_wire365;
   assign  _add_all_x_data_in366 = data_wire366;
   assign  _add_all_x_data_in367 = data_wire367;
   assign  _add_all_x_data_in368 = data_wire368;
   assign  _add_all_x_data_in369 = data_wire369;
   assign  _add_all_x_data_in370 = data_wire370;
   assign  _add_all_x_data_in371 = data_wire371;
   assign  _add_all_x_data_in372 = data_wire372;
   assign  _add_all_x_data_in373 = data_wire373;
   assign  _add_all_x_data_in374 = data_wire374;
   assign  _add_all_x_data_in375 = data_wire375;
   assign  _add_all_x_data_in376 = data_wire376;
   assign  _add_all_x_data_in377 = data_wire377;
   assign  _add_all_x_data_in378 = data_wire378;
   assign  _add_all_x_data_in379 = data_wire379;
   assign  _add_all_x_data_in380 = data_wire380;
   assign  _add_all_x_data_in381 = data_wire381;
   assign  _add_all_x_data_in382 = data_wire382;
   assign  _add_all_x_data_in385 = data_wire385;
   assign  _add_all_x_data_in386 = data_wire386;
   assign  _add_all_x_data_in387 = data_wire387;
   assign  _add_all_x_data_in388 = data_wire388;
   assign  _add_all_x_data_in389 = data_wire389;
   assign  _add_all_x_data_in390 = data_wire390;
   assign  _add_all_x_data_in391 = data_wire391;
   assign  _add_all_x_data_in392 = data_wire392;
   assign  _add_all_x_data_in393 = data_wire393;
   assign  _add_all_x_data_in394 = data_wire394;
   assign  _add_all_x_data_in395 = data_wire395;
   assign  _add_all_x_data_in396 = data_wire396;
   assign  _add_all_x_data_in397 = data_wire397;
   assign  _add_all_x_data_in398 = data_wire398;
   assign  _add_all_x_data_in399 = data_wire399;
   assign  _add_all_x_data_in400 = data_wire400;
   assign  _add_all_x_data_in401 = data_wire401;
   assign  _add_all_x_data_in402 = data_wire402;
   assign  _add_all_x_data_in403 = data_wire403;
   assign  _add_all_x_data_in404 = data_wire404;
   assign  _add_all_x_data_in405 = data_wire405;
   assign  _add_all_x_data_in406 = data_wire406;
   assign  _add_all_x_data_in407 = data_wire407;
   assign  _add_all_x_data_in408 = data_wire408;
   assign  _add_all_x_data_in409 = data_wire409;
   assign  _add_all_x_data_in410 = data_wire410;
   assign  _add_all_x_data_in411 = data_wire411;
   assign  _add_all_x_data_in412 = data_wire412;
   assign  _add_all_x_data_in413 = data_wire413;
   assign  _add_all_x_data_in414 = data_wire414;
   assign  _add_all_x_data_in417 = data_wire417;
   assign  _add_all_x_data_in418 = data_wire418;
   assign  _add_all_x_data_in419 = data_wire419;
   assign  _add_all_x_data_in420 = data_wire420;
   assign  _add_all_x_data_in421 = data_wire421;
   assign  _add_all_x_data_in422 = data_wire422;
   assign  _add_all_x_data_in423 = data_wire423;
   assign  _add_all_x_data_in424 = data_wire424;
   assign  _add_all_x_data_in425 = data_wire425;
   assign  _add_all_x_data_in426 = data_wire426;
   assign  _add_all_x_data_in427 = data_wire427;
   assign  _add_all_x_data_in428 = data_wire428;
   assign  _add_all_x_data_in429 = data_wire429;
   assign  _add_all_x_data_in430 = data_wire430;
   assign  _add_all_x_data_in431 = data_wire431;
   assign  _add_all_x_data_in432 = data_wire432;
   assign  _add_all_x_data_in433 = data_wire433;
   assign  _add_all_x_data_in434 = data_wire434;
   assign  _add_all_x_data_in435 = data_wire435;
   assign  _add_all_x_data_in436 = data_wire436;
   assign  _add_all_x_data_in437 = data_wire437;
   assign  _add_all_x_data_in438 = data_wire438;
   assign  _add_all_x_data_in439 = data_wire439;
   assign  _add_all_x_data_in440 = data_wire440;
   assign  _add_all_x_data_in441 = data_wire441;
   assign  _add_all_x_data_in442 = data_wire442;
   assign  _add_all_x_data_in443 = data_wire443;
   assign  _add_all_x_data_in444 = data_wire444;
   assign  _add_all_x_data_in445 = data_wire445;
   assign  _add_all_x_data_in446 = data_wire446;
   assign  _add_all_x_data_in449 = data_wire449;
   assign  _add_all_x_data_in450 = data_wire450;
   assign  _add_all_x_data_in451 = data_wire451;
   assign  _add_all_x_data_in452 = data_wire452;
   assign  _add_all_x_data_in453 = data_wire453;
   assign  _add_all_x_data_in454 = data_wire454;
   assign  _add_all_x_data_in455 = data_wire455;
   assign  _add_all_x_data_in456 = data_wire456;
   assign  _add_all_x_data_in457 = data_wire457;
   assign  _add_all_x_data_in458 = data_wire458;
   assign  _add_all_x_data_in459 = data_wire459;
   assign  _add_all_x_data_in460 = data_wire460;
   assign  _add_all_x_data_in461 = data_wire461;
   assign  _add_all_x_data_in462 = data_wire462;
   assign  _add_all_x_data_in463 = data_wire463;
   assign  _add_all_x_data_in464 = data_wire464;
   assign  _add_all_x_data_in465 = data_wire465;
   assign  _add_all_x_data_in466 = data_wire466;
   assign  _add_all_x_data_in467 = data_wire467;
   assign  _add_all_x_data_in468 = data_wire468;
   assign  _add_all_x_data_in469 = data_wire469;
   assign  _add_all_x_data_in470 = data_wire470;
   assign  _add_all_x_data_in471 = data_wire471;
   assign  _add_all_x_data_in472 = data_wire472;
   assign  _add_all_x_data_in473 = data_wire473;
   assign  _add_all_x_data_in474 = data_wire474;
   assign  _add_all_x_data_in475 = data_wire475;
   assign  _add_all_x_data_in476 = data_wire476;
   assign  _add_all_x_data_in477 = data_wire477;
   assign  _add_all_x_data_in478 = data_wire478;
   assign  _add_all_x_data_in_org33 = data_out_org33;
   assign  _add_all_x_data_in_org34 = data_out_org34;
   assign  _add_all_x_data_in_org35 = data_out_org35;
   assign  _add_all_x_data_in_org36 = data_out_org36;
   assign  _add_all_x_data_in_org37 = data_out_org37;
   assign  _add_all_x_data_in_org38 = data_out_org38;
   assign  _add_all_x_data_in_org39 = data_out_org39;
   assign  _add_all_x_data_in_org40 = data_out_org40;
   assign  _add_all_x_data_in_org41 = data_out_org41;
   assign  _add_all_x_data_in_org42 = data_out_org42;
   assign  _add_all_x_data_in_org43 = data_out_org43;
   assign  _add_all_x_data_in_org44 = data_out_org44;
   assign  _add_all_x_data_in_org45 = data_out_org45;
   assign  _add_all_x_data_in_org46 = data_out_org46;
   assign  _add_all_x_data_in_org47 = data_out_org47;
   assign  _add_all_x_data_in_org48 = data_out_org48;
   assign  _add_all_x_data_in_org49 = data_out_org49;
   assign  _add_all_x_data_in_org50 = data_out_org50;
   assign  _add_all_x_data_in_org51 = data_out_org51;
   assign  _add_all_x_data_in_org52 = data_out_org52;
   assign  _add_all_x_data_in_org53 = data_out_org53;
   assign  _add_all_x_data_in_org54 = data_out_org54;
   assign  _add_all_x_data_in_org55 = data_out_org55;
   assign  _add_all_x_data_in_org56 = data_out_org56;
   assign  _add_all_x_data_in_org57 = data_out_org57;
   assign  _add_all_x_data_in_org58 = data_out_org58;
   assign  _add_all_x_data_in_org59 = data_out_org59;
   assign  _add_all_x_data_in_org60 = data_out_org60;
   assign  _add_all_x_data_in_org61 = data_out_org61;
   assign  _add_all_x_data_in_org62 = data_out_org62;
   assign  _add_all_x_data_in_org65 = data_out_org65;
   assign  _add_all_x_data_in_org66 = data_out_org66;
   assign  _add_all_x_data_in_org67 = data_out_org67;
   assign  _add_all_x_data_in_org68 = data_out_org68;
   assign  _add_all_x_data_in_org69 = data_out_org69;
   assign  _add_all_x_data_in_org70 = data_out_org70;
   assign  _add_all_x_data_in_org71 = data_out_org71;
   assign  _add_all_x_data_in_org72 = data_out_org72;
   assign  _add_all_x_data_in_org73 = data_out_org73;
   assign  _add_all_x_data_in_org74 = data_out_org74;
   assign  _add_all_x_data_in_org75 = data_out_org75;
   assign  _add_all_x_data_in_org76 = data_out_org76;
   assign  _add_all_x_data_in_org77 = data_out_org77;
   assign  _add_all_x_data_in_org78 = data_out_org78;
   assign  _add_all_x_data_in_org79 = data_out_org79;
   assign  _add_all_x_data_in_org80 = data_out_org80;
   assign  _add_all_x_data_in_org81 = data_out_org81;
   assign  _add_all_x_data_in_org82 = data_out_org82;
   assign  _add_all_x_data_in_org83 = data_out_org83;
   assign  _add_all_x_data_in_org84 = data_out_org84;
   assign  _add_all_x_data_in_org85 = data_out_org85;
   assign  _add_all_x_data_in_org86 = data_out_org86;
   assign  _add_all_x_data_in_org87 = data_out_org87;
   assign  _add_all_x_data_in_org88 = data_out_org88;
   assign  _add_all_x_data_in_org89 = data_out_org89;
   assign  _add_all_x_data_in_org90 = data_out_org90;
   assign  _add_all_x_data_in_org91 = data_out_org91;
   assign  _add_all_x_data_in_org92 = data_out_org92;
   assign  _add_all_x_data_in_org93 = data_out_org93;
   assign  _add_all_x_data_in_org94 = data_out_org94;
   assign  _add_all_x_data_in_org97 = data_out_org97;
   assign  _add_all_x_data_in_org98 = data_out_org98;
   assign  _add_all_x_data_in_org99 = data_out_org99;
   assign  _add_all_x_data_in_org100 = data_out_org100;
   assign  _add_all_x_data_in_org101 = data_out_org101;
   assign  _add_all_x_data_in_org102 = data_out_org102;
   assign  _add_all_x_data_in_org103 = data_out_org103;
   assign  _add_all_x_data_in_org104 = data_out_org104;
   assign  _add_all_x_data_in_org105 = data_out_org105;
   assign  _add_all_x_data_in_org106 = data_out_org106;
   assign  _add_all_x_data_in_org107 = data_out_org107;
   assign  _add_all_x_data_in_org108 = data_out_org108;
   assign  _add_all_x_data_in_org109 = data_out_org109;
   assign  _add_all_x_data_in_org110 = data_out_org110;
   assign  _add_all_x_data_in_org111 = data_out_org111;
   assign  _add_all_x_data_in_org112 = data_out_org112;
   assign  _add_all_x_data_in_org113 = data_out_org113;
   assign  _add_all_x_data_in_org114 = data_out_org114;
   assign  _add_all_x_data_in_org115 = data_out_org115;
   assign  _add_all_x_data_in_org116 = data_out_org116;
   assign  _add_all_x_data_in_org117 = data_out_org117;
   assign  _add_all_x_data_in_org118 = data_out_org118;
   assign  _add_all_x_data_in_org119 = data_out_org119;
   assign  _add_all_x_data_in_org120 = data_out_org120;
   assign  _add_all_x_data_in_org121 = data_out_org121;
   assign  _add_all_x_data_in_org122 = data_out_org122;
   assign  _add_all_x_data_in_org123 = data_out_org123;
   assign  _add_all_x_data_in_org124 = data_out_org124;
   assign  _add_all_x_data_in_org125 = data_out_org125;
   assign  _add_all_x_data_in_org126 = data_out_org126;
   assign  _add_all_x_data_in_org129 = data_out_org129;
   assign  _add_all_x_data_in_org130 = data_out_org130;
   assign  _add_all_x_data_in_org131 = data_out_org131;
   assign  _add_all_x_data_in_org132 = data_out_org132;
   assign  _add_all_x_data_in_org133 = data_out_org133;
   assign  _add_all_x_data_in_org134 = data_out_org134;
   assign  _add_all_x_data_in_org135 = data_out_org135;
   assign  _add_all_x_data_in_org136 = data_out_org136;
   assign  _add_all_x_data_in_org137 = data_out_org137;
   assign  _add_all_x_data_in_org138 = data_out_org138;
   assign  _add_all_x_data_in_org139 = data_out_org139;
   assign  _add_all_x_data_in_org140 = data_out_org140;
   assign  _add_all_x_data_in_org141 = data_out_org141;
   assign  _add_all_x_data_in_org142 = data_out_org142;
   assign  _add_all_x_data_in_org143 = data_out_org143;
   assign  _add_all_x_data_in_org144 = data_out_org144;
   assign  _add_all_x_data_in_org145 = data_out_org145;
   assign  _add_all_x_data_in_org146 = data_out_org146;
   assign  _add_all_x_data_in_org147 = data_out_org147;
   assign  _add_all_x_data_in_org148 = data_out_org148;
   assign  _add_all_x_data_in_org149 = data_out_org149;
   assign  _add_all_x_data_in_org150 = data_out_org150;
   assign  _add_all_x_data_in_org151 = data_out_org151;
   assign  _add_all_x_data_in_org152 = data_out_org152;
   assign  _add_all_x_data_in_org153 = data_out_org153;
   assign  _add_all_x_data_in_org154 = data_out_org154;
   assign  _add_all_x_data_in_org155 = data_out_org155;
   assign  _add_all_x_data_in_org156 = data_out_org156;
   assign  _add_all_x_data_in_org157 = data_out_org157;
   assign  _add_all_x_data_in_org158 = data_out_org158;
   assign  _add_all_x_data_in_org161 = data_out_org161;
   assign  _add_all_x_data_in_org162 = data_out_org162;
   assign  _add_all_x_data_in_org163 = data_out_org163;
   assign  _add_all_x_data_in_org164 = data_out_org164;
   assign  _add_all_x_data_in_org165 = data_out_org165;
   assign  _add_all_x_data_in_org166 = data_out_org166;
   assign  _add_all_x_data_in_org167 = data_out_org167;
   assign  _add_all_x_data_in_org168 = data_out_org168;
   assign  _add_all_x_data_in_org169 = data_out_org169;
   assign  _add_all_x_data_in_org170 = data_out_org170;
   assign  _add_all_x_data_in_org171 = data_out_org171;
   assign  _add_all_x_data_in_org172 = data_out_org172;
   assign  _add_all_x_data_in_org173 = data_out_org173;
   assign  _add_all_x_data_in_org174 = data_out_org174;
   assign  _add_all_x_data_in_org175 = data_out_org175;
   assign  _add_all_x_data_in_org176 = data_out_org176;
   assign  _add_all_x_data_in_org177 = data_out_org177;
   assign  _add_all_x_data_in_org178 = data_out_org178;
   assign  _add_all_x_data_in_org179 = data_out_org179;
   assign  _add_all_x_data_in_org180 = data_out_org180;
   assign  _add_all_x_data_in_org181 = data_out_org181;
   assign  _add_all_x_data_in_org182 = data_out_org182;
   assign  _add_all_x_data_in_org183 = data_out_org183;
   assign  _add_all_x_data_in_org184 = data_out_org184;
   assign  _add_all_x_data_in_org185 = data_out_org185;
   assign  _add_all_x_data_in_org186 = data_out_org186;
   assign  _add_all_x_data_in_org187 = data_out_org187;
   assign  _add_all_x_data_in_org188 = data_out_org188;
   assign  _add_all_x_data_in_org189 = data_out_org189;
   assign  _add_all_x_data_in_org190 = data_out_org190;
   assign  _add_all_x_data_in_org193 = data_out_org193;
   assign  _add_all_x_data_in_org194 = data_out_org194;
   assign  _add_all_x_data_in_org195 = data_out_org195;
   assign  _add_all_x_data_in_org196 = data_out_org196;
   assign  _add_all_x_data_in_org197 = data_out_org197;
   assign  _add_all_x_data_in_org198 = data_out_org198;
   assign  _add_all_x_data_in_org199 = data_out_org199;
   assign  _add_all_x_data_in_org200 = data_out_org200;
   assign  _add_all_x_data_in_org201 = data_out_org201;
   assign  _add_all_x_data_in_org202 = data_out_org202;
   assign  _add_all_x_data_in_org203 = data_out_org203;
   assign  _add_all_x_data_in_org204 = data_out_org204;
   assign  _add_all_x_data_in_org205 = data_out_org205;
   assign  _add_all_x_data_in_org206 = data_out_org206;
   assign  _add_all_x_data_in_org207 = data_out_org207;
   assign  _add_all_x_data_in_org208 = data_out_org208;
   assign  _add_all_x_data_in_org209 = data_out_org209;
   assign  _add_all_x_data_in_org210 = data_out_org210;
   assign  _add_all_x_data_in_org211 = data_out_org211;
   assign  _add_all_x_data_in_org212 = data_out_org212;
   assign  _add_all_x_data_in_org213 = data_out_org213;
   assign  _add_all_x_data_in_org214 = data_out_org214;
   assign  _add_all_x_data_in_org215 = data_out_org215;
   assign  _add_all_x_data_in_org216 = data_out_org216;
   assign  _add_all_x_data_in_org217 = data_out_org217;
   assign  _add_all_x_data_in_org218 = data_out_org218;
   assign  _add_all_x_data_in_org219 = data_out_org219;
   assign  _add_all_x_data_in_org220 = data_out_org220;
   assign  _add_all_x_data_in_org221 = data_out_org221;
   assign  _add_all_x_data_in_org222 = data_out_org222;
   assign  _add_all_x_data_in_org225 = data_out_org225;
   assign  _add_all_x_data_in_org226 = data_out_org226;
   assign  _add_all_x_data_in_org227 = data_out_org227;
   assign  _add_all_x_data_in_org228 = data_out_org228;
   assign  _add_all_x_data_in_org229 = data_out_org229;
   assign  _add_all_x_data_in_org230 = data_out_org230;
   assign  _add_all_x_data_in_org231 = data_out_org231;
   assign  _add_all_x_data_in_org232 = data_out_org232;
   assign  _add_all_x_data_in_org233 = data_out_org233;
   assign  _add_all_x_data_in_org234 = data_out_org234;
   assign  _add_all_x_data_in_org235 = data_out_org235;
   assign  _add_all_x_data_in_org236 = data_out_org236;
   assign  _add_all_x_data_in_org237 = data_out_org237;
   assign  _add_all_x_data_in_org238 = data_out_org238;
   assign  _add_all_x_data_in_org239 = data_out_org239;
   assign  _add_all_x_data_in_org240 = data_out_org240;
   assign  _add_all_x_data_in_org241 = data_out_org241;
   assign  _add_all_x_data_in_org242 = data_out_org242;
   assign  _add_all_x_data_in_org243 = data_out_org243;
   assign  _add_all_x_data_in_org244 = data_out_org244;
   assign  _add_all_x_data_in_org245 = data_out_org245;
   assign  _add_all_x_data_in_org246 = data_out_org246;
   assign  _add_all_x_data_in_org247 = data_out_org247;
   assign  _add_all_x_data_in_org248 = data_out_org248;
   assign  _add_all_x_data_in_org249 = data_out_org249;
   assign  _add_all_x_data_in_org250 = data_out_org250;
   assign  _add_all_x_data_in_org251 = data_out_org251;
   assign  _add_all_x_data_in_org252 = data_out_org252;
   assign  _add_all_x_data_in_org253 = data_out_org253;
   assign  _add_all_x_data_in_org254 = data_out_org254;
   assign  _add_all_x_data_in_org257 = data_out_org257;
   assign  _add_all_x_data_in_org258 = data_out_org258;
   assign  _add_all_x_data_in_org259 = data_out_org259;
   assign  _add_all_x_data_in_org260 = data_out_org260;
   assign  _add_all_x_data_in_org261 = data_out_org261;
   assign  _add_all_x_data_in_org262 = data_out_org262;
   assign  _add_all_x_data_in_org263 = data_out_org263;
   assign  _add_all_x_data_in_org264 = data_out_org264;
   assign  _add_all_x_data_in_org265 = data_out_org265;
   assign  _add_all_x_data_in_org266 = data_out_org266;
   assign  _add_all_x_data_in_org267 = data_out_org267;
   assign  _add_all_x_data_in_org268 = data_out_org268;
   assign  _add_all_x_data_in_org269 = data_out_org269;
   assign  _add_all_x_data_in_org270 = data_out_org270;
   assign  _add_all_x_data_in_org271 = data_out_org271;
   assign  _add_all_x_data_in_org272 = data_out_org272;
   assign  _add_all_x_data_in_org273 = data_out_org273;
   assign  _add_all_x_data_in_org274 = data_out_org274;
   assign  _add_all_x_data_in_org275 = data_out_org275;
   assign  _add_all_x_data_in_org276 = data_out_org276;
   assign  _add_all_x_data_in_org277 = data_out_org277;
   assign  _add_all_x_data_in_org278 = data_out_org278;
   assign  _add_all_x_data_in_org279 = data_out_org279;
   assign  _add_all_x_data_in_org280 = data_out_org280;
   assign  _add_all_x_data_in_org281 = data_out_org281;
   assign  _add_all_x_data_in_org282 = data_out_org282;
   assign  _add_all_x_data_in_org283 = data_out_org283;
   assign  _add_all_x_data_in_org284 = data_out_org284;
   assign  _add_all_x_data_in_org285 = data_out_org285;
   assign  _add_all_x_data_in_org286 = data_out_org286;
   assign  _add_all_x_data_in_org289 = data_out_org289;
   assign  _add_all_x_data_in_org290 = data_out_org290;
   assign  _add_all_x_data_in_org291 = data_out_org291;
   assign  _add_all_x_data_in_org292 = data_out_org292;
   assign  _add_all_x_data_in_org293 = data_out_org293;
   assign  _add_all_x_data_in_org294 = data_out_org294;
   assign  _add_all_x_data_in_org295 = data_out_org295;
   assign  _add_all_x_data_in_org296 = data_out_org296;
   assign  _add_all_x_data_in_org297 = data_out_org297;
   assign  _add_all_x_data_in_org298 = data_out_org298;
   assign  _add_all_x_data_in_org299 = data_out_org299;
   assign  _add_all_x_data_in_org300 = data_out_org300;
   assign  _add_all_x_data_in_org301 = data_out_org301;
   assign  _add_all_x_data_in_org302 = data_out_org302;
   assign  _add_all_x_data_in_org303 = data_out_org303;
   assign  _add_all_x_data_in_org304 = data_out_org304;
   assign  _add_all_x_data_in_org305 = data_out_org305;
   assign  _add_all_x_data_in_org306 = data_out_org306;
   assign  _add_all_x_data_in_org307 = data_out_org307;
   assign  _add_all_x_data_in_org308 = data_out_org308;
   assign  _add_all_x_data_in_org309 = data_out_org309;
   assign  _add_all_x_data_in_org310 = data_out_org310;
   assign  _add_all_x_data_in_org311 = data_out_org311;
   assign  _add_all_x_data_in_org312 = data_out_org312;
   assign  _add_all_x_data_in_org313 = data_out_org313;
   assign  _add_all_x_data_in_org314 = data_out_org314;
   assign  _add_all_x_data_in_org315 = data_out_org315;
   assign  _add_all_x_data_in_org316 = data_out_org316;
   assign  _add_all_x_data_in_org317 = data_out_org317;
   assign  _add_all_x_data_in_org318 = data_out_org318;
   assign  _add_all_x_data_in_org321 = data_out_org321;
   assign  _add_all_x_data_in_org322 = data_out_org322;
   assign  _add_all_x_data_in_org323 = data_out_org323;
   assign  _add_all_x_data_in_org324 = data_out_org324;
   assign  _add_all_x_data_in_org325 = data_out_org325;
   assign  _add_all_x_data_in_org326 = data_out_org326;
   assign  _add_all_x_data_in_org327 = data_out_org327;
   assign  _add_all_x_data_in_org328 = data_out_org328;
   assign  _add_all_x_data_in_org329 = data_out_org329;
   assign  _add_all_x_data_in_org330 = data_out_org330;
   assign  _add_all_x_data_in_org331 = data_out_org331;
   assign  _add_all_x_data_in_org332 = data_out_org332;
   assign  _add_all_x_data_in_org333 = data_out_org333;
   assign  _add_all_x_data_in_org334 = data_out_org334;
   assign  _add_all_x_data_in_org335 = data_out_org335;
   assign  _add_all_x_data_in_org336 = data_out_org336;
   assign  _add_all_x_data_in_org337 = data_out_org337;
   assign  _add_all_x_data_in_org338 = data_out_org338;
   assign  _add_all_x_data_in_org339 = data_out_org339;
   assign  _add_all_x_data_in_org340 = data_out_org340;
   assign  _add_all_x_data_in_org341 = data_out_org341;
   assign  _add_all_x_data_in_org342 = data_out_org342;
   assign  _add_all_x_data_in_org343 = data_out_org343;
   assign  _add_all_x_data_in_org344 = data_out_org344;
   assign  _add_all_x_data_in_org345 = data_out_org345;
   assign  _add_all_x_data_in_org346 = data_out_org346;
   assign  _add_all_x_data_in_org347 = data_out_org347;
   assign  _add_all_x_data_in_org348 = data_out_org348;
   assign  _add_all_x_data_in_org349 = data_out_org349;
   assign  _add_all_x_data_in_org350 = data_out_org350;
   assign  _add_all_x_data_in_org353 = data_out_org353;
   assign  _add_all_x_data_in_org354 = data_out_org354;
   assign  _add_all_x_data_in_org355 = data_out_org355;
   assign  _add_all_x_data_in_org356 = data_out_org356;
   assign  _add_all_x_data_in_org357 = data_out_org357;
   assign  _add_all_x_data_in_org358 = data_out_org358;
   assign  _add_all_x_data_in_org359 = data_out_org359;
   assign  _add_all_x_data_in_org360 = data_out_org360;
   assign  _add_all_x_data_in_org361 = data_out_org361;
   assign  _add_all_x_data_in_org362 = data_out_org362;
   assign  _add_all_x_data_in_org363 = data_out_org363;
   assign  _add_all_x_data_in_org364 = data_out_org364;
   assign  _add_all_x_data_in_org365 = data_out_org365;
   assign  _add_all_x_data_in_org366 = data_out_org366;
   assign  _add_all_x_data_in_org367 = data_out_org367;
   assign  _add_all_x_data_in_org368 = data_out_org368;
   assign  _add_all_x_data_in_org369 = data_out_org369;
   assign  _add_all_x_data_in_org370 = data_out_org370;
   assign  _add_all_x_data_in_org371 = data_out_org371;
   assign  _add_all_x_data_in_org372 = data_out_org372;
   assign  _add_all_x_data_in_org373 = data_out_org373;
   assign  _add_all_x_data_in_org374 = data_out_org374;
   assign  _add_all_x_data_in_org375 = data_out_org375;
   assign  _add_all_x_data_in_org376 = data_out_org376;
   assign  _add_all_x_data_in_org377 = data_out_org377;
   assign  _add_all_x_data_in_org378 = data_out_org378;
   assign  _add_all_x_data_in_org379 = data_out_org379;
   assign  _add_all_x_data_in_org380 = data_out_org380;
   assign  _add_all_x_data_in_org381 = data_out_org381;
   assign  _add_all_x_data_in_org382 = data_out_org382;
   assign  _add_all_x_data_in_org385 = data_out_org385;
   assign  _add_all_x_data_in_org386 = data_out_org386;
   assign  _add_all_x_data_in_org387 = data_out_org387;
   assign  _add_all_x_data_in_org388 = data_out_org388;
   assign  _add_all_x_data_in_org389 = data_out_org389;
   assign  _add_all_x_data_in_org390 = data_out_org390;
   assign  _add_all_x_data_in_org391 = data_out_org391;
   assign  _add_all_x_data_in_org392 = data_out_org392;
   assign  _add_all_x_data_in_org393 = data_out_org393;
   assign  _add_all_x_data_in_org394 = data_out_org394;
   assign  _add_all_x_data_in_org395 = data_out_org395;
   assign  _add_all_x_data_in_org396 = data_out_org396;
   assign  _add_all_x_data_in_org397 = data_out_org397;
   assign  _add_all_x_data_in_org398 = data_out_org398;
   assign  _add_all_x_data_in_org399 = data_out_org399;
   assign  _add_all_x_data_in_org400 = data_out_org400;
   assign  _add_all_x_data_in_org401 = data_out_org401;
   assign  _add_all_x_data_in_org402 = data_out_org402;
   assign  _add_all_x_data_in_org403 = data_out_org403;
   assign  _add_all_x_data_in_org404 = data_out_org404;
   assign  _add_all_x_data_in_org405 = data_out_org405;
   assign  _add_all_x_data_in_org406 = data_out_org406;
   assign  _add_all_x_data_in_org407 = data_out_org407;
   assign  _add_all_x_data_in_org408 = data_out_org408;
   assign  _add_all_x_data_in_org409 = data_out_org409;
   assign  _add_all_x_data_in_org410 = data_out_org410;
   assign  _add_all_x_data_in_org411 = data_out_org411;
   assign  _add_all_x_data_in_org412 = data_out_org412;
   assign  _add_all_x_data_in_org413 = data_out_org413;
   assign  _add_all_x_data_in_org414 = data_out_org414;
   assign  _add_all_x_data_in_org417 = data_out_org417;
   assign  _add_all_x_data_in_org418 = data_out_org418;
   assign  _add_all_x_data_in_org419 = data_out_org419;
   assign  _add_all_x_data_in_org420 = data_out_org420;
   assign  _add_all_x_data_in_org421 = data_out_org421;
   assign  _add_all_x_data_in_org422 = data_out_org422;
   assign  _add_all_x_data_in_org423 = data_out_org423;
   assign  _add_all_x_data_in_org424 = data_out_org424;
   assign  _add_all_x_data_in_org425 = data_out_org425;
   assign  _add_all_x_data_in_org426 = data_out_org426;
   assign  _add_all_x_data_in_org427 = data_out_org427;
   assign  _add_all_x_data_in_org428 = data_out_org428;
   assign  _add_all_x_data_in_org429 = data_out_org429;
   assign  _add_all_x_data_in_org430 = data_out_org430;
   assign  _add_all_x_data_in_org431 = data_out_org431;
   assign  _add_all_x_data_in_org432 = data_out_org432;
   assign  _add_all_x_data_in_org433 = data_out_org433;
   assign  _add_all_x_data_in_org434 = data_out_org434;
   assign  _add_all_x_data_in_org435 = data_out_org435;
   assign  _add_all_x_data_in_org436 = data_out_org436;
   assign  _add_all_x_data_in_org437 = data_out_org437;
   assign  _add_all_x_data_in_org438 = data_out_org438;
   assign  _add_all_x_data_in_org439 = data_out_org439;
   assign  _add_all_x_data_in_org440 = data_out_org440;
   assign  _add_all_x_data_in_org441 = data_out_org441;
   assign  _add_all_x_data_in_org442 = data_out_org442;
   assign  _add_all_x_data_in_org443 = data_out_org443;
   assign  _add_all_x_data_in_org444 = data_out_org444;
   assign  _add_all_x_data_in_org445 = data_out_org445;
   assign  _add_all_x_data_in_org446 = data_out_org446;
   assign  _add_all_x_data_in_org449 = data_out_org449;
   assign  _add_all_x_data_in_org450 = data_out_org450;
   assign  _add_all_x_data_in_org451 = data_out_org451;
   assign  _add_all_x_data_in_org452 = data_out_org452;
   assign  _add_all_x_data_in_org453 = data_out_org453;
   assign  _add_all_x_data_in_org454 = data_out_org454;
   assign  _add_all_x_data_in_org455 = data_out_org455;
   assign  _add_all_x_data_in_org456 = data_out_org456;
   assign  _add_all_x_data_in_org457 = data_out_org457;
   assign  _add_all_x_data_in_org458 = data_out_org458;
   assign  _add_all_x_data_in_org459 = data_out_org459;
   assign  _add_all_x_data_in_org460 = data_out_org460;
   assign  _add_all_x_data_in_org461 = data_out_org461;
   assign  _add_all_x_data_in_org462 = data_out_org462;
   assign  _add_all_x_data_in_org463 = data_out_org463;
   assign  _add_all_x_data_in_org464 = data_out_org464;
   assign  _add_all_x_data_in_org465 = data_out_org465;
   assign  _add_all_x_data_in_org466 = data_out_org466;
   assign  _add_all_x_data_in_org467 = data_out_org467;
   assign  _add_all_x_data_in_org468 = data_out_org468;
   assign  _add_all_x_data_in_org469 = data_out_org469;
   assign  _add_all_x_data_in_org470 = data_out_org470;
   assign  _add_all_x_data_in_org471 = data_out_org471;
   assign  _add_all_x_data_in_org472 = data_out_org472;
   assign  _add_all_x_data_in_org473 = data_out_org473;
   assign  _add_all_x_data_in_org474 = data_out_org474;
   assign  _add_all_x_data_in_org475 = data_out_org475;
   assign  _add_all_x_data_in_org476 = data_out_org476;
   assign  _add_all_x_data_in_org477 = data_out_org477;
   assign  _add_all_x_data_in_org478 = data_out_org478;
   assign  _add_all_x_sg_in33 = sg33;
   assign  _add_all_x_sg_in34 = sg34;
   assign  _add_all_x_sg_in35 = sg35;
   assign  _add_all_x_sg_in36 = sg36;
   assign  _add_all_x_sg_in37 = sg37;
   assign  _add_all_x_sg_in38 = sg38;
   assign  _add_all_x_sg_in39 = sg39;
   assign  _add_all_x_sg_in40 = sg40;
   assign  _add_all_x_sg_in41 = sg41;
   assign  _add_all_x_sg_in42 = sg42;
   assign  _add_all_x_sg_in43 = sg43;
   assign  _add_all_x_sg_in44 = sg44;
   assign  _add_all_x_sg_in45 = sg45;
   assign  _add_all_x_sg_in46 = sg46;
   assign  _add_all_x_sg_in47 = sg47;
   assign  _add_all_x_sg_in48 = sg48;
   assign  _add_all_x_sg_in49 = sg49;
   assign  _add_all_x_sg_in50 = sg50;
   assign  _add_all_x_sg_in51 = sg51;
   assign  _add_all_x_sg_in52 = sg52;
   assign  _add_all_x_sg_in53 = sg53;
   assign  _add_all_x_sg_in54 = sg54;
   assign  _add_all_x_sg_in55 = sg55;
   assign  _add_all_x_sg_in56 = sg56;
   assign  _add_all_x_sg_in57 = sg57;
   assign  _add_all_x_sg_in58 = sg58;
   assign  _add_all_x_sg_in59 = sg59;
   assign  _add_all_x_sg_in60 = sg60;
   assign  _add_all_x_sg_in61 = sg61;
   assign  _add_all_x_sg_in62 = sg62;
   assign  _add_all_x_sg_in65 = sg65;
   assign  _add_all_x_sg_in66 = sg66;
   assign  _add_all_x_sg_in67 = sg67;
   assign  _add_all_x_sg_in68 = sg68;
   assign  _add_all_x_sg_in69 = sg69;
   assign  _add_all_x_sg_in70 = sg70;
   assign  _add_all_x_sg_in71 = sg71;
   assign  _add_all_x_sg_in72 = sg72;
   assign  _add_all_x_sg_in73 = sg73;
   assign  _add_all_x_sg_in74 = sg74;
   assign  _add_all_x_sg_in75 = sg75;
   assign  _add_all_x_sg_in76 = sg76;
   assign  _add_all_x_sg_in77 = sg77;
   assign  _add_all_x_sg_in78 = sg78;
   assign  _add_all_x_sg_in79 = sg79;
   assign  _add_all_x_sg_in80 = sg80;
   assign  _add_all_x_sg_in81 = sg81;
   assign  _add_all_x_sg_in82 = sg82;
   assign  _add_all_x_sg_in83 = sg83;
   assign  _add_all_x_sg_in84 = sg84;
   assign  _add_all_x_sg_in85 = sg85;
   assign  _add_all_x_sg_in86 = sg86;
   assign  _add_all_x_sg_in87 = sg87;
   assign  _add_all_x_sg_in88 = sg88;
   assign  _add_all_x_sg_in89 = sg89;
   assign  _add_all_x_sg_in90 = sg90;
   assign  _add_all_x_sg_in91 = sg91;
   assign  _add_all_x_sg_in92 = sg92;
   assign  _add_all_x_sg_in93 = sg93;
   assign  _add_all_x_sg_in94 = sg94;
   assign  _add_all_x_sg_in97 = sg97;
   assign  _add_all_x_sg_in98 = sg98;
   assign  _add_all_x_sg_in99 = sg99;
   assign  _add_all_x_sg_in100 = sg100;
   assign  _add_all_x_sg_in101 = sg101;
   assign  _add_all_x_sg_in102 = sg102;
   assign  _add_all_x_sg_in103 = sg103;
   assign  _add_all_x_sg_in104 = sg104;
   assign  _add_all_x_sg_in105 = sg105;
   assign  _add_all_x_sg_in106 = sg106;
   assign  _add_all_x_sg_in107 = sg107;
   assign  _add_all_x_sg_in108 = sg108;
   assign  _add_all_x_sg_in109 = sg109;
   assign  _add_all_x_sg_in110 = sg110;
   assign  _add_all_x_sg_in111 = sg111;
   assign  _add_all_x_sg_in112 = sg112;
   assign  _add_all_x_sg_in113 = sg113;
   assign  _add_all_x_sg_in114 = sg114;
   assign  _add_all_x_sg_in115 = sg115;
   assign  _add_all_x_sg_in116 = sg116;
   assign  _add_all_x_sg_in117 = sg117;
   assign  _add_all_x_sg_in118 = sg118;
   assign  _add_all_x_sg_in119 = sg119;
   assign  _add_all_x_sg_in120 = sg120;
   assign  _add_all_x_sg_in121 = sg121;
   assign  _add_all_x_sg_in122 = sg122;
   assign  _add_all_x_sg_in123 = sg123;
   assign  _add_all_x_sg_in124 = sg124;
   assign  _add_all_x_sg_in125 = sg125;
   assign  _add_all_x_sg_in126 = sg126;
   assign  _add_all_x_sg_in129 = sg129;
   assign  _add_all_x_sg_in130 = sg130;
   assign  _add_all_x_sg_in131 = sg131;
   assign  _add_all_x_sg_in132 = sg132;
   assign  _add_all_x_sg_in133 = sg133;
   assign  _add_all_x_sg_in134 = sg134;
   assign  _add_all_x_sg_in135 = sg135;
   assign  _add_all_x_sg_in136 = sg136;
   assign  _add_all_x_sg_in137 = sg137;
   assign  _add_all_x_sg_in138 = sg138;
   assign  _add_all_x_sg_in139 = sg139;
   assign  _add_all_x_sg_in140 = sg140;
   assign  _add_all_x_sg_in141 = sg141;
   assign  _add_all_x_sg_in142 = sg142;
   assign  _add_all_x_sg_in143 = sg143;
   assign  _add_all_x_sg_in144 = sg144;
   assign  _add_all_x_sg_in145 = sg145;
   assign  _add_all_x_sg_in146 = sg146;
   assign  _add_all_x_sg_in147 = sg147;
   assign  _add_all_x_sg_in148 = sg148;
   assign  _add_all_x_sg_in149 = sg149;
   assign  _add_all_x_sg_in150 = sg150;
   assign  _add_all_x_sg_in151 = sg151;
   assign  _add_all_x_sg_in152 = sg152;
   assign  _add_all_x_sg_in153 = sg153;
   assign  _add_all_x_sg_in154 = sg154;
   assign  _add_all_x_sg_in155 = sg155;
   assign  _add_all_x_sg_in156 = sg156;
   assign  _add_all_x_sg_in157 = sg157;
   assign  _add_all_x_sg_in158 = sg158;
   assign  _add_all_x_sg_in161 = sg161;
   assign  _add_all_x_sg_in162 = sg162;
   assign  _add_all_x_sg_in163 = sg163;
   assign  _add_all_x_sg_in164 = sg164;
   assign  _add_all_x_sg_in165 = sg165;
   assign  _add_all_x_sg_in166 = sg166;
   assign  _add_all_x_sg_in167 = sg167;
   assign  _add_all_x_sg_in168 = sg168;
   assign  _add_all_x_sg_in169 = sg169;
   assign  _add_all_x_sg_in170 = sg170;
   assign  _add_all_x_sg_in171 = sg171;
   assign  _add_all_x_sg_in172 = sg172;
   assign  _add_all_x_sg_in173 = sg173;
   assign  _add_all_x_sg_in174 = sg174;
   assign  _add_all_x_sg_in175 = sg175;
   assign  _add_all_x_sg_in176 = sg176;
   assign  _add_all_x_sg_in177 = sg177;
   assign  _add_all_x_sg_in178 = sg178;
   assign  _add_all_x_sg_in179 = sg179;
   assign  _add_all_x_sg_in180 = sg180;
   assign  _add_all_x_sg_in181 = sg181;
   assign  _add_all_x_sg_in182 = sg182;
   assign  _add_all_x_sg_in183 = sg183;
   assign  _add_all_x_sg_in184 = sg184;
   assign  _add_all_x_sg_in185 = sg185;
   assign  _add_all_x_sg_in186 = sg186;
   assign  _add_all_x_sg_in187 = sg187;
   assign  _add_all_x_sg_in188 = sg188;
   assign  _add_all_x_sg_in189 = sg189;
   assign  _add_all_x_sg_in190 = sg190;
   assign  _add_all_x_sg_in193 = sg193;
   assign  _add_all_x_sg_in194 = sg194;
   assign  _add_all_x_sg_in195 = sg195;
   assign  _add_all_x_sg_in196 = sg196;
   assign  _add_all_x_sg_in197 = sg197;
   assign  _add_all_x_sg_in198 = sg198;
   assign  _add_all_x_sg_in199 = sg199;
   assign  _add_all_x_sg_in200 = sg200;
   assign  _add_all_x_sg_in201 = sg201;
   assign  _add_all_x_sg_in202 = sg202;
   assign  _add_all_x_sg_in203 = sg203;
   assign  _add_all_x_sg_in204 = sg204;
   assign  _add_all_x_sg_in205 = sg205;
   assign  _add_all_x_sg_in206 = sg206;
   assign  _add_all_x_sg_in207 = sg207;
   assign  _add_all_x_sg_in208 = sg208;
   assign  _add_all_x_sg_in209 = sg209;
   assign  _add_all_x_sg_in210 = sg210;
   assign  _add_all_x_sg_in211 = sg211;
   assign  _add_all_x_sg_in212 = sg212;
   assign  _add_all_x_sg_in213 = sg213;
   assign  _add_all_x_sg_in214 = sg214;
   assign  _add_all_x_sg_in215 = sg215;
   assign  _add_all_x_sg_in216 = sg216;
   assign  _add_all_x_sg_in217 = sg217;
   assign  _add_all_x_sg_in218 = sg218;
   assign  _add_all_x_sg_in219 = sg219;
   assign  _add_all_x_sg_in220 = sg220;
   assign  _add_all_x_sg_in221 = sg221;
   assign  _add_all_x_sg_in222 = sg222;
   assign  _add_all_x_sg_in225 = sg225;
   assign  _add_all_x_sg_in226 = sg226;
   assign  _add_all_x_sg_in227 = sg227;
   assign  _add_all_x_sg_in228 = sg228;
   assign  _add_all_x_sg_in229 = sg229;
   assign  _add_all_x_sg_in230 = sg230;
   assign  _add_all_x_sg_in231 = sg231;
   assign  _add_all_x_sg_in232 = sg232;
   assign  _add_all_x_sg_in233 = sg233;
   assign  _add_all_x_sg_in234 = sg234;
   assign  _add_all_x_sg_in235 = sg235;
   assign  _add_all_x_sg_in236 = sg236;
   assign  _add_all_x_sg_in237 = sg237;
   assign  _add_all_x_sg_in238 = sg238;
   assign  _add_all_x_sg_in239 = sg239;
   assign  _add_all_x_sg_in240 = sg240;
   assign  _add_all_x_sg_in241 = sg241;
   assign  _add_all_x_sg_in242 = sg242;
   assign  _add_all_x_sg_in243 = sg243;
   assign  _add_all_x_sg_in244 = sg244;
   assign  _add_all_x_sg_in245 = sg245;
   assign  _add_all_x_sg_in246 = sg246;
   assign  _add_all_x_sg_in247 = sg247;
   assign  _add_all_x_sg_in248 = sg248;
   assign  _add_all_x_sg_in249 = sg249;
   assign  _add_all_x_sg_in250 = sg250;
   assign  _add_all_x_sg_in251 = sg251;
   assign  _add_all_x_sg_in252 = sg252;
   assign  _add_all_x_sg_in253 = sg253;
   assign  _add_all_x_sg_in254 = sg254;
   assign  _add_all_x_sg_in257 = sg257;
   assign  _add_all_x_sg_in258 = sg258;
   assign  _add_all_x_sg_in259 = sg259;
   assign  _add_all_x_sg_in260 = sg260;
   assign  _add_all_x_sg_in261 = sg261;
   assign  _add_all_x_sg_in262 = sg262;
   assign  _add_all_x_sg_in263 = sg263;
   assign  _add_all_x_sg_in264 = sg264;
   assign  _add_all_x_sg_in265 = sg265;
   assign  _add_all_x_sg_in266 = sg266;
   assign  _add_all_x_sg_in267 = sg267;
   assign  _add_all_x_sg_in268 = sg268;
   assign  _add_all_x_sg_in269 = sg269;
   assign  _add_all_x_sg_in270 = sg270;
   assign  _add_all_x_sg_in271 = sg271;
   assign  _add_all_x_sg_in272 = sg272;
   assign  _add_all_x_sg_in273 = sg273;
   assign  _add_all_x_sg_in274 = sg274;
   assign  _add_all_x_sg_in275 = sg275;
   assign  _add_all_x_sg_in276 = sg276;
   assign  _add_all_x_sg_in277 = sg277;
   assign  _add_all_x_sg_in278 = sg278;
   assign  _add_all_x_sg_in279 = sg279;
   assign  _add_all_x_sg_in280 = sg280;
   assign  _add_all_x_sg_in281 = sg281;
   assign  _add_all_x_sg_in282 = sg282;
   assign  _add_all_x_sg_in283 = sg283;
   assign  _add_all_x_sg_in284 = sg284;
   assign  _add_all_x_sg_in285 = sg285;
   assign  _add_all_x_sg_in286 = sg286;
   assign  _add_all_x_sg_in289 = sg289;
   assign  _add_all_x_sg_in290 = sg290;
   assign  _add_all_x_sg_in291 = sg291;
   assign  _add_all_x_sg_in292 = sg292;
   assign  _add_all_x_sg_in293 = sg293;
   assign  _add_all_x_sg_in294 = sg294;
   assign  _add_all_x_sg_in295 = sg295;
   assign  _add_all_x_sg_in296 = sg296;
   assign  _add_all_x_sg_in297 = sg297;
   assign  _add_all_x_sg_in298 = sg298;
   assign  _add_all_x_sg_in299 = sg299;
   assign  _add_all_x_sg_in300 = sg300;
   assign  _add_all_x_sg_in301 = sg301;
   assign  _add_all_x_sg_in302 = sg302;
   assign  _add_all_x_sg_in303 = sg303;
   assign  _add_all_x_sg_in304 = sg304;
   assign  _add_all_x_sg_in305 = sg305;
   assign  _add_all_x_sg_in306 = sg306;
   assign  _add_all_x_sg_in307 = sg307;
   assign  _add_all_x_sg_in308 = sg308;
   assign  _add_all_x_sg_in309 = sg309;
   assign  _add_all_x_sg_in310 = sg310;
   assign  _add_all_x_sg_in311 = sg311;
   assign  _add_all_x_sg_in312 = sg312;
   assign  _add_all_x_sg_in313 = sg313;
   assign  _add_all_x_sg_in314 = sg314;
   assign  _add_all_x_sg_in315 = sg315;
   assign  _add_all_x_sg_in316 = sg316;
   assign  _add_all_x_sg_in317 = sg317;
   assign  _add_all_x_sg_in318 = sg318;
   assign  _add_all_x_sg_in321 = sg321;
   assign  _add_all_x_sg_in322 = sg322;
   assign  _add_all_x_sg_in323 = sg323;
   assign  _add_all_x_sg_in324 = sg324;
   assign  _add_all_x_sg_in325 = sg325;
   assign  _add_all_x_sg_in326 = sg326;
   assign  _add_all_x_sg_in327 = sg327;
   assign  _add_all_x_sg_in328 = sg328;
   assign  _add_all_x_sg_in329 = sg329;
   assign  _add_all_x_sg_in330 = sg330;
   assign  _add_all_x_sg_in331 = sg331;
   assign  _add_all_x_sg_in332 = sg332;
   assign  _add_all_x_sg_in333 = sg333;
   assign  _add_all_x_sg_in334 = sg334;
   assign  _add_all_x_sg_in335 = sg335;
   assign  _add_all_x_sg_in336 = sg336;
   assign  _add_all_x_sg_in337 = sg337;
   assign  _add_all_x_sg_in338 = sg338;
   assign  _add_all_x_sg_in339 = sg339;
   assign  _add_all_x_sg_in340 = sg340;
   assign  _add_all_x_sg_in341 = sg341;
   assign  _add_all_x_sg_in342 = sg342;
   assign  _add_all_x_sg_in343 = sg343;
   assign  _add_all_x_sg_in344 = sg344;
   assign  _add_all_x_sg_in345 = sg345;
   assign  _add_all_x_sg_in346 = sg346;
   assign  _add_all_x_sg_in347 = sg347;
   assign  _add_all_x_sg_in348 = sg348;
   assign  _add_all_x_sg_in349 = sg349;
   assign  _add_all_x_sg_in350 = sg350;
   assign  _add_all_x_sg_in353 = sg353;
   assign  _add_all_x_sg_in354 = sg354;
   assign  _add_all_x_sg_in355 = sg355;
   assign  _add_all_x_sg_in356 = sg356;
   assign  _add_all_x_sg_in357 = sg357;
   assign  _add_all_x_sg_in358 = sg358;
   assign  _add_all_x_sg_in359 = sg359;
   assign  _add_all_x_sg_in360 = sg360;
   assign  _add_all_x_sg_in361 = sg361;
   assign  _add_all_x_sg_in362 = sg362;
   assign  _add_all_x_sg_in363 = sg363;
   assign  _add_all_x_sg_in364 = sg364;
   assign  _add_all_x_sg_in365 = sg365;
   assign  _add_all_x_sg_in366 = sg366;
   assign  _add_all_x_sg_in367 = sg367;
   assign  _add_all_x_sg_in368 = sg368;
   assign  _add_all_x_sg_in369 = sg369;
   assign  _add_all_x_sg_in370 = sg370;
   assign  _add_all_x_sg_in371 = sg371;
   assign  _add_all_x_sg_in372 = sg372;
   assign  _add_all_x_sg_in373 = sg373;
   assign  _add_all_x_sg_in374 = sg374;
   assign  _add_all_x_sg_in375 = sg375;
   assign  _add_all_x_sg_in376 = sg376;
   assign  _add_all_x_sg_in377 = sg377;
   assign  _add_all_x_sg_in378 = sg378;
   assign  _add_all_x_sg_in379 = sg379;
   assign  _add_all_x_sg_in380 = sg380;
   assign  _add_all_x_sg_in381 = sg381;
   assign  _add_all_x_sg_in382 = sg382;
   assign  _add_all_x_sg_in385 = sg385;
   assign  _add_all_x_sg_in386 = sg386;
   assign  _add_all_x_sg_in387 = sg387;
   assign  _add_all_x_sg_in388 = sg388;
   assign  _add_all_x_sg_in389 = sg389;
   assign  _add_all_x_sg_in390 = sg390;
   assign  _add_all_x_sg_in391 = sg391;
   assign  _add_all_x_sg_in392 = sg392;
   assign  _add_all_x_sg_in393 = sg393;
   assign  _add_all_x_sg_in394 = sg394;
   assign  _add_all_x_sg_in395 = sg395;
   assign  _add_all_x_sg_in396 = sg396;
   assign  _add_all_x_sg_in397 = sg397;
   assign  _add_all_x_sg_in398 = sg398;
   assign  _add_all_x_sg_in399 = sg399;
   assign  _add_all_x_sg_in400 = sg400;
   assign  _add_all_x_sg_in401 = sg401;
   assign  _add_all_x_sg_in402 = sg402;
   assign  _add_all_x_sg_in403 = sg403;
   assign  _add_all_x_sg_in404 = sg404;
   assign  _add_all_x_sg_in405 = sg405;
   assign  _add_all_x_sg_in406 = sg406;
   assign  _add_all_x_sg_in407 = sg407;
   assign  _add_all_x_sg_in408 = sg408;
   assign  _add_all_x_sg_in409 = sg409;
   assign  _add_all_x_sg_in410 = sg410;
   assign  _add_all_x_sg_in411 = sg411;
   assign  _add_all_x_sg_in412 = sg412;
   assign  _add_all_x_sg_in413 = sg413;
   assign  _add_all_x_sg_in414 = sg414;
   assign  _add_all_x_sg_in417 = sg417;
   assign  _add_all_x_sg_in418 = sg418;
   assign  _add_all_x_sg_in419 = sg419;
   assign  _add_all_x_sg_in420 = sg420;
   assign  _add_all_x_sg_in421 = sg421;
   assign  _add_all_x_sg_in422 = sg422;
   assign  _add_all_x_sg_in423 = sg423;
   assign  _add_all_x_sg_in424 = sg424;
   assign  _add_all_x_sg_in425 = sg425;
   assign  _add_all_x_sg_in426 = sg426;
   assign  _add_all_x_sg_in427 = sg427;
   assign  _add_all_x_sg_in428 = sg428;
   assign  _add_all_x_sg_in429 = sg429;
   assign  _add_all_x_sg_in430 = sg430;
   assign  _add_all_x_sg_in431 = sg431;
   assign  _add_all_x_sg_in432 = sg432;
   assign  _add_all_x_sg_in433 = sg433;
   assign  _add_all_x_sg_in434 = sg434;
   assign  _add_all_x_sg_in435 = sg435;
   assign  _add_all_x_sg_in436 = sg436;
   assign  _add_all_x_sg_in437 = sg437;
   assign  _add_all_x_sg_in438 = sg438;
   assign  _add_all_x_sg_in439 = sg439;
   assign  _add_all_x_sg_in440 = sg440;
   assign  _add_all_x_sg_in441 = sg441;
   assign  _add_all_x_sg_in442 = sg442;
   assign  _add_all_x_sg_in443 = sg443;
   assign  _add_all_x_sg_in444 = sg444;
   assign  _add_all_x_sg_in445 = sg445;
   assign  _add_all_x_sg_in446 = sg446;
   assign  _add_all_x_sg_in449 = sg449;
   assign  _add_all_x_sg_in450 = sg450;
   assign  _add_all_x_sg_in451 = sg451;
   assign  _add_all_x_sg_in452 = sg452;
   assign  _add_all_x_sg_in453 = sg453;
   assign  _add_all_x_sg_in454 = sg454;
   assign  _add_all_x_sg_in455 = sg455;
   assign  _add_all_x_sg_in456 = sg456;
   assign  _add_all_x_sg_in457 = sg457;
   assign  _add_all_x_sg_in458 = sg458;
   assign  _add_all_x_sg_in459 = sg459;
   assign  _add_all_x_sg_in460 = sg460;
   assign  _add_all_x_sg_in461 = sg461;
   assign  _add_all_x_sg_in462 = sg462;
   assign  _add_all_x_sg_in463 = sg463;
   assign  _add_all_x_sg_in464 = sg464;
   assign  _add_all_x_sg_in465 = sg465;
   assign  _add_all_x_sg_in466 = sg466;
   assign  _add_all_x_sg_in467 = sg467;
   assign  _add_all_x_sg_in468 = sg468;
   assign  _add_all_x_sg_in469 = sg469;
   assign  _add_all_x_sg_in470 = sg470;
   assign  _add_all_x_sg_in471 = sg471;
   assign  _add_all_x_sg_in472 = sg472;
   assign  _add_all_x_sg_in473 = sg473;
   assign  _add_all_x_sg_in474 = sg474;
   assign  _add_all_x_sg_in475 = sg475;
   assign  _add_all_x_sg_in476 = sg476;
   assign  _add_all_x_sg_in477 = sg477;
   assign  _add_all_x_sg_in478 = sg478;
   assign  _add_all_x_in_do = kanwa_s;
   assign  _add_all_x_p_reset = p_reset;
   assign  _add_all_x_m_clock = m_clock;
   assign  _sub_x_data_in33 = ((_net_3181)?_add_all_x_data_out_index34:10'b0)|
    ((_net_2760)?_add_all_x_data_out_index33:10'b0);
   assign  _sub_x_data_in35 = ((_net_3180)?_add_all_x_data_out_index36:10'b0)|
    ((_net_2759)?_add_all_x_data_out_index35:10'b0);
   assign  _sub_x_data_in37 = ((_net_3179)?_add_all_x_data_out_index38:10'b0)|
    ((_net_2758)?_add_all_x_data_out_index37:10'b0);
   assign  _sub_x_data_in39 = ((_net_3178)?_add_all_x_data_out_index40:10'b0)|
    ((_net_2757)?_add_all_x_data_out_index39:10'b0);
   assign  _sub_x_data_in41 = ((_net_3177)?_add_all_x_data_out_index42:10'b0)|
    ((_net_2756)?_add_all_x_data_out_index41:10'b0);
   assign  _sub_x_data_in43 = ((_net_3176)?_add_all_x_data_out_index44:10'b0)|
    ((_net_2755)?_add_all_x_data_out_index43:10'b0);
   assign  _sub_x_data_in45 = ((_net_3175)?_add_all_x_data_out_index46:10'b0)|
    ((_net_2754)?_add_all_x_data_out_index45:10'b0);
   assign  _sub_x_data_in47 = ((_net_3174)?_add_all_x_data_out_index48:10'b0)|
    ((_net_2753)?_add_all_x_data_out_index47:10'b0);
   assign  _sub_x_data_in49 = ((_net_3173)?_add_all_x_data_out_index50:10'b0)|
    ((_net_2752)?_add_all_x_data_out_index49:10'b0);
   assign  _sub_x_data_in51 = ((_net_3172)?_add_all_x_data_out_index52:10'b0)|
    ((_net_2751)?_add_all_x_data_out_index51:10'b0);
   assign  _sub_x_data_in53 = ((_net_3171)?_add_all_x_data_out_index54:10'b0)|
    ((_net_2750)?_add_all_x_data_out_index53:10'b0);
   assign  _sub_x_data_in55 = ((_net_3170)?_add_all_x_data_out_index56:10'b0)|
    ((_net_2749)?_add_all_x_data_out_index55:10'b0);
   assign  _sub_x_data_in57 = ((_net_3169)?_add_all_x_data_out_index58:10'b0)|
    ((_net_2748)?_add_all_x_data_out_index57:10'b0);
   assign  _sub_x_data_in59 = ((_net_3168)?_add_all_x_data_out_index60:10'b0)|
    ((_net_2747)?_add_all_x_data_out_index59:10'b0);
   assign  _sub_x_data_in61 = ((_net_3167)?_add_all_x_data_out_index62:10'b0)|
    ((_net_2746)?_add_all_x_data_out_index61:10'b0);
   assign  _sub_x_data_in65 = ((_net_3166)?_add_all_x_data_out_index65:10'b0)|
    ((_net_2745)?_add_all_x_data_out_index66:10'b0);
   assign  _sub_x_data_in67 = ((_net_3165)?_add_all_x_data_out_index67:10'b0)|
    ((_net_2744)?_add_all_x_data_out_index68:10'b0);
   assign  _sub_x_data_in69 = ((_net_3164)?_add_all_x_data_out_index69:10'b0)|
    ((_net_2743)?_add_all_x_data_out_index70:10'b0);
   assign  _sub_x_data_in71 = ((_net_3163)?_add_all_x_data_out_index71:10'b0)|
    ((_net_2742)?_add_all_x_data_out_index72:10'b0);
   assign  _sub_x_data_in73 = ((_net_3162)?_add_all_x_data_out_index73:10'b0)|
    ((_net_2741)?_add_all_x_data_out_index74:10'b0);
   assign  _sub_x_data_in75 = ((_net_3161)?_add_all_x_data_out_index75:10'b0)|
    ((_net_2740)?_add_all_x_data_out_index76:10'b0);
   assign  _sub_x_data_in77 = ((_net_3160)?_add_all_x_data_out_index77:10'b0)|
    ((_net_2739)?_add_all_x_data_out_index78:10'b0);
   assign  _sub_x_data_in79 = ((_net_3159)?_add_all_x_data_out_index79:10'b0)|
    ((_net_2738)?_add_all_x_data_out_index80:10'b0);
   assign  _sub_x_data_in81 = ((_net_3158)?_add_all_x_data_out_index81:10'b0)|
    ((_net_2737)?_add_all_x_data_out_index82:10'b0);
   assign  _sub_x_data_in83 = ((_net_3157)?_add_all_x_data_out_index83:10'b0)|
    ((_net_2736)?_add_all_x_data_out_index84:10'b0);
   assign  _sub_x_data_in85 = ((_net_3156)?_add_all_x_data_out_index85:10'b0)|
    ((_net_2735)?_add_all_x_data_out_index86:10'b0);
   assign  _sub_x_data_in87 = ((_net_3155)?_add_all_x_data_out_index87:10'b0)|
    ((_net_2734)?_add_all_x_data_out_index88:10'b0);
   assign  _sub_x_data_in89 = ((_net_3154)?_add_all_x_data_out_index89:10'b0)|
    ((_net_2733)?_add_all_x_data_out_index90:10'b0);
   assign  _sub_x_data_in91 = ((_net_3153)?_add_all_x_data_out_index91:10'b0)|
    ((_net_2732)?_add_all_x_data_out_index92:10'b0);
   assign  _sub_x_data_in93 = ((_net_3152)?_add_all_x_data_out_index93:10'b0)|
    ((_net_2731)?_add_all_x_data_out_index94:10'b0);
   assign  _sub_x_data_in97 = ((_net_3151)?_add_all_x_data_out_index98:10'b0)|
    ((_net_2730)?_add_all_x_data_out_index97:10'b0);
   assign  _sub_x_data_in99 = ((_net_3150)?_add_all_x_data_out_index100:10'b0)|
    ((_net_2729)?_add_all_x_data_out_index99:10'b0);
   assign  _sub_x_data_in101 = ((_net_3149)?_add_all_x_data_out_index102:10'b0)|
    ((_net_2728)?_add_all_x_data_out_index101:10'b0);
   assign  _sub_x_data_in103 = ((_net_3148)?_add_all_x_data_out_index104:10'b0)|
    ((_net_2727)?_add_all_x_data_out_index103:10'b0);
   assign  _sub_x_data_in105 = ((_net_3147)?_add_all_x_data_out_index106:10'b0)|
    ((_net_2726)?_add_all_x_data_out_index105:10'b0);
   assign  _sub_x_data_in107 = ((_net_3146)?_add_all_x_data_out_index108:10'b0)|
    ((_net_2725)?_add_all_x_data_out_index107:10'b0);
   assign  _sub_x_data_in109 = ((_net_3145)?_add_all_x_data_out_index110:10'b0)|
    ((_net_2724)?_add_all_x_data_out_index109:10'b0);
   assign  _sub_x_data_in111 = ((_net_3144)?_add_all_x_data_out_index112:10'b0)|
    ((_net_2723)?_add_all_x_data_out_index111:10'b0);
   assign  _sub_x_data_in113 = ((_net_3143)?_add_all_x_data_out_index114:10'b0)|
    ((_net_2722)?_add_all_x_data_out_index113:10'b0);
   assign  _sub_x_data_in115 = ((_net_3142)?_add_all_x_data_out_index116:10'b0)|
    ((_net_2721)?_add_all_x_data_out_index115:10'b0);
   assign  _sub_x_data_in117 = ((_net_3141)?_add_all_x_data_out_index118:10'b0)|
    ((_net_2720)?_add_all_x_data_out_index117:10'b0);
   assign  _sub_x_data_in119 = ((_net_3140)?_add_all_x_data_out_index120:10'b0)|
    ((_net_2719)?_add_all_x_data_out_index119:10'b0);
   assign  _sub_x_data_in121 = ((_net_3139)?_add_all_x_data_out_index122:10'b0)|
    ((_net_2718)?_add_all_x_data_out_index121:10'b0);
   assign  _sub_x_data_in123 = ((_net_3138)?_add_all_x_data_out_index124:10'b0)|
    ((_net_2717)?_add_all_x_data_out_index123:10'b0);
   assign  _sub_x_data_in125 = ((_net_3137)?_add_all_x_data_out_index126:10'b0)|
    ((_net_2716)?_add_all_x_data_out_index125:10'b0);
   assign  _sub_x_data_in129 = ((_net_3136)?_add_all_x_data_out_index129:10'b0)|
    ((_net_2715)?_add_all_x_data_out_index130:10'b0);
   assign  _sub_x_data_in131 = ((_net_3135)?_add_all_x_data_out_index131:10'b0)|
    ((_net_2714)?_add_all_x_data_out_index132:10'b0);
   assign  _sub_x_data_in133 = ((_net_3134)?_add_all_x_data_out_index133:10'b0)|
    ((_net_2713)?_add_all_x_data_out_index134:10'b0);
   assign  _sub_x_data_in135 = ((_net_3133)?_add_all_x_data_out_index135:10'b0)|
    ((_net_2712)?_add_all_x_data_out_index136:10'b0);
   assign  _sub_x_data_in137 = ((_net_3132)?_add_all_x_data_out_index137:10'b0)|
    ((_net_2711)?_add_all_x_data_out_index138:10'b0);
   assign  _sub_x_data_in139 = ((_net_3131)?_add_all_x_data_out_index139:10'b0)|
    ((_net_2710)?_add_all_x_data_out_index140:10'b0);
   assign  _sub_x_data_in141 = ((_net_3130)?_add_all_x_data_out_index141:10'b0)|
    ((_net_2709)?_add_all_x_data_out_index142:10'b0);
   assign  _sub_x_data_in143 = ((_net_3129)?_add_all_x_data_out_index143:10'b0)|
    ((_net_2708)?_add_all_x_data_out_index144:10'b0);
   assign  _sub_x_data_in145 = ((_net_3128)?_add_all_x_data_out_index145:10'b0)|
    ((_net_2707)?_add_all_x_data_out_index146:10'b0);
   assign  _sub_x_data_in147 = ((_net_3127)?_add_all_x_data_out_index147:10'b0)|
    ((_net_2706)?_add_all_x_data_out_index148:10'b0);
   assign  _sub_x_data_in149 = ((_net_3126)?_add_all_x_data_out_index149:10'b0)|
    ((_net_2705)?_add_all_x_data_out_index150:10'b0);
   assign  _sub_x_data_in151 = ((_net_3125)?_add_all_x_data_out_index151:10'b0)|
    ((_net_2704)?_add_all_x_data_out_index152:10'b0);
   assign  _sub_x_data_in153 = ((_net_3124)?_add_all_x_data_out_index153:10'b0)|
    ((_net_2703)?_add_all_x_data_out_index154:10'b0);
   assign  _sub_x_data_in155 = ((_net_3123)?_add_all_x_data_out_index155:10'b0)|
    ((_net_2702)?_add_all_x_data_out_index156:10'b0);
   assign  _sub_x_data_in157 = ((_net_3122)?_add_all_x_data_out_index157:10'b0)|
    ((_net_2701)?_add_all_x_data_out_index158:10'b0);
   assign  _sub_x_data_in161 = ((_net_3121)?_add_all_x_data_out_index162:10'b0)|
    ((_net_2700)?_add_all_x_data_out_index161:10'b0);
   assign  _sub_x_data_in163 = ((_net_3120)?_add_all_x_data_out_index164:10'b0)|
    ((_net_2699)?_add_all_x_data_out_index163:10'b0);
   assign  _sub_x_data_in165 = ((_net_3119)?_add_all_x_data_out_index166:10'b0)|
    ((_net_2698)?_add_all_x_data_out_index165:10'b0);
   assign  _sub_x_data_in167 = ((_net_3118)?_add_all_x_data_out_index168:10'b0)|
    ((_net_2697)?_add_all_x_data_out_index167:10'b0);
   assign  _sub_x_data_in169 = ((_net_3117)?_add_all_x_data_out_index170:10'b0)|
    ((_net_2696)?_add_all_x_data_out_index169:10'b0);
   assign  _sub_x_data_in171 = ((_net_3116)?_add_all_x_data_out_index172:10'b0)|
    ((_net_2695)?_add_all_x_data_out_index171:10'b0);
   assign  _sub_x_data_in173 = ((_net_3115)?_add_all_x_data_out_index174:10'b0)|
    ((_net_2694)?_add_all_x_data_out_index173:10'b0);
   assign  _sub_x_data_in175 = ((_net_3114)?_add_all_x_data_out_index176:10'b0)|
    ((_net_2693)?_add_all_x_data_out_index175:10'b0);
   assign  _sub_x_data_in177 = ((_net_3113)?_add_all_x_data_out_index178:10'b0)|
    ((_net_2692)?_add_all_x_data_out_index177:10'b0);
   assign  _sub_x_data_in179 = ((_net_3112)?_add_all_x_data_out_index180:10'b0)|
    ((_net_2691)?_add_all_x_data_out_index179:10'b0);
   assign  _sub_x_data_in181 = ((_net_3111)?_add_all_x_data_out_index182:10'b0)|
    ((_net_2690)?_add_all_x_data_out_index181:10'b0);
   assign  _sub_x_data_in183 = ((_net_3110)?_add_all_x_data_out_index184:10'b0)|
    ((_net_2689)?_add_all_x_data_out_index183:10'b0);
   assign  _sub_x_data_in185 = ((_net_3109)?_add_all_x_data_out_index186:10'b0)|
    ((_net_2688)?_add_all_x_data_out_index185:10'b0);
   assign  _sub_x_data_in187 = ((_net_3108)?_add_all_x_data_out_index188:10'b0)|
    ((_net_2687)?_add_all_x_data_out_index187:10'b0);
   assign  _sub_x_data_in189 = ((_net_3107)?_add_all_x_data_out_index190:10'b0)|
    ((_net_2686)?_add_all_x_data_out_index189:10'b0);
   assign  _sub_x_data_in193 = ((_net_3106)?_add_all_x_data_out_index193:10'b0)|
    ((_net_2685)?_add_all_x_data_out_index194:10'b0);
   assign  _sub_x_data_in195 = ((_net_3105)?_add_all_x_data_out_index195:10'b0)|
    ((_net_2684)?_add_all_x_data_out_index196:10'b0);
   assign  _sub_x_data_in197 = ((_net_3104)?_add_all_x_data_out_index197:10'b0)|
    ((_net_2683)?_add_all_x_data_out_index198:10'b0);
   assign  _sub_x_data_in199 = ((_net_3103)?_add_all_x_data_out_index199:10'b0)|
    ((_net_2682)?_add_all_x_data_out_index200:10'b0);
   assign  _sub_x_data_in201 = ((_net_3102)?_add_all_x_data_out_index201:10'b0)|
    ((_net_2681)?_add_all_x_data_out_index202:10'b0);
   assign  _sub_x_data_in203 = ((_net_3101)?_add_all_x_data_out_index203:10'b0)|
    ((_net_2680)?_add_all_x_data_out_index204:10'b0);
   assign  _sub_x_data_in205 = ((_net_3100)?_add_all_x_data_out_index205:10'b0)|
    ((_net_2679)?_add_all_x_data_out_index206:10'b0);
   assign  _sub_x_data_in207 = ((_net_3099)?_add_all_x_data_out_index207:10'b0)|
    ((_net_2678)?_add_all_x_data_out_index208:10'b0);
   assign  _sub_x_data_in209 = ((_net_3098)?_add_all_x_data_out_index209:10'b0)|
    ((_net_2677)?_add_all_x_data_out_index210:10'b0);
   assign  _sub_x_data_in211 = ((_net_3097)?_add_all_x_data_out_index211:10'b0)|
    ((_net_2676)?_add_all_x_data_out_index212:10'b0);
   assign  _sub_x_data_in213 = ((_net_3096)?_add_all_x_data_out_index213:10'b0)|
    ((_net_2675)?_add_all_x_data_out_index214:10'b0);
   assign  _sub_x_data_in215 = ((_net_3095)?_add_all_x_data_out_index215:10'b0)|
    ((_net_2674)?_add_all_x_data_out_index216:10'b0);
   assign  _sub_x_data_in217 = ((_net_3094)?_add_all_x_data_out_index217:10'b0)|
    ((_net_2673)?_add_all_x_data_out_index218:10'b0);
   assign  _sub_x_data_in219 = ((_net_3093)?_add_all_x_data_out_index219:10'b0)|
    ((_net_2672)?_add_all_x_data_out_index220:10'b0);
   assign  _sub_x_data_in221 = ((_net_3092)?_add_all_x_data_out_index221:10'b0)|
    ((_net_2671)?_add_all_x_data_out_index222:10'b0);
   assign  _sub_x_data_in225 = ((_net_3091)?_add_all_x_data_out_index226:10'b0)|
    ((_net_2670)?_add_all_x_data_out_index225:10'b0);
   assign  _sub_x_data_in227 = ((_net_3090)?_add_all_x_data_out_index228:10'b0)|
    ((_net_2669)?_add_all_x_data_out_index227:10'b0);
   assign  _sub_x_data_in229 = ((_net_3089)?_add_all_x_data_out_index230:10'b0)|
    ((_net_2668)?_add_all_x_data_out_index229:10'b0);
   assign  _sub_x_data_in231 = ((_net_3088)?_add_all_x_data_out_index232:10'b0)|
    ((_net_2667)?_add_all_x_data_out_index231:10'b0);
   assign  _sub_x_data_in233 = ((_net_3087)?_add_all_x_data_out_index234:10'b0)|
    ((_net_2666)?_add_all_x_data_out_index233:10'b0);
   assign  _sub_x_data_in235 = ((_net_3086)?_add_all_x_data_out_index236:10'b0)|
    ((_net_2665)?_add_all_x_data_out_index235:10'b0);
   assign  _sub_x_data_in237 = ((_net_3085)?_add_all_x_data_out_index238:10'b0)|
    ((_net_2664)?_add_all_x_data_out_index237:10'b0);
   assign  _sub_x_data_in239 = ((_net_3084)?_add_all_x_data_out_index240:10'b0)|
    ((_net_2663)?_add_all_x_data_out_index239:10'b0);
   assign  _sub_x_data_in241 = ((_net_3083)?_add_all_x_data_out_index242:10'b0)|
    ((_net_2662)?_add_all_x_data_out_index241:10'b0);
   assign  _sub_x_data_in243 = ((_net_3082)?_add_all_x_data_out_index244:10'b0)|
    ((_net_2661)?_add_all_x_data_out_index243:10'b0);
   assign  _sub_x_data_in245 = ((_net_3081)?_add_all_x_data_out_index246:10'b0)|
    ((_net_2660)?_add_all_x_data_out_index245:10'b0);
   assign  _sub_x_data_in247 = ((_net_3080)?_add_all_x_data_out_index248:10'b0)|
    ((_net_2659)?_add_all_x_data_out_index247:10'b0);
   assign  _sub_x_data_in249 = ((_net_3079)?_add_all_x_data_out_index250:10'b0)|
    ((_net_2658)?_add_all_x_data_out_index249:10'b0);
   assign  _sub_x_data_in251 = ((_net_3078)?_add_all_x_data_out_index252:10'b0)|
    ((_net_2657)?_add_all_x_data_out_index251:10'b0);
   assign  _sub_x_data_in253 = ((_net_3077)?_add_all_x_data_out_index254:10'b0)|
    ((_net_2656)?_add_all_x_data_out_index253:10'b0);
   assign  _sub_x_data_in257 = ((_net_3076)?_add_all_x_data_out_index257:10'b0)|
    ((_net_2655)?_add_all_x_data_out_index258:10'b0);
   assign  _sub_x_data_in259 = ((_net_3075)?_add_all_x_data_out_index259:10'b0)|
    ((_net_2654)?_add_all_x_data_out_index260:10'b0);
   assign  _sub_x_data_in261 = ((_net_3074)?_add_all_x_data_out_index261:10'b0)|
    ((_net_2653)?_add_all_x_data_out_index262:10'b0);
   assign  _sub_x_data_in263 = ((_net_3073)?_add_all_x_data_out_index263:10'b0)|
    ((_net_2652)?_add_all_x_data_out_index264:10'b0);
   assign  _sub_x_data_in265 = ((_net_3072)?_add_all_x_data_out_index265:10'b0)|
    ((_net_2651)?_add_all_x_data_out_index266:10'b0);
   assign  _sub_x_data_in267 = ((_net_3071)?_add_all_x_data_out_index267:10'b0)|
    ((_net_2650)?_add_all_x_data_out_index268:10'b0);
   assign  _sub_x_data_in269 = ((_net_3070)?_add_all_x_data_out_index269:10'b0)|
    ((_net_2649)?_add_all_x_data_out_index270:10'b0);
   assign  _sub_x_data_in271 = ((_net_3069)?_add_all_x_data_out_index271:10'b0)|
    ((_net_2648)?_add_all_x_data_out_index272:10'b0);
   assign  _sub_x_data_in273 = ((_net_3068)?_add_all_x_data_out_index273:10'b0)|
    ((_net_2647)?_add_all_x_data_out_index274:10'b0);
   assign  _sub_x_data_in275 = ((_net_3067)?_add_all_x_data_out_index275:10'b0)|
    ((_net_2646)?_add_all_x_data_out_index276:10'b0);
   assign  _sub_x_data_in277 = ((_net_3066)?_add_all_x_data_out_index277:10'b0)|
    ((_net_2645)?_add_all_x_data_out_index278:10'b0);
   assign  _sub_x_data_in279 = ((_net_3065)?_add_all_x_data_out_index279:10'b0)|
    ((_net_2644)?_add_all_x_data_out_index280:10'b0);
   assign  _sub_x_data_in281 = ((_net_3064)?_add_all_x_data_out_index281:10'b0)|
    ((_net_2643)?_add_all_x_data_out_index282:10'b0);
   assign  _sub_x_data_in283 = ((_net_3063)?_add_all_x_data_out_index283:10'b0)|
    ((_net_2642)?_add_all_x_data_out_index284:10'b0);
   assign  _sub_x_data_in285 = ((_net_3062)?_add_all_x_data_out_index285:10'b0)|
    ((_net_2641)?_add_all_x_data_out_index286:10'b0);
   assign  _sub_x_data_in289 = ((_net_3061)?_add_all_x_data_out_index290:10'b0)|
    ((_net_2640)?_add_all_x_data_out_index289:10'b0);
   assign  _sub_x_data_in291 = ((_net_3060)?_add_all_x_data_out_index292:10'b0)|
    ((_net_2639)?_add_all_x_data_out_index291:10'b0);
   assign  _sub_x_data_in293 = ((_net_3059)?_add_all_x_data_out_index294:10'b0)|
    ((_net_2638)?_add_all_x_data_out_index293:10'b0);
   assign  _sub_x_data_in295 = ((_net_3058)?_add_all_x_data_out_index296:10'b0)|
    ((_net_2637)?_add_all_x_data_out_index295:10'b0);
   assign  _sub_x_data_in297 = ((_net_3057)?_add_all_x_data_out_index298:10'b0)|
    ((_net_2636)?_add_all_x_data_out_index297:10'b0);
   assign  _sub_x_data_in299 = ((_net_3056)?_add_all_x_data_out_index300:10'b0)|
    ((_net_2635)?_add_all_x_data_out_index299:10'b0);
   assign  _sub_x_data_in301 = ((_net_3055)?_add_all_x_data_out_index302:10'b0)|
    ((_net_2634)?_add_all_x_data_out_index301:10'b0);
   assign  _sub_x_data_in303 = ((_net_3054)?_add_all_x_data_out_index304:10'b0)|
    ((_net_2633)?_add_all_x_data_out_index303:10'b0);
   assign  _sub_x_data_in305 = ((_net_3053)?_add_all_x_data_out_index306:10'b0)|
    ((_net_2632)?_add_all_x_data_out_index305:10'b0);
   assign  _sub_x_data_in307 = ((_net_3052)?_add_all_x_data_out_index308:10'b0)|
    ((_net_2631)?_add_all_x_data_out_index307:10'b0);
   assign  _sub_x_data_in309 = ((_net_3051)?_add_all_x_data_out_index310:10'b0)|
    ((_net_2630)?_add_all_x_data_out_index309:10'b0);
   assign  _sub_x_data_in311 = ((_net_3050)?_add_all_x_data_out_index312:10'b0)|
    ((_net_2629)?_add_all_x_data_out_index311:10'b0);
   assign  _sub_x_data_in313 = ((_net_3049)?_add_all_x_data_out_index314:10'b0)|
    ((_net_2628)?_add_all_x_data_out_index313:10'b0);
   assign  _sub_x_data_in315 = ((_net_3048)?_add_all_x_data_out_index316:10'b0)|
    ((_net_2627)?_add_all_x_data_out_index315:10'b0);
   assign  _sub_x_data_in317 = ((_net_3047)?_add_all_x_data_out_index318:10'b0)|
    ((_net_2626)?_add_all_x_data_out_index317:10'b0);
   assign  _sub_x_data_in321 = ((_net_3046)?_add_all_x_data_out_index321:10'b0)|
    ((_net_2625)?_add_all_x_data_out_index322:10'b0);
   assign  _sub_x_data_in323 = ((_net_3045)?_add_all_x_data_out_index323:10'b0)|
    ((_net_2624)?_add_all_x_data_out_index324:10'b0);
   assign  _sub_x_data_in325 = ((_net_3044)?_add_all_x_data_out_index325:10'b0)|
    ((_net_2623)?_add_all_x_data_out_index326:10'b0);
   assign  _sub_x_data_in327 = ((_net_3043)?_add_all_x_data_out_index327:10'b0)|
    ((_net_2622)?_add_all_x_data_out_index328:10'b0);
   assign  _sub_x_data_in329 = ((_net_3042)?_add_all_x_data_out_index329:10'b0)|
    ((_net_2621)?_add_all_x_data_out_index330:10'b0);
   assign  _sub_x_data_in331 = ((_net_3041)?_add_all_x_data_out_index331:10'b0)|
    ((_net_2620)?_add_all_x_data_out_index332:10'b0);
   assign  _sub_x_data_in333 = ((_net_3040)?_add_all_x_data_out_index333:10'b0)|
    ((_net_2619)?_add_all_x_data_out_index334:10'b0);
   assign  _sub_x_data_in335 = ((_net_3039)?_add_all_x_data_out_index335:10'b0)|
    ((_net_2618)?_add_all_x_data_out_index336:10'b0);
   assign  _sub_x_data_in337 = ((_net_3038)?_add_all_x_data_out_index337:10'b0)|
    ((_net_2617)?_add_all_x_data_out_index338:10'b0);
   assign  _sub_x_data_in339 = ((_net_3037)?_add_all_x_data_out_index339:10'b0)|
    ((_net_2616)?_add_all_x_data_out_index340:10'b0);
   assign  _sub_x_data_in341 = ((_net_3036)?_add_all_x_data_out_index341:10'b0)|
    ((_net_2615)?_add_all_x_data_out_index342:10'b0);
   assign  _sub_x_data_in343 = ((_net_3035)?_add_all_x_data_out_index343:10'b0)|
    ((_net_2614)?_add_all_x_data_out_index344:10'b0);
   assign  _sub_x_data_in345 = ((_net_3034)?_add_all_x_data_out_index345:10'b0)|
    ((_net_2613)?_add_all_x_data_out_index346:10'b0);
   assign  _sub_x_data_in347 = ((_net_3033)?_add_all_x_data_out_index347:10'b0)|
    ((_net_2612)?_add_all_x_data_out_index348:10'b0);
   assign  _sub_x_data_in349 = ((_net_3032)?_add_all_x_data_out_index349:10'b0)|
    ((_net_2611)?_add_all_x_data_out_index350:10'b0);
   assign  _sub_x_data_in353 = ((_net_3031)?_add_all_x_data_out_index354:10'b0)|
    ((_net_2610)?_add_all_x_data_out_index353:10'b0);
   assign  _sub_x_data_in355 = ((_net_3030)?_add_all_x_data_out_index356:10'b0)|
    ((_net_2609)?_add_all_x_data_out_index355:10'b0);
   assign  _sub_x_data_in357 = ((_net_3029)?_add_all_x_data_out_index358:10'b0)|
    ((_net_2608)?_add_all_x_data_out_index357:10'b0);
   assign  _sub_x_data_in359 = ((_net_3028)?_add_all_x_data_out_index360:10'b0)|
    ((_net_2607)?_add_all_x_data_out_index359:10'b0);
   assign  _sub_x_data_in361 = ((_net_3027)?_add_all_x_data_out_index362:10'b0)|
    ((_net_2606)?_add_all_x_data_out_index361:10'b0);
   assign  _sub_x_data_in363 = ((_net_3026)?_add_all_x_data_out_index364:10'b0)|
    ((_net_2605)?_add_all_x_data_out_index363:10'b0);
   assign  _sub_x_data_in365 = ((_net_3025)?_add_all_x_data_out_index366:10'b0)|
    ((_net_2604)?_add_all_x_data_out_index365:10'b0);
   assign  _sub_x_data_in367 = ((_net_3024)?_add_all_x_data_out_index368:10'b0)|
    ((_net_2603)?_add_all_x_data_out_index367:10'b0);
   assign  _sub_x_data_in369 = ((_net_3023)?_add_all_x_data_out_index370:10'b0)|
    ((_net_2602)?_add_all_x_data_out_index369:10'b0);
   assign  _sub_x_data_in371 = ((_net_3022)?_add_all_x_data_out_index372:10'b0)|
    ((_net_2601)?_add_all_x_data_out_index371:10'b0);
   assign  _sub_x_data_in373 = ((_net_3021)?_add_all_x_data_out_index374:10'b0)|
    ((_net_2600)?_add_all_x_data_out_index373:10'b0);
   assign  _sub_x_data_in375 = ((_net_3020)?_add_all_x_data_out_index376:10'b0)|
    ((_net_2599)?_add_all_x_data_out_index375:10'b0);
   assign  _sub_x_data_in377 = ((_net_3019)?_add_all_x_data_out_index378:10'b0)|
    ((_net_2598)?_add_all_x_data_out_index377:10'b0);
   assign  _sub_x_data_in379 = ((_net_3018)?_add_all_x_data_out_index380:10'b0)|
    ((_net_2597)?_add_all_x_data_out_index379:10'b0);
   assign  _sub_x_data_in381 = ((_net_3017)?_add_all_x_data_out_index382:10'b0)|
    ((_net_2596)?_add_all_x_data_out_index381:10'b0);
   assign  _sub_x_data_in385 = ((_net_3016)?_add_all_x_data_out_index385:10'b0)|
    ((_net_2595)?_add_all_x_data_out_index386:10'b0);
   assign  _sub_x_data_in387 = ((_net_3015)?_add_all_x_data_out_index387:10'b0)|
    ((_net_2594)?_add_all_x_data_out_index388:10'b0);
   assign  _sub_x_data_in389 = ((_net_3014)?_add_all_x_data_out_index389:10'b0)|
    ((_net_2593)?_add_all_x_data_out_index390:10'b0);
   assign  _sub_x_data_in391 = ((_net_3013)?_add_all_x_data_out_index391:10'b0)|
    ((_net_2592)?_add_all_x_data_out_index392:10'b0);
   assign  _sub_x_data_in393 = ((_net_3012)?_add_all_x_data_out_index393:10'b0)|
    ((_net_2591)?_add_all_x_data_out_index394:10'b0);
   assign  _sub_x_data_in395 = ((_net_3011)?_add_all_x_data_out_index395:10'b0)|
    ((_net_2590)?_add_all_x_data_out_index396:10'b0);
   assign  _sub_x_data_in397 = ((_net_3010)?_add_all_x_data_out_index397:10'b0)|
    ((_net_2589)?_add_all_x_data_out_index398:10'b0);
   assign  _sub_x_data_in399 = ((_net_3009)?_add_all_x_data_out_index399:10'b0)|
    ((_net_2588)?_add_all_x_data_out_index400:10'b0);
   assign  _sub_x_data_in401 = ((_net_3008)?_add_all_x_data_out_index401:10'b0)|
    ((_net_2587)?_add_all_x_data_out_index402:10'b0);
   assign  _sub_x_data_in403 = ((_net_3007)?_add_all_x_data_out_index403:10'b0)|
    ((_net_2586)?_add_all_x_data_out_index404:10'b0);
   assign  _sub_x_data_in405 = ((_net_3006)?_add_all_x_data_out_index405:10'b0)|
    ((_net_2585)?_add_all_x_data_out_index406:10'b0);
   assign  _sub_x_data_in407 = ((_net_3005)?_add_all_x_data_out_index407:10'b0)|
    ((_net_2584)?_add_all_x_data_out_index408:10'b0);
   assign  _sub_x_data_in409 = ((_net_3004)?_add_all_x_data_out_index409:10'b0)|
    ((_net_2583)?_add_all_x_data_out_index410:10'b0);
   assign  _sub_x_data_in411 = ((_net_3003)?_add_all_x_data_out_index411:10'b0)|
    ((_net_2582)?_add_all_x_data_out_index412:10'b0);
   assign  _sub_x_data_in413 = ((_net_3002)?_add_all_x_data_out_index413:10'b0)|
    ((_net_2581)?_add_all_x_data_out_index414:10'b0);
   assign  _sub_x_data_in417 = ((_net_3001)?_add_all_x_data_out_index418:10'b0)|
    ((_net_2580)?_add_all_x_data_out_index417:10'b0);
   assign  _sub_x_data_in419 = ((_net_3000)?_add_all_x_data_out_index420:10'b0)|
    ((_net_2579)?_add_all_x_data_out_index419:10'b0);
   assign  _sub_x_data_in421 = ((_net_2999)?_add_all_x_data_out_index422:10'b0)|
    ((_net_2578)?_add_all_x_data_out_index421:10'b0);
   assign  _sub_x_data_in423 = ((_net_2998)?_add_all_x_data_out_index424:10'b0)|
    ((_net_2577)?_add_all_x_data_out_index423:10'b0);
   assign  _sub_x_data_in425 = ((_net_2997)?_add_all_x_data_out_index426:10'b0)|
    ((_net_2576)?_add_all_x_data_out_index425:10'b0);
   assign  _sub_x_data_in427 = ((_net_2996)?_add_all_x_data_out_index428:10'b0)|
    ((_net_2575)?_add_all_x_data_out_index427:10'b0);
   assign  _sub_x_data_in429 = ((_net_2995)?_add_all_x_data_out_index430:10'b0)|
    ((_net_2574)?_add_all_x_data_out_index429:10'b0);
   assign  _sub_x_data_in431 = ((_net_2994)?_add_all_x_data_out_index432:10'b0)|
    ((_net_2573)?_add_all_x_data_out_index431:10'b0);
   assign  _sub_x_data_in433 = ((_net_2993)?_add_all_x_data_out_index434:10'b0)|
    ((_net_2572)?_add_all_x_data_out_index433:10'b0);
   assign  _sub_x_data_in435 = ((_net_2992)?_add_all_x_data_out_index436:10'b0)|
    ((_net_2571)?_add_all_x_data_out_index435:10'b0);
   assign  _sub_x_data_in437 = ((_net_2991)?_add_all_x_data_out_index438:10'b0)|
    ((_net_2570)?_add_all_x_data_out_index437:10'b0);
   assign  _sub_x_data_in439 = ((_net_2990)?_add_all_x_data_out_index440:10'b0)|
    ((_net_2569)?_add_all_x_data_out_index439:10'b0);
   assign  _sub_x_data_in441 = ((_net_2989)?_add_all_x_data_out_index442:10'b0)|
    ((_net_2568)?_add_all_x_data_out_index441:10'b0);
   assign  _sub_x_data_in443 = ((_net_2988)?_add_all_x_data_out_index444:10'b0)|
    ((_net_2567)?_add_all_x_data_out_index443:10'b0);
   assign  _sub_x_data_in445 = ((_net_2987)?_add_all_x_data_out_index446:10'b0)|
    ((_net_2566)?_add_all_x_data_out_index445:10'b0);
   assign  _sub_x_data_in449 = ((_net_2986)?_add_all_x_data_out_index449:10'b0)|
    ((_net_2565)?_add_all_x_data_out_index450:10'b0);
   assign  _sub_x_data_in451 = ((_net_2985)?_add_all_x_data_out_index451:10'b0)|
    ((_net_2564)?_add_all_x_data_out_index452:10'b0);
   assign  _sub_x_data_in453 = ((_net_2984)?_add_all_x_data_out_index453:10'b0)|
    ((_net_2563)?_add_all_x_data_out_index454:10'b0);
   assign  _sub_x_data_in455 = ((_net_2983)?_add_all_x_data_out_index455:10'b0)|
    ((_net_2562)?_add_all_x_data_out_index456:10'b0);
   assign  _sub_x_data_in457 = ((_net_2982)?_add_all_x_data_out_index457:10'b0)|
    ((_net_2561)?_add_all_x_data_out_index458:10'b0);
   assign  _sub_x_data_in459 = ((_net_2981)?_add_all_x_data_out_index459:10'b0)|
    ((_net_2560)?_add_all_x_data_out_index460:10'b0);
   assign  _sub_x_data_in461 = ((_net_2980)?_add_all_x_data_out_index461:10'b0)|
    ((_net_2559)?_add_all_x_data_out_index462:10'b0);
   assign  _sub_x_data_in463 = ((_net_2979)?_add_all_x_data_out_index463:10'b0)|
    ((_net_2558)?_add_all_x_data_out_index464:10'b0);
   assign  _sub_x_data_in465 = ((_net_2978)?_add_all_x_data_out_index465:10'b0)|
    ((_net_2557)?_add_all_x_data_out_index466:10'b0);
   assign  _sub_x_data_in467 = ((_net_2977)?_add_all_x_data_out_index467:10'b0)|
    ((_net_2556)?_add_all_x_data_out_index468:10'b0);
   assign  _sub_x_data_in469 = ((_net_2976)?_add_all_x_data_out_index469:10'b0)|
    ((_net_2555)?_add_all_x_data_out_index470:10'b0);
   assign  _sub_x_data_in471 = ((_net_2975)?_add_all_x_data_out_index471:10'b0)|
    ((_net_2554)?_add_all_x_data_out_index472:10'b0);
   assign  _sub_x_data_in473 = ((_net_2974)?_add_all_x_data_out_index473:10'b0)|
    ((_net_2553)?_add_all_x_data_out_index474:10'b0);
   assign  _sub_x_data_in475 = ((_net_2973)?_add_all_x_data_out_index475:10'b0)|
    ((_net_2552)?_add_all_x_data_out_index476:10'b0);
   assign  _sub_x_data_in477 = ((_net_2972)?_add_all_x_data_out_index477:10'b0)|
    ((_net_2551)?_add_all_x_data_out_index478:10'b0);
   assign  _sub_x_data_in_index33 = ((_net_3391)?_add_all_x_data_out34:10'b0)|
    ((_net_2970)?_add_all_x_data_out33:10'b0);
   assign  _sub_x_data_in_index35 = ((_net_3390)?_add_all_x_data_out36:10'b0)|
    ((_net_2969)?_add_all_x_data_out35:10'b0);
   assign  _sub_x_data_in_index37 = ((_net_3389)?_add_all_x_data_out38:10'b0)|
    ((_net_2968)?_add_all_x_data_out37:10'b0);
   assign  _sub_x_data_in_index39 = ((_net_3388)?_add_all_x_data_out40:10'b0)|
    ((_net_2967)?_add_all_x_data_out39:10'b0);
   assign  _sub_x_data_in_index41 = ((_net_3387)?_add_all_x_data_out42:10'b0)|
    ((_net_2966)?_add_all_x_data_out41:10'b0);
   assign  _sub_x_data_in_index43 = ((_net_3386)?_add_all_x_data_out44:10'b0)|
    ((_net_2965)?_add_all_x_data_out43:10'b0);
   assign  _sub_x_data_in_index45 = ((_net_3385)?_add_all_x_data_out46:10'b0)|
    ((_net_2964)?_add_all_x_data_out45:10'b0);
   assign  _sub_x_data_in_index47 = ((_net_3384)?_add_all_x_data_out48:10'b0)|
    ((_net_2963)?_add_all_x_data_out47:10'b0);
   assign  _sub_x_data_in_index49 = ((_net_3383)?_add_all_x_data_out50:10'b0)|
    ((_net_2962)?_add_all_x_data_out49:10'b0);
   assign  _sub_x_data_in_index51 = ((_net_3382)?_add_all_x_data_out52:10'b0)|
    ((_net_2961)?_add_all_x_data_out51:10'b0);
   assign  _sub_x_data_in_index53 = ((_net_3381)?_add_all_x_data_out54:10'b0)|
    ((_net_2960)?_add_all_x_data_out53:10'b0);
   assign  _sub_x_data_in_index55 = ((_net_3380)?_add_all_x_data_out56:10'b0)|
    ((_net_2959)?_add_all_x_data_out55:10'b0);
   assign  _sub_x_data_in_index57 = ((_net_3379)?_add_all_x_data_out58:10'b0)|
    ((_net_2958)?_add_all_x_data_out57:10'b0);
   assign  _sub_x_data_in_index59 = ((_net_3378)?_add_all_x_data_out60:10'b0)|
    ((_net_2957)?_add_all_x_data_out59:10'b0);
   assign  _sub_x_data_in_index61 = ((_net_3377)?_add_all_x_data_out62:10'b0)|
    ((_net_2956)?_add_all_x_data_out61:10'b0);
   assign  _sub_x_data_in_index65 = ((_net_3376)?_add_all_x_data_out65:10'b0)|
    ((_net_2955)?_add_all_x_data_out66:10'b0);
   assign  _sub_x_data_in_index67 = ((_net_3375)?_add_all_x_data_out67:10'b0)|
    ((_net_2954)?_add_all_x_data_out68:10'b0);
   assign  _sub_x_data_in_index69 = ((_net_3374)?_add_all_x_data_out69:10'b0)|
    ((_net_2953)?_add_all_x_data_out70:10'b0);
   assign  _sub_x_data_in_index71 = ((_net_3373)?_add_all_x_data_out71:10'b0)|
    ((_net_2952)?_add_all_x_data_out72:10'b0);
   assign  _sub_x_data_in_index73 = ((_net_3372)?_add_all_x_data_out73:10'b0)|
    ((_net_2951)?_add_all_x_data_out74:10'b0);
   assign  _sub_x_data_in_index75 = ((_net_3371)?_add_all_x_data_out75:10'b0)|
    ((_net_2950)?_add_all_x_data_out76:10'b0);
   assign  _sub_x_data_in_index77 = ((_net_3370)?_add_all_x_data_out77:10'b0)|
    ((_net_2949)?_add_all_x_data_out78:10'b0);
   assign  _sub_x_data_in_index79 = ((_net_3369)?_add_all_x_data_out79:10'b0)|
    ((_net_2948)?_add_all_x_data_out80:10'b0);
   assign  _sub_x_data_in_index81 = ((_net_3368)?_add_all_x_data_out81:10'b0)|
    ((_net_2947)?_add_all_x_data_out82:10'b0);
   assign  _sub_x_data_in_index83 = ((_net_3367)?_add_all_x_data_out83:10'b0)|
    ((_net_2946)?_add_all_x_data_out84:10'b0);
   assign  _sub_x_data_in_index85 = ((_net_3366)?_add_all_x_data_out85:10'b0)|
    ((_net_2945)?_add_all_x_data_out86:10'b0);
   assign  _sub_x_data_in_index87 = ((_net_3365)?_add_all_x_data_out87:10'b0)|
    ((_net_2944)?_add_all_x_data_out88:10'b0);
   assign  _sub_x_data_in_index89 = ((_net_3364)?_add_all_x_data_out89:10'b0)|
    ((_net_2943)?_add_all_x_data_out90:10'b0);
   assign  _sub_x_data_in_index91 = ((_net_3363)?_add_all_x_data_out91:10'b0)|
    ((_net_2942)?_add_all_x_data_out92:10'b0);
   assign  _sub_x_data_in_index93 = ((_net_3362)?_add_all_x_data_out93:10'b0)|
    ((_net_2941)?_add_all_x_data_out94:10'b0);
   assign  _sub_x_data_in_index97 = ((_net_3361)?_add_all_x_data_out98:10'b0)|
    ((_net_2940)?_add_all_x_data_out97:10'b0);
   assign  _sub_x_data_in_index99 = ((_net_3360)?_add_all_x_data_out100:10'b0)|
    ((_net_2939)?_add_all_x_data_out99:10'b0);
   assign  _sub_x_data_in_index101 = ((_net_3359)?_add_all_x_data_out102:10'b0)|
    ((_net_2938)?_add_all_x_data_out101:10'b0);
   assign  _sub_x_data_in_index103 = ((_net_3358)?_add_all_x_data_out104:10'b0)|
    ((_net_2937)?_add_all_x_data_out103:10'b0);
   assign  _sub_x_data_in_index105 = ((_net_3357)?_add_all_x_data_out106:10'b0)|
    ((_net_2936)?_add_all_x_data_out105:10'b0);
   assign  _sub_x_data_in_index107 = ((_net_3356)?_add_all_x_data_out108:10'b0)|
    ((_net_2935)?_add_all_x_data_out107:10'b0);
   assign  _sub_x_data_in_index109 = ((_net_3355)?_add_all_x_data_out110:10'b0)|
    ((_net_2934)?_add_all_x_data_out109:10'b0);
   assign  _sub_x_data_in_index111 = ((_net_3354)?_add_all_x_data_out112:10'b0)|
    ((_net_2933)?_add_all_x_data_out111:10'b0);
   assign  _sub_x_data_in_index113 = ((_net_3353)?_add_all_x_data_out114:10'b0)|
    ((_net_2932)?_add_all_x_data_out113:10'b0);
   assign  _sub_x_data_in_index115 = ((_net_3352)?_add_all_x_data_out116:10'b0)|
    ((_net_2931)?_add_all_x_data_out115:10'b0);
   assign  _sub_x_data_in_index117 = ((_net_3351)?_add_all_x_data_out118:10'b0)|
    ((_net_2930)?_add_all_x_data_out117:10'b0);
   assign  _sub_x_data_in_index119 = ((_net_3350)?_add_all_x_data_out120:10'b0)|
    ((_net_2929)?_add_all_x_data_out119:10'b0);
   assign  _sub_x_data_in_index121 = ((_net_3349)?_add_all_x_data_out122:10'b0)|
    ((_net_2928)?_add_all_x_data_out121:10'b0);
   assign  _sub_x_data_in_index123 = ((_net_3348)?_add_all_x_data_out124:10'b0)|
    ((_net_2927)?_add_all_x_data_out123:10'b0);
   assign  _sub_x_data_in_index125 = ((_net_3347)?_add_all_x_data_out126:10'b0)|
    ((_net_2926)?_add_all_x_data_out125:10'b0);
   assign  _sub_x_data_in_index129 = ((_net_3346)?_add_all_x_data_out129:10'b0)|
    ((_net_2925)?_add_all_x_data_out130:10'b0);
   assign  _sub_x_data_in_index131 = ((_net_3345)?_add_all_x_data_out131:10'b0)|
    ((_net_2924)?_add_all_x_data_out132:10'b0);
   assign  _sub_x_data_in_index133 = ((_net_3344)?_add_all_x_data_out133:10'b0)|
    ((_net_2923)?_add_all_x_data_out134:10'b0);
   assign  _sub_x_data_in_index135 = ((_net_3343)?_add_all_x_data_out135:10'b0)|
    ((_net_2922)?_add_all_x_data_out136:10'b0);
   assign  _sub_x_data_in_index137 = ((_net_3342)?_add_all_x_data_out137:10'b0)|
    ((_net_2921)?_add_all_x_data_out138:10'b0);
   assign  _sub_x_data_in_index139 = ((_net_3341)?_add_all_x_data_out139:10'b0)|
    ((_net_2920)?_add_all_x_data_out140:10'b0);
   assign  _sub_x_data_in_index141 = ((_net_3340)?_add_all_x_data_out141:10'b0)|
    ((_net_2919)?_add_all_x_data_out142:10'b0);
   assign  _sub_x_data_in_index143 = ((_net_3339)?_add_all_x_data_out143:10'b0)|
    ((_net_2918)?_add_all_x_data_out144:10'b0);
   assign  _sub_x_data_in_index145 = ((_net_3338)?_add_all_x_data_out145:10'b0)|
    ((_net_2917)?_add_all_x_data_out146:10'b0);
   assign  _sub_x_data_in_index147 = ((_net_3337)?_add_all_x_data_out147:10'b0)|
    ((_net_2916)?_add_all_x_data_out148:10'b0);
   assign  _sub_x_data_in_index149 = ((_net_3336)?_add_all_x_data_out149:10'b0)|
    ((_net_2915)?_add_all_x_data_out150:10'b0);
   assign  _sub_x_data_in_index151 = ((_net_3335)?_add_all_x_data_out151:10'b0)|
    ((_net_2914)?_add_all_x_data_out152:10'b0);
   assign  _sub_x_data_in_index153 = ((_net_3334)?_add_all_x_data_out153:10'b0)|
    ((_net_2913)?_add_all_x_data_out154:10'b0);
   assign  _sub_x_data_in_index155 = ((_net_3333)?_add_all_x_data_out155:10'b0)|
    ((_net_2912)?_add_all_x_data_out156:10'b0);
   assign  _sub_x_data_in_index157 = ((_net_3332)?_add_all_x_data_out157:10'b0)|
    ((_net_2911)?_add_all_x_data_out158:10'b0);
   assign  _sub_x_data_in_index161 = ((_net_3331)?_add_all_x_data_out162:10'b0)|
    ((_net_2910)?_add_all_x_data_out161:10'b0);
   assign  _sub_x_data_in_index163 = ((_net_3330)?_add_all_x_data_out164:10'b0)|
    ((_net_2909)?_add_all_x_data_out163:10'b0);
   assign  _sub_x_data_in_index165 = ((_net_3329)?_add_all_x_data_out166:10'b0)|
    ((_net_2908)?_add_all_x_data_out165:10'b0);
   assign  _sub_x_data_in_index167 = ((_net_3328)?_add_all_x_data_out168:10'b0)|
    ((_net_2907)?_add_all_x_data_out167:10'b0);
   assign  _sub_x_data_in_index169 = ((_net_3327)?_add_all_x_data_out170:10'b0)|
    ((_net_2906)?_add_all_x_data_out169:10'b0);
   assign  _sub_x_data_in_index171 = ((_net_3326)?_add_all_x_data_out172:10'b0)|
    ((_net_2905)?_add_all_x_data_out171:10'b0);
   assign  _sub_x_data_in_index173 = ((_net_3325)?_add_all_x_data_out174:10'b0)|
    ((_net_2904)?_add_all_x_data_out173:10'b0);
   assign  _sub_x_data_in_index175 = ((_net_3324)?_add_all_x_data_out176:10'b0)|
    ((_net_2903)?_add_all_x_data_out175:10'b0);
   assign  _sub_x_data_in_index177 = ((_net_3323)?_add_all_x_data_out178:10'b0)|
    ((_net_2902)?_add_all_x_data_out177:10'b0);
   assign  _sub_x_data_in_index179 = ((_net_3322)?_add_all_x_data_out180:10'b0)|
    ((_net_2901)?_add_all_x_data_out179:10'b0);
   assign  _sub_x_data_in_index181 = ((_net_3321)?_add_all_x_data_out182:10'b0)|
    ((_net_2900)?_add_all_x_data_out181:10'b0);
   assign  _sub_x_data_in_index183 = ((_net_3320)?_add_all_x_data_out184:10'b0)|
    ((_net_2899)?_add_all_x_data_out183:10'b0);
   assign  _sub_x_data_in_index185 = ((_net_3319)?_add_all_x_data_out186:10'b0)|
    ((_net_2898)?_add_all_x_data_out185:10'b0);
   assign  _sub_x_data_in_index187 = ((_net_3318)?_add_all_x_data_out188:10'b0)|
    ((_net_2897)?_add_all_x_data_out187:10'b0);
   assign  _sub_x_data_in_index189 = ((_net_3317)?_add_all_x_data_out190:10'b0)|
    ((_net_2896)?_add_all_x_data_out189:10'b0);
   assign  _sub_x_data_in_index193 = ((_net_3316)?_add_all_x_data_out193:10'b0)|
    ((_net_2895)?_add_all_x_data_out194:10'b0);
   assign  _sub_x_data_in_index195 = ((_net_3315)?_add_all_x_data_out195:10'b0)|
    ((_net_2894)?_add_all_x_data_out196:10'b0);
   assign  _sub_x_data_in_index197 = ((_net_3314)?_add_all_x_data_out197:10'b0)|
    ((_net_2893)?_add_all_x_data_out198:10'b0);
   assign  _sub_x_data_in_index199 = ((_net_3313)?_add_all_x_data_out199:10'b0)|
    ((_net_2892)?_add_all_x_data_out200:10'b0);
   assign  _sub_x_data_in_index201 = ((_net_3312)?_add_all_x_data_out201:10'b0)|
    ((_net_2891)?_add_all_x_data_out202:10'b0);
   assign  _sub_x_data_in_index203 = ((_net_3311)?_add_all_x_data_out203:10'b0)|
    ((_net_2890)?_add_all_x_data_out204:10'b0);
   assign  _sub_x_data_in_index205 = ((_net_3310)?_add_all_x_data_out205:10'b0)|
    ((_net_2889)?_add_all_x_data_out206:10'b0);
   assign  _sub_x_data_in_index207 = ((_net_3309)?_add_all_x_data_out207:10'b0)|
    ((_net_2888)?_add_all_x_data_out208:10'b0);
   assign  _sub_x_data_in_index209 = ((_net_3308)?_add_all_x_data_out209:10'b0)|
    ((_net_2887)?_add_all_x_data_out210:10'b0);
   assign  _sub_x_data_in_index211 = ((_net_3307)?_add_all_x_data_out211:10'b0)|
    ((_net_2886)?_add_all_x_data_out212:10'b0);
   assign  _sub_x_data_in_index213 = ((_net_3306)?_add_all_x_data_out213:10'b0)|
    ((_net_2885)?_add_all_x_data_out214:10'b0);
   assign  _sub_x_data_in_index215 = ((_net_3305)?_add_all_x_data_out215:10'b0)|
    ((_net_2884)?_add_all_x_data_out216:10'b0);
   assign  _sub_x_data_in_index217 = ((_net_3304)?_add_all_x_data_out217:10'b0)|
    ((_net_2883)?_add_all_x_data_out218:10'b0);
   assign  _sub_x_data_in_index219 = ((_net_3303)?_add_all_x_data_out219:10'b0)|
    ((_net_2882)?_add_all_x_data_out220:10'b0);
   assign  _sub_x_data_in_index221 = ((_net_3302)?_add_all_x_data_out221:10'b0)|
    ((_net_2881)?_add_all_x_data_out222:10'b0);
   assign  _sub_x_data_in_index225 = ((_net_3301)?_add_all_x_data_out226:10'b0)|
    ((_net_2880)?_add_all_x_data_out225:10'b0);
   assign  _sub_x_data_in_index227 = ((_net_3300)?_add_all_x_data_out228:10'b0)|
    ((_net_2879)?_add_all_x_data_out227:10'b0);
   assign  _sub_x_data_in_index229 = ((_net_3299)?_add_all_x_data_out230:10'b0)|
    ((_net_2878)?_add_all_x_data_out229:10'b0);
   assign  _sub_x_data_in_index231 = ((_net_3298)?_add_all_x_data_out232:10'b0)|
    ((_net_2877)?_add_all_x_data_out231:10'b0);
   assign  _sub_x_data_in_index233 = ((_net_3297)?_add_all_x_data_out234:10'b0)|
    ((_net_2876)?_add_all_x_data_out233:10'b0);
   assign  _sub_x_data_in_index235 = ((_net_3296)?_add_all_x_data_out236:10'b0)|
    ((_net_2875)?_add_all_x_data_out235:10'b0);
   assign  _sub_x_data_in_index237 = ((_net_3295)?_add_all_x_data_out238:10'b0)|
    ((_net_2874)?_add_all_x_data_out237:10'b0);
   assign  _sub_x_data_in_index239 = ((_net_3294)?_add_all_x_data_out240:10'b0)|
    ((_net_2873)?_add_all_x_data_out239:10'b0);
   assign  _sub_x_data_in_index241 = ((_net_3293)?_add_all_x_data_out242:10'b0)|
    ((_net_2872)?_add_all_x_data_out241:10'b0);
   assign  _sub_x_data_in_index243 = ((_net_3292)?_add_all_x_data_out244:10'b0)|
    ((_net_2871)?_add_all_x_data_out243:10'b0);
   assign  _sub_x_data_in_index245 = ((_net_3291)?_add_all_x_data_out246:10'b0)|
    ((_net_2870)?_add_all_x_data_out245:10'b0);
   assign  _sub_x_data_in_index247 = ((_net_3290)?_add_all_x_data_out248:10'b0)|
    ((_net_2869)?_add_all_x_data_out247:10'b0);
   assign  _sub_x_data_in_index249 = ((_net_3289)?_add_all_x_data_out250:10'b0)|
    ((_net_2868)?_add_all_x_data_out249:10'b0);
   assign  _sub_x_data_in_index251 = ((_net_3288)?_add_all_x_data_out252:10'b0)|
    ((_net_2867)?_add_all_x_data_out251:10'b0);
   assign  _sub_x_data_in_index253 = ((_net_3287)?_add_all_x_data_out254:10'b0)|
    ((_net_2866)?_add_all_x_data_out253:10'b0);
   assign  _sub_x_data_in_index257 = ((_net_3286)?_add_all_x_data_out257:10'b0)|
    ((_net_2865)?_add_all_x_data_out258:10'b0);
   assign  _sub_x_data_in_index259 = ((_net_3285)?_add_all_x_data_out259:10'b0)|
    ((_net_2864)?_add_all_x_data_out260:10'b0);
   assign  _sub_x_data_in_index261 = ((_net_3284)?_add_all_x_data_out261:10'b0)|
    ((_net_2863)?_add_all_x_data_out262:10'b0);
   assign  _sub_x_data_in_index263 = ((_net_3283)?_add_all_x_data_out263:10'b0)|
    ((_net_2862)?_add_all_x_data_out264:10'b0);
   assign  _sub_x_data_in_index265 = ((_net_3282)?_add_all_x_data_out265:10'b0)|
    ((_net_2861)?_add_all_x_data_out266:10'b0);
   assign  _sub_x_data_in_index267 = ((_net_3281)?_add_all_x_data_out267:10'b0)|
    ((_net_2860)?_add_all_x_data_out268:10'b0);
   assign  _sub_x_data_in_index269 = ((_net_3280)?_add_all_x_data_out269:10'b0)|
    ((_net_2859)?_add_all_x_data_out270:10'b0);
   assign  _sub_x_data_in_index271 = ((_net_3279)?_add_all_x_data_out271:10'b0)|
    ((_net_2858)?_add_all_x_data_out272:10'b0);
   assign  _sub_x_data_in_index273 = ((_net_3278)?_add_all_x_data_out273:10'b0)|
    ((_net_2857)?_add_all_x_data_out274:10'b0);
   assign  _sub_x_data_in_index275 = ((_net_3277)?_add_all_x_data_out275:10'b0)|
    ((_net_2856)?_add_all_x_data_out276:10'b0);
   assign  _sub_x_data_in_index277 = ((_net_3276)?_add_all_x_data_out277:10'b0)|
    ((_net_2855)?_add_all_x_data_out278:10'b0);
   assign  _sub_x_data_in_index279 = ((_net_3275)?_add_all_x_data_out279:10'b0)|
    ((_net_2854)?_add_all_x_data_out280:10'b0);
   assign  _sub_x_data_in_index281 = ((_net_3274)?_add_all_x_data_out281:10'b0)|
    ((_net_2853)?_add_all_x_data_out282:10'b0);
   assign  _sub_x_data_in_index283 = ((_net_3273)?_add_all_x_data_out283:10'b0)|
    ((_net_2852)?_add_all_x_data_out284:10'b0);
   assign  _sub_x_data_in_index285 = ((_net_3272)?_add_all_x_data_out285:10'b0)|
    ((_net_2851)?_add_all_x_data_out286:10'b0);
   assign  _sub_x_data_in_index289 = ((_net_3271)?_add_all_x_data_out290:10'b0)|
    ((_net_2850)?_add_all_x_data_out289:10'b0);
   assign  _sub_x_data_in_index291 = ((_net_3270)?_add_all_x_data_out292:10'b0)|
    ((_net_2849)?_add_all_x_data_out291:10'b0);
   assign  _sub_x_data_in_index293 = ((_net_3269)?_add_all_x_data_out294:10'b0)|
    ((_net_2848)?_add_all_x_data_out293:10'b0);
   assign  _sub_x_data_in_index295 = ((_net_3268)?_add_all_x_data_out296:10'b0)|
    ((_net_2847)?_add_all_x_data_out295:10'b0);
   assign  _sub_x_data_in_index297 = ((_net_3267)?_add_all_x_data_out298:10'b0)|
    ((_net_2846)?_add_all_x_data_out297:10'b0);
   assign  _sub_x_data_in_index299 = ((_net_3266)?_add_all_x_data_out300:10'b0)|
    ((_net_2845)?_add_all_x_data_out299:10'b0);
   assign  _sub_x_data_in_index301 = ((_net_3265)?_add_all_x_data_out302:10'b0)|
    ((_net_2844)?_add_all_x_data_out301:10'b0);
   assign  _sub_x_data_in_index303 = ((_net_3264)?_add_all_x_data_out304:10'b0)|
    ((_net_2843)?_add_all_x_data_out303:10'b0);
   assign  _sub_x_data_in_index305 = ((_net_3263)?_add_all_x_data_out306:10'b0)|
    ((_net_2842)?_add_all_x_data_out305:10'b0);
   assign  _sub_x_data_in_index307 = ((_net_3262)?_add_all_x_data_out308:10'b0)|
    ((_net_2841)?_add_all_x_data_out307:10'b0);
   assign  _sub_x_data_in_index309 = ((_net_3261)?_add_all_x_data_out310:10'b0)|
    ((_net_2840)?_add_all_x_data_out309:10'b0);
   assign  _sub_x_data_in_index311 = ((_net_3260)?_add_all_x_data_out312:10'b0)|
    ((_net_2839)?_add_all_x_data_out311:10'b0);
   assign  _sub_x_data_in_index313 = ((_net_3259)?_add_all_x_data_out314:10'b0)|
    ((_net_2838)?_add_all_x_data_out313:10'b0);
   assign  _sub_x_data_in_index315 = ((_net_3258)?_add_all_x_data_out316:10'b0)|
    ((_net_2837)?_add_all_x_data_out315:10'b0);
   assign  _sub_x_data_in_index317 = ((_net_3257)?_add_all_x_data_out318:10'b0)|
    ((_net_2836)?_add_all_x_data_out317:10'b0);
   assign  _sub_x_data_in_index321 = ((_net_3256)?_add_all_x_data_out321:10'b0)|
    ((_net_2835)?_add_all_x_data_out322:10'b0);
   assign  _sub_x_data_in_index323 = ((_net_3255)?_add_all_x_data_out323:10'b0)|
    ((_net_2834)?_add_all_x_data_out324:10'b0);
   assign  _sub_x_data_in_index325 = ((_net_3254)?_add_all_x_data_out325:10'b0)|
    ((_net_2833)?_add_all_x_data_out326:10'b0);
   assign  _sub_x_data_in_index327 = ((_net_3253)?_add_all_x_data_out327:10'b0)|
    ((_net_2832)?_add_all_x_data_out328:10'b0);
   assign  _sub_x_data_in_index329 = ((_net_3252)?_add_all_x_data_out329:10'b0)|
    ((_net_2831)?_add_all_x_data_out330:10'b0);
   assign  _sub_x_data_in_index331 = ((_net_3251)?_add_all_x_data_out331:10'b0)|
    ((_net_2830)?_add_all_x_data_out332:10'b0);
   assign  _sub_x_data_in_index333 = ((_net_3250)?_add_all_x_data_out333:10'b0)|
    ((_net_2829)?_add_all_x_data_out334:10'b0);
   assign  _sub_x_data_in_index335 = ((_net_3249)?_add_all_x_data_out335:10'b0)|
    ((_net_2828)?_add_all_x_data_out336:10'b0);
   assign  _sub_x_data_in_index337 = ((_net_3248)?_add_all_x_data_out337:10'b0)|
    ((_net_2827)?_add_all_x_data_out338:10'b0);
   assign  _sub_x_data_in_index339 = ((_net_3247)?_add_all_x_data_out339:10'b0)|
    ((_net_2826)?_add_all_x_data_out340:10'b0);
   assign  _sub_x_data_in_index341 = ((_net_3246)?_add_all_x_data_out341:10'b0)|
    ((_net_2825)?_add_all_x_data_out342:10'b0);
   assign  _sub_x_data_in_index343 = ((_net_3245)?_add_all_x_data_out343:10'b0)|
    ((_net_2824)?_add_all_x_data_out344:10'b0);
   assign  _sub_x_data_in_index345 = ((_net_3244)?_add_all_x_data_out345:10'b0)|
    ((_net_2823)?_add_all_x_data_out346:10'b0);
   assign  _sub_x_data_in_index347 = ((_net_3243)?_add_all_x_data_out347:10'b0)|
    ((_net_2822)?_add_all_x_data_out348:10'b0);
   assign  _sub_x_data_in_index349 = ((_net_3242)?_add_all_x_data_out349:10'b0)|
    ((_net_2821)?_add_all_x_data_out350:10'b0);
   assign  _sub_x_data_in_index353 = ((_net_3241)?_add_all_x_data_out354:10'b0)|
    ((_net_2820)?_add_all_x_data_out353:10'b0);
   assign  _sub_x_data_in_index355 = ((_net_3240)?_add_all_x_data_out356:10'b0)|
    ((_net_2819)?_add_all_x_data_out355:10'b0);
   assign  _sub_x_data_in_index357 = ((_net_3239)?_add_all_x_data_out358:10'b0)|
    ((_net_2818)?_add_all_x_data_out357:10'b0);
   assign  _sub_x_data_in_index359 = ((_net_3238)?_add_all_x_data_out360:10'b0)|
    ((_net_2817)?_add_all_x_data_out359:10'b0);
   assign  _sub_x_data_in_index361 = ((_net_3237)?_add_all_x_data_out362:10'b0)|
    ((_net_2816)?_add_all_x_data_out361:10'b0);
   assign  _sub_x_data_in_index363 = ((_net_3236)?_add_all_x_data_out364:10'b0)|
    ((_net_2815)?_add_all_x_data_out363:10'b0);
   assign  _sub_x_data_in_index365 = ((_net_3235)?_add_all_x_data_out366:10'b0)|
    ((_net_2814)?_add_all_x_data_out365:10'b0);
   assign  _sub_x_data_in_index367 = ((_net_3234)?_add_all_x_data_out368:10'b0)|
    ((_net_2813)?_add_all_x_data_out367:10'b0);
   assign  _sub_x_data_in_index369 = ((_net_3233)?_add_all_x_data_out370:10'b0)|
    ((_net_2812)?_add_all_x_data_out369:10'b0);
   assign  _sub_x_data_in_index371 = ((_net_3232)?_add_all_x_data_out372:10'b0)|
    ((_net_2811)?_add_all_x_data_out371:10'b0);
   assign  _sub_x_data_in_index373 = ((_net_3231)?_add_all_x_data_out374:10'b0)|
    ((_net_2810)?_add_all_x_data_out373:10'b0);
   assign  _sub_x_data_in_index375 = ((_net_3230)?_add_all_x_data_out376:10'b0)|
    ((_net_2809)?_add_all_x_data_out375:10'b0);
   assign  _sub_x_data_in_index377 = ((_net_3229)?_add_all_x_data_out378:10'b0)|
    ((_net_2808)?_add_all_x_data_out377:10'b0);
   assign  _sub_x_data_in_index379 = ((_net_3228)?_add_all_x_data_out380:10'b0)|
    ((_net_2807)?_add_all_x_data_out379:10'b0);
   assign  _sub_x_data_in_index381 = ((_net_3227)?_add_all_x_data_out382:10'b0)|
    ((_net_2806)?_add_all_x_data_out381:10'b0);
   assign  _sub_x_data_in_index385 = ((_net_3226)?_add_all_x_data_out385:10'b0)|
    ((_net_2805)?_add_all_x_data_out386:10'b0);
   assign  _sub_x_data_in_index387 = ((_net_3225)?_add_all_x_data_out387:10'b0)|
    ((_net_2804)?_add_all_x_data_out388:10'b0);
   assign  _sub_x_data_in_index389 = ((_net_3224)?_add_all_x_data_out389:10'b0)|
    ((_net_2803)?_add_all_x_data_out390:10'b0);
   assign  _sub_x_data_in_index391 = ((_net_3223)?_add_all_x_data_out391:10'b0)|
    ((_net_2802)?_add_all_x_data_out392:10'b0);
   assign  _sub_x_data_in_index393 = ((_net_3222)?_add_all_x_data_out393:10'b0)|
    ((_net_2801)?_add_all_x_data_out394:10'b0);
   assign  _sub_x_data_in_index395 = ((_net_3221)?_add_all_x_data_out395:10'b0)|
    ((_net_2800)?_add_all_x_data_out396:10'b0);
   assign  _sub_x_data_in_index397 = ((_net_3220)?_add_all_x_data_out397:10'b0)|
    ((_net_2799)?_add_all_x_data_out398:10'b0);
   assign  _sub_x_data_in_index399 = ((_net_3219)?_add_all_x_data_out399:10'b0)|
    ((_net_2798)?_add_all_x_data_out400:10'b0);
   assign  _sub_x_data_in_index401 = ((_net_3218)?_add_all_x_data_out401:10'b0)|
    ((_net_2797)?_add_all_x_data_out402:10'b0);
   assign  _sub_x_data_in_index403 = ((_net_3217)?_add_all_x_data_out403:10'b0)|
    ((_net_2796)?_add_all_x_data_out404:10'b0);
   assign  _sub_x_data_in_index405 = ((_net_3216)?_add_all_x_data_out405:10'b0)|
    ((_net_2795)?_add_all_x_data_out406:10'b0);
   assign  _sub_x_data_in_index407 = ((_net_3215)?_add_all_x_data_out407:10'b0)|
    ((_net_2794)?_add_all_x_data_out408:10'b0);
   assign  _sub_x_data_in_index409 = ((_net_3214)?_add_all_x_data_out409:10'b0)|
    ((_net_2793)?_add_all_x_data_out410:10'b0);
   assign  _sub_x_data_in_index411 = ((_net_3213)?_add_all_x_data_out411:10'b0)|
    ((_net_2792)?_add_all_x_data_out412:10'b0);
   assign  _sub_x_data_in_index413 = ((_net_3212)?_add_all_x_data_out413:10'b0)|
    ((_net_2791)?_add_all_x_data_out414:10'b0);
   assign  _sub_x_data_in_index417 = ((_net_3211)?_add_all_x_data_out418:10'b0)|
    ((_net_2790)?_add_all_x_data_out417:10'b0);
   assign  _sub_x_data_in_index419 = ((_net_3210)?_add_all_x_data_out420:10'b0)|
    ((_net_2789)?_add_all_x_data_out419:10'b0);
   assign  _sub_x_data_in_index421 = ((_net_3209)?_add_all_x_data_out422:10'b0)|
    ((_net_2788)?_add_all_x_data_out421:10'b0);
   assign  _sub_x_data_in_index423 = ((_net_3208)?_add_all_x_data_out424:10'b0)|
    ((_net_2787)?_add_all_x_data_out423:10'b0);
   assign  _sub_x_data_in_index425 = ((_net_3207)?_add_all_x_data_out426:10'b0)|
    ((_net_2786)?_add_all_x_data_out425:10'b0);
   assign  _sub_x_data_in_index427 = ((_net_3206)?_add_all_x_data_out428:10'b0)|
    ((_net_2785)?_add_all_x_data_out427:10'b0);
   assign  _sub_x_data_in_index429 = ((_net_3205)?_add_all_x_data_out430:10'b0)|
    ((_net_2784)?_add_all_x_data_out429:10'b0);
   assign  _sub_x_data_in_index431 = ((_net_3204)?_add_all_x_data_out432:10'b0)|
    ((_net_2783)?_add_all_x_data_out431:10'b0);
   assign  _sub_x_data_in_index433 = ((_net_3203)?_add_all_x_data_out434:10'b0)|
    ((_net_2782)?_add_all_x_data_out433:10'b0);
   assign  _sub_x_data_in_index435 = ((_net_3202)?_add_all_x_data_out436:10'b0)|
    ((_net_2781)?_add_all_x_data_out435:10'b0);
   assign  _sub_x_data_in_index437 = ((_net_3201)?_add_all_x_data_out438:10'b0)|
    ((_net_2780)?_add_all_x_data_out437:10'b0);
   assign  _sub_x_data_in_index439 = ((_net_3200)?_add_all_x_data_out440:10'b0)|
    ((_net_2779)?_add_all_x_data_out439:10'b0);
   assign  _sub_x_data_in_index441 = ((_net_3199)?_add_all_x_data_out442:10'b0)|
    ((_net_2778)?_add_all_x_data_out441:10'b0);
   assign  _sub_x_data_in_index443 = ((_net_3198)?_add_all_x_data_out444:10'b0)|
    ((_net_2777)?_add_all_x_data_out443:10'b0);
   assign  _sub_x_data_in_index445 = ((_net_3197)?_add_all_x_data_out446:10'b0)|
    ((_net_2776)?_add_all_x_data_out445:10'b0);
   assign  _sub_x_data_in_index449 = ((_net_3196)?_add_all_x_data_out449:10'b0)|
    ((_net_2775)?_add_all_x_data_out450:10'b0);
   assign  _sub_x_data_in_index451 = ((_net_3195)?_add_all_x_data_out451:10'b0)|
    ((_net_2774)?_add_all_x_data_out452:10'b0);
   assign  _sub_x_data_in_index453 = ((_net_3194)?_add_all_x_data_out453:10'b0)|
    ((_net_2773)?_add_all_x_data_out454:10'b0);
   assign  _sub_x_data_in_index455 = ((_net_3193)?_add_all_x_data_out455:10'b0)|
    ((_net_2772)?_add_all_x_data_out456:10'b0);
   assign  _sub_x_data_in_index457 = ((_net_3192)?_add_all_x_data_out457:10'b0)|
    ((_net_2771)?_add_all_x_data_out458:10'b0);
   assign  _sub_x_data_in_index459 = ((_net_3191)?_add_all_x_data_out459:10'b0)|
    ((_net_2770)?_add_all_x_data_out460:10'b0);
   assign  _sub_x_data_in_index461 = ((_net_3190)?_add_all_x_data_out461:10'b0)|
    ((_net_2769)?_add_all_x_data_out462:10'b0);
   assign  _sub_x_data_in_index463 = ((_net_3189)?_add_all_x_data_out463:10'b0)|
    ((_net_2768)?_add_all_x_data_out464:10'b0);
   assign  _sub_x_data_in_index465 = ((_net_3188)?_add_all_x_data_out465:10'b0)|
    ((_net_2767)?_add_all_x_data_out466:10'b0);
   assign  _sub_x_data_in_index467 = ((_net_3187)?_add_all_x_data_out467:10'b0)|
    ((_net_2766)?_add_all_x_data_out468:10'b0);
   assign  _sub_x_data_in_index469 = ((_net_3186)?_add_all_x_data_out469:10'b0)|
    ((_net_2765)?_add_all_x_data_out470:10'b0);
   assign  _sub_x_data_in_index471 = ((_net_3185)?_add_all_x_data_out471:10'b0)|
    ((_net_2764)?_add_all_x_data_out472:10'b0);
   assign  _sub_x_data_in_index473 = ((_net_3184)?_add_all_x_data_out473:10'b0)|
    ((_net_2763)?_add_all_x_data_out474:10'b0);
   assign  _sub_x_data_in_index475 = ((_net_3183)?_add_all_x_data_out475:10'b0)|
    ((_net_2762)?_add_all_x_data_out476:10'b0);
   assign  _sub_x_data_in_index477 = ((_net_3182)?_add_all_x_data_out477:10'b0)|
    ((_net_2761)?_add_all_x_data_out478:10'b0);
   assign  _sub_x_subs_exe = (_net_2971|_net_2550);
   assign  _sub_x_p_reset = p_reset;
   assign  _sub_x_m_clock = m_clock;
   assign  _net_4 = ((((((kanwa_exit < 2'b10)|(dig_exit==1'b0))&(start_reg != (goal_reg-10'b0000000001)))&(start_reg != (goal_reg+10'b0000000001)))&(start_reg != (goal_reg-10'b0000100000)))&(start_reg != (goal_reg+10'b0000100000)));
   assign  _net_5 = (_reg_1&_net_4);
   assign  _net_6 = (_reg_1&_net_4);
   assign  _net_7 = (_reg_1&_net_4);
   assign  _net_8 = (_reg_1&_net_4);
   assign  _net_9 = (_reg_1&_net_4);
   assign  _net_10 = (_reg_1&_net_4);
   assign  _net_11 = (_reg_1&_net_4);
   assign  _net_12 = (_reg_1&_net_4);
   assign  _net_13 = (_reg_1&_net_4);
   assign  _net_14 = (_reg_1&_net_4);
   assign  _net_15 = (_reg_1&_net_4);
   assign  _net_16 = (_reg_1&_net_4);
   assign  _net_17 = (_reg_1&_net_4);
   assign  _net_18 = (_reg_1&_net_4);
   assign  _net_19 = (_reg_1&_net_4);
   assign  _net_20 = (_reg_1&_net_4);
   assign  _net_21 = (_reg_1&_net_4);
   assign  _net_22 = (_reg_1&_net_4);
   assign  _net_23 = (_reg_1&_net_4);
   assign  _net_24 = (_reg_1&_net_4);
   assign  _net_25 = (_reg_1&_net_4);
   assign  _net_26 = (_reg_1&_net_4);
   assign  _net_27 = (_reg_1&_net_4);
   assign  _net_28 = (_reg_1&_net_4);
   assign  _net_29 = (_reg_1&_net_4);
   assign  _net_30 = (_reg_1&_net_4);
   assign  _net_31 = (_reg_1&_net_4);
   assign  _net_32 = (_reg_1&_net_4);
   assign  _net_33 = (_reg_1&_net_4);
   assign  _net_34 = (_reg_1&_net_4);
   assign  _net_35 = (_reg_1&_net_4);
   assign  _net_36 = (_reg_1&_net_4);
   assign  _net_37 = (_reg_1&_net_4);
   assign  _net_38 = (_reg_1&_net_4);
   assign  _net_39 = (_reg_1&_net_4);
   assign  _net_40 = (_reg_1&_net_4);
   assign  _net_41 = (_reg_1&_net_4);
   assign  _net_42 = (_reg_1&_net_4);
   assign  _net_43 = (_reg_1&_net_4);
   assign  _net_44 = (_reg_1&_net_4);
   assign  _net_45 = (_reg_1&_net_4);
   assign  _net_46 = (_reg_1&_net_4);
   assign  _net_47 = (_reg_1&_net_4);
   assign  _net_48 = (_reg_1&_net_4);
   assign  _net_49 = (_reg_1&_net_4);
   assign  _net_50 = (_reg_1&_net_4);
   assign  _net_51 = (_reg_1&_net_4);
   assign  _net_52 = (_reg_1&_net_4);
   assign  _net_53 = (_reg_1&_net_4);
   assign  _net_54 = (_reg_1&_net_4);
   assign  _net_55 = (_reg_1&_net_4);
   assign  _net_56 = (_reg_1&_net_4);
   assign  _net_57 = (_reg_1&_net_4);
   assign  _net_58 = (_reg_1&_net_4);
   assign  _net_59 = (_reg_1&_net_4);
   assign  _net_60 = (_reg_1&_net_4);
   assign  _net_61 = (_reg_1&_net_4);
   assign  _net_62 = (_reg_1&_net_4);
   assign  _net_63 = (_reg_1&_net_4);
   assign  _net_64 = (_reg_1&_net_4);
   assign  _net_65 = (_reg_1&_net_4);
   assign  _net_66 = (_reg_1&_net_4);
   assign  _net_67 = (_reg_1&_net_4);
   assign  _net_68 = (_reg_1&_net_4);
   assign  _net_69 = (_reg_1&_net_4);
   assign  _net_70 = (_reg_1&_net_4);
   assign  _net_71 = (_reg_1&_net_4);
   assign  _net_72 = (_reg_1&_net_4);
   assign  _net_73 = (_reg_1&_net_4);
   assign  _net_74 = (_reg_1&_net_4);
   assign  _net_75 = (_reg_1&_net_4);
   assign  _net_76 = (_reg_1&_net_4);
   assign  _net_77 = (_reg_1&_net_4);
   assign  _net_78 = (_reg_1&_net_4);
   assign  _net_79 = (_reg_1&_net_4);
   assign  _net_80 = (_reg_1&_net_4);
   assign  _net_81 = (_reg_1&_net_4);
   assign  _net_82 = (_reg_1&_net_4);
   assign  _net_83 = (_reg_1&_net_4);
   assign  _net_84 = (_reg_1&_net_4);
   assign  _net_85 = (_reg_1&_net_4);
   assign  _net_86 = (_reg_1&_net_4);
   assign  _net_87 = (_reg_1&_net_4);
   assign  _net_88 = (_reg_1&_net_4);
   assign  _net_89 = (_reg_1&_net_4);
   assign  _net_90 = (_reg_1&_net_4);
   assign  _net_91 = (_reg_1&_net_4);
   assign  _net_92 = (_reg_1&_net_4);
   assign  _net_93 = (_reg_1&_net_4);
   assign  _net_94 = (_reg_1&_net_4);
   assign  _net_95 = (_reg_1&_net_4);
   assign  _net_96 = (_reg_1&_net_4);
   assign  _net_97 = (_reg_1&_net_4);
   assign  _net_98 = (_reg_1&_net_4);
   assign  _net_99 = (_reg_1&_net_4);
   assign  _net_100 = (_reg_1&_net_4);
   assign  _net_101 = (_reg_1&_net_4);
   assign  _net_102 = (_reg_1&_net_4);
   assign  _net_103 = (_reg_1&_net_4);
   assign  _net_104 = (_reg_1&_net_4);
   assign  _net_105 = (_reg_1&_net_4);
   assign  _net_106 = (_reg_1&_net_4);
   assign  _net_107 = (_reg_1&_net_4);
   assign  _net_108 = (_reg_1&_net_4);
   assign  _net_109 = (_reg_1&_net_4);
   assign  _net_110 = (_reg_1&_net_4);
   assign  _net_111 = (_reg_1&_net_4);
   assign  _net_112 = (_reg_1&_net_4);
   assign  _net_113 = (_reg_1&_net_4);
   assign  _net_114 = (_reg_1&_net_4);
   assign  _net_115 = (_reg_1&_net_4);
   assign  _net_116 = (_reg_1&_net_4);
   assign  _net_117 = (_reg_1&_net_4);
   assign  _net_118 = (_reg_1&_net_4);
   assign  _net_119 = (_reg_1&_net_4);
   assign  _net_120 = (_reg_1&_net_4);
   assign  _net_121 = (_reg_1&_net_4);
   assign  _net_122 = (_reg_1&_net_4);
   assign  _net_123 = (_reg_1&_net_4);
   assign  _net_124 = (_reg_1&_net_4);
   assign  _net_125 = (_reg_1&_net_4);
   assign  _net_126 = (_reg_1&_net_4);
   assign  _net_127 = (_reg_1&_net_4);
   assign  _net_128 = (_reg_1&_net_4);
   assign  _net_129 = (_reg_1&_net_4);
   assign  _net_130 = (_reg_1&_net_4);
   assign  _net_131 = (_reg_1&_net_4);
   assign  _net_132 = (_reg_1&_net_4);
   assign  _net_133 = (_reg_1&_net_4);
   assign  _net_134 = (_reg_1&_net_4);
   assign  _net_135 = (_reg_1&_net_4);
   assign  _net_136 = (_reg_1&_net_4);
   assign  _net_137 = (_reg_1&_net_4);
   assign  _net_138 = (_reg_1&_net_4);
   assign  _net_139 = (_reg_1&_net_4);
   assign  _net_140 = (_reg_1&_net_4);
   assign  _net_141 = (_reg_1&_net_4);
   assign  _net_142 = (_reg_1&_net_4);
   assign  _net_143 = (_reg_1&_net_4);
   assign  _net_144 = (_reg_1&_net_4);
   assign  _net_145 = (_reg_1&_net_4);
   assign  _net_146 = (_reg_1&_net_4);
   assign  _net_147 = (_reg_1&_net_4);
   assign  _net_148 = (_reg_1&_net_4);
   assign  _net_149 = (_reg_1&_net_4);
   assign  _net_150 = (_reg_1&_net_4);
   assign  _net_151 = (_reg_1&_net_4);
   assign  _net_152 = (_reg_1&_net_4);
   assign  _net_153 = (_reg_1&_net_4);
   assign  _net_154 = (_reg_1&_net_4);
   assign  _net_155 = (_reg_1&_net_4);
   assign  _net_156 = (_reg_1&_net_4);
   assign  _net_157 = (_reg_1&_net_4);
   assign  _net_158 = (_reg_1&_net_4);
   assign  _net_159 = (_reg_1&_net_4);
   assign  _net_160 = (_reg_1&_net_4);
   assign  _net_161 = (_reg_1&_net_4);
   assign  _net_162 = (_reg_1&_net_4);
   assign  _net_163 = (_reg_1&_net_4);
   assign  _net_164 = (_reg_1&_net_4);
   assign  _net_165 = (_reg_1&_net_4);
   assign  _net_166 = (_reg_1&_net_4);
   assign  _net_167 = (_reg_1&_net_4);
   assign  _net_168 = (_reg_1&_net_4);
   assign  _net_169 = (_reg_1&_net_4);
   assign  _net_170 = (_reg_1&_net_4);
   assign  _net_171 = (_reg_1&_net_4);
   assign  _net_172 = (_reg_1&_net_4);
   assign  _net_173 = (_reg_1&_net_4);
   assign  _net_174 = (_reg_1&_net_4);
   assign  _net_175 = (_reg_1&_net_4);
   assign  _net_176 = (_reg_1&_net_4);
   assign  _net_177 = (_reg_1&_net_4);
   assign  _net_178 = (_reg_1&_net_4);
   assign  _net_179 = (_reg_1&_net_4);
   assign  _net_180 = (_reg_1&_net_4);
   assign  _net_181 = (_reg_1&_net_4);
   assign  _net_182 = (_reg_1&_net_4);
   assign  _net_183 = (_reg_1&_net_4);
   assign  _net_184 = (_reg_1&_net_4);
   assign  _net_185 = (_reg_1&_net_4);
   assign  _net_186 = (_reg_1&_net_4);
   assign  _net_187 = (_reg_1&_net_4);
   assign  _net_188 = (_reg_1&_net_4);
   assign  _net_189 = (_reg_1&_net_4);
   assign  _net_190 = (_reg_1&_net_4);
   assign  _net_191 = (_reg_1&_net_4);
   assign  _net_192 = (_reg_1&_net_4);
   assign  _net_193 = (_reg_1&_net_4);
   assign  _net_194 = (_reg_1&_net_4);
   assign  _net_195 = (_reg_1&_net_4);
   assign  _net_196 = (_reg_1&_net_4);
   assign  _net_197 = (_reg_1&_net_4);
   assign  _net_198 = (_reg_1&_net_4);
   assign  _net_199 = (_reg_1&_net_4);
   assign  _net_200 = (_reg_1&_net_4);
   assign  _net_201 = (_reg_1&_net_4);
   assign  _net_202 = (_reg_1&_net_4);
   assign  _net_203 = (_reg_1&_net_4);
   assign  _net_204 = (_reg_1&_net_4);
   assign  _net_205 = (_reg_1&_net_4);
   assign  _net_206 = (_reg_1&_net_4);
   assign  _net_207 = (_reg_1&_net_4);
   assign  _net_208 = (_reg_1&_net_4);
   assign  _net_209 = (_reg_1&_net_4);
   assign  _net_210 = (_reg_1&_net_4);
   assign  _net_211 = (_reg_1&_net_4);
   assign  _net_212 = (_reg_1&_net_4);
   assign  _net_213 = (_reg_1&_net_4);
   assign  _net_214 = (_reg_1&_net_4);
   assign  _net_215 = (_reg_1&_net_4);
   assign  _net_216 = (_reg_1&_net_4);
   assign  _net_217 = (_reg_1&_net_4);
   assign  _net_218 = (_reg_1&_net_4);
   assign  _net_219 = (_reg_1&_net_4);
   assign  _net_220 = (_reg_1&_net_4);
   assign  _net_221 = (_reg_1&_net_4);
   assign  _net_222 = (_reg_1&_net_4);
   assign  _net_223 = (_reg_1&_net_4);
   assign  _net_224 = (_reg_1&_net_4);
   assign  _net_225 = (_reg_1&_net_4);
   assign  _net_226 = (_reg_1&_net_4);
   assign  _net_227 = (_reg_1&_net_4);
   assign  _net_228 = (_reg_1&_net_4);
   assign  _net_229 = (_reg_1&_net_4);
   assign  _net_230 = (_reg_1&_net_4);
   assign  _net_231 = (_reg_1&_net_4);
   assign  _net_232 = (_reg_1&_net_4);
   assign  _net_233 = (_reg_1&_net_4);
   assign  _net_234 = (_reg_1&_net_4);
   assign  _net_235 = (_reg_1&_net_4);
   assign  _net_236 = (_reg_1&_net_4);
   assign  _net_237 = (_reg_1&_net_4);
   assign  _net_238 = (_reg_1&_net_4);
   assign  _net_239 = (_reg_1&_net_4);
   assign  _net_240 = (_reg_1&_net_4);
   assign  _net_241 = (_reg_1&_net_4);
   assign  _net_242 = (_reg_1&_net_4);
   assign  _net_243 = (_reg_1&_net_4);
   assign  _net_244 = (_reg_1&_net_4);
   assign  _net_245 = (_reg_1&_net_4);
   assign  _net_246 = (_reg_1&_net_4);
   assign  _net_247 = (_reg_1&_net_4);
   assign  _net_248 = (_reg_1&_net_4);
   assign  _net_249 = (_reg_1&_net_4);
   assign  _net_250 = (_reg_1&_net_4);
   assign  _net_251 = (_reg_1&_net_4);
   assign  _net_252 = (_reg_1&_net_4);
   assign  _net_253 = (_reg_1&_net_4);
   assign  _net_254 = (_reg_1&_net_4);
   assign  _net_255 = (_reg_1&_net_4);
   assign  _net_256 = (_reg_1&_net_4);
   assign  _net_257 = (_reg_1&_net_4);
   assign  _net_258 = (_reg_1&_net_4);
   assign  _net_259 = (_reg_1&_net_4);
   assign  _net_260 = (_reg_1&_net_4);
   assign  _net_261 = (_reg_1&_net_4);
   assign  _net_262 = (_reg_1&_net_4);
   assign  _net_263 = (_reg_1&_net_4);
   assign  _net_264 = (_reg_1&_net_4);
   assign  _net_265 = (_reg_1&_net_4);
   assign  _net_266 = (_reg_1&_net_4);
   assign  _net_267 = (_reg_1&_net_4);
   assign  _net_268 = (_reg_1&_net_4);
   assign  _net_269 = (_reg_1&_net_4);
   assign  _net_270 = (_reg_1&_net_4);
   assign  _net_271 = (_reg_1&_net_4);
   assign  _net_272 = (_reg_1&_net_4);
   assign  _net_273 = (_reg_1&_net_4);
   assign  _net_274 = (_reg_1&_net_4);
   assign  _net_275 = (_reg_1&_net_4);
   assign  _net_276 = (_reg_1&_net_4);
   assign  _net_277 = (_reg_1&_net_4);
   assign  _net_278 = (_reg_1&_net_4);
   assign  _net_279 = (_reg_1&_net_4);
   assign  _net_280 = (_reg_1&_net_4);
   assign  _net_281 = (_reg_1&_net_4);
   assign  _net_282 = (_reg_1&_net_4);
   assign  _net_283 = (_reg_1&_net_4);
   assign  _net_284 = (_reg_1&_net_4);
   assign  _net_285 = (_reg_1&_net_4);
   assign  _net_286 = (_reg_1&_net_4);
   assign  _net_287 = (_reg_1&_net_4);
   assign  _net_288 = (_reg_1&_net_4);
   assign  _net_289 = (_reg_1&_net_4);
   assign  _net_290 = (_reg_1&_net_4);
   assign  _net_291 = (_reg_1&_net_4);
   assign  _net_292 = (_reg_1&_net_4);
   assign  _net_293 = (_reg_1&_net_4);
   assign  _net_294 = (_reg_1&_net_4);
   assign  _net_295 = (_reg_1&_net_4);
   assign  _net_296 = (_reg_1&_net_4);
   assign  _net_297 = (_reg_1&_net_4);
   assign  _net_298 = (_reg_1&_net_4);
   assign  _net_299 = (_reg_1&_net_4);
   assign  _net_300 = (_reg_1&_net_4);
   assign  _net_301 = (_reg_1&_net_4);
   assign  _net_302 = (_reg_1&_net_4);
   assign  _net_303 = (_reg_1&_net_4);
   assign  _net_304 = (_reg_1&_net_4);
   assign  _net_305 = (_reg_1&_net_4);
   assign  _net_306 = (_reg_1&_net_4);
   assign  _net_307 = (_reg_1&_net_4);
   assign  _net_308 = (_reg_1&_net_4);
   assign  _net_309 = (_reg_1&_net_4);
   assign  _net_310 = (_reg_1&_net_4);
   assign  _net_311 = (_reg_1&_net_4);
   assign  _net_312 = (_reg_1&_net_4);
   assign  _net_313 = (_reg_1&_net_4);
   assign  _net_314 = (_reg_1&_net_4);
   assign  _net_315 = (_reg_1&_net_4);
   assign  _net_316 = (_reg_1&_net_4);
   assign  _net_317 = (_reg_1&_net_4);
   assign  _net_318 = (_reg_1&_net_4);
   assign  _net_319 = (_reg_1&_net_4);
   assign  _net_320 = (_reg_1&_net_4);
   assign  _net_321 = (_reg_1&_net_4);
   assign  _net_322 = (_reg_1&_net_4);
   assign  _net_323 = (_reg_1&_net_4);
   assign  _net_324 = (_reg_1&_net_4);
   assign  _net_325 = (_reg_1&_net_4);
   assign  _net_326 = (_reg_1&_net_4);
   assign  _net_327 = (_reg_1&_net_4);
   assign  _net_328 = (_reg_1&_net_4);
   assign  _net_329 = (_reg_1&_net_4);
   assign  _net_330 = (_reg_1&_net_4);
   assign  _net_331 = (_reg_1&_net_4);
   assign  _net_332 = (_reg_1&_net_4);
   assign  _net_333 = (_reg_1&_net_4);
   assign  _net_334 = (_reg_1&_net_4);
   assign  _net_335 = (_reg_1&_net_4);
   assign  _net_336 = (_reg_1&_net_4);
   assign  _net_337 = (_reg_1&_net_4);
   assign  _net_338 = (_reg_1&_net_4);
   assign  _net_339 = (_reg_1&_net_4);
   assign  _net_340 = (_reg_1&_net_4);
   assign  _net_341 = (_reg_1&_net_4);
   assign  _net_342 = (_reg_1&_net_4);
   assign  _net_343 = (_reg_1&_net_4);
   assign  _net_344 = (_reg_1&_net_4);
   assign  _net_345 = (_reg_1&_net_4);
   assign  _net_346 = (_reg_1&_net_4);
   assign  _net_347 = (_reg_1&_net_4);
   assign  _net_348 = (_reg_1&_net_4);
   assign  _net_349 = (_reg_1&_net_4);
   assign  _net_350 = (_reg_1&_net_4);
   assign  _net_351 = (_reg_1&_net_4);
   assign  _net_352 = (_reg_1&_net_4);
   assign  _net_353 = (_reg_1&_net_4);
   assign  _net_354 = (_reg_1&_net_4);
   assign  _net_355 = (_reg_1&_net_4);
   assign  _net_356 = (_reg_1&_net_4);
   assign  _net_357 = (_reg_1&_net_4);
   assign  _net_358 = (_reg_1&_net_4);
   assign  _net_359 = (_reg_1&_net_4);
   assign  _net_360 = (_reg_1&_net_4);
   assign  _net_361 = (_reg_1&_net_4);
   assign  _net_362 = (_reg_1&_net_4);
   assign  _net_363 = (_reg_1&_net_4);
   assign  _net_364 = (_reg_1&_net_4);
   assign  _net_365 = (_reg_1&_net_4);
   assign  _net_366 = (_reg_1&_net_4);
   assign  _net_367 = (_reg_1&_net_4);
   assign  _net_368 = (_reg_1&_net_4);
   assign  _net_369 = (_reg_1&_net_4);
   assign  _net_370 = (_reg_1&_net_4);
   assign  _net_371 = (_reg_1&_net_4);
   assign  _net_372 = (_reg_1&_net_4);
   assign  _net_373 = (_reg_1&_net_4);
   assign  _net_374 = (_reg_1&_net_4);
   assign  _net_375 = (_reg_1&_net_4);
   assign  _net_376 = (_reg_1&_net_4);
   assign  _net_377 = (_reg_1&_net_4);
   assign  _net_378 = (_reg_1&_net_4);
   assign  _net_379 = (_reg_1&_net_4);
   assign  _net_380 = (_reg_1&_net_4);
   assign  _net_381 = (_reg_1&_net_4);
   assign  _net_382 = (_reg_1&_net_4);
   assign  _net_383 = (_reg_1&_net_4);
   assign  _net_384 = (_reg_1&_net_4);
   assign  _net_385 = (_reg_1&_net_4);
   assign  _net_386 = (_reg_1&_net_4);
   assign  _net_387 = (_reg_1&_net_4);
   assign  _net_388 = (_reg_1&_net_4);
   assign  _net_389 = (_reg_1&_net_4);
   assign  _net_390 = (_reg_1&_net_4);
   assign  _net_391 = (_reg_1&_net_4);
   assign  _net_392 = (_reg_1&_net_4);
   assign  _net_393 = (_reg_1&_net_4);
   assign  _net_394 = (_reg_1&_net_4);
   assign  _net_395 = (_reg_1&_net_4);
   assign  _net_396 = (_reg_1&_net_4);
   assign  _net_397 = (_reg_1&_net_4);
   assign  _net_398 = (_reg_1&_net_4);
   assign  _net_399 = (_reg_1&_net_4);
   assign  _net_400 = (_reg_1&_net_4);
   assign  _net_401 = (_reg_1&_net_4);
   assign  _net_402 = (_reg_1&_net_4);
   assign  _net_403 = (_reg_1&_net_4);
   assign  _net_404 = (_reg_1&_net_4);
   assign  _net_405 = (_reg_1&_net_4);
   assign  _net_406 = (_reg_1&_net_4);
   assign  _net_407 = (_reg_1&_net_4);
   assign  _net_408 = (_reg_1&_net_4);
   assign  _net_409 = (_reg_1&_net_4);
   assign  _net_410 = (_reg_1&_net_4);
   assign  _net_411 = (_reg_1&_net_4);
   assign  _net_412 = (_reg_1&_net_4);
   assign  _net_413 = (_reg_1&_net_4);
   assign  _net_414 = (_reg_1&_net_4);
   assign  _net_415 = (_reg_1&_net_4);
   assign  _net_416 = (_reg_1&_net_4);
   assign  _net_417 = (_reg_1&_net_4);
   assign  _net_418 = (_reg_1&_net_4);
   assign  _net_419 = (_reg_1&_net_4);
   assign  _net_420 = (_reg_1&_net_4);
   assign  _net_421 = (_reg_1&_net_4);
   assign  _net_422 = (_reg_1&_net_4);
   assign  _net_423 = (_reg_1&_net_4);
   assign  _net_424 = (_reg_1&_net_4);
   assign  _net_425 = (_reg_1&_net_4);
   assign  _net_426 = (_reg_1&_net_4);
   assign  _net_427 = (_reg_1&_net_4);
   assign  _net_428 = (_reg_1&_net_4);
   assign  _net_429 = (_reg_1&_net_4);
   assign  _net_430 = (_reg_1&_net_4);
   assign  _net_431 = (_reg_1&_net_4);
   assign  _net_432 = (_reg_1&_net_4);
   assign  _net_433 = (_reg_1&_net_4);
   assign  _net_434 = (_reg_1&_net_4);
   assign  _net_435 = (_reg_1&_net_4);
   assign  _net_436 = (_reg_1&_net_4);
   assign  _net_437 = (_reg_1&_net_4);
   assign  _net_438 = (_reg_1&_net_4);
   assign  _net_439 = (_reg_1&_net_4);
   assign  _net_440 = (_reg_1&_net_4);
   assign  _net_441 = (_reg_1&_net_4);
   assign  _net_442 = (_reg_1&_net_4);
   assign  _net_443 = (_reg_1&_net_4);
   assign  _net_444 = (_reg_1&_net_4);
   assign  _net_445 = (_reg_1&_net_4);
   assign  _net_446 = (_reg_1&_net_4);
   assign  _net_447 = (_reg_1&_net_4);
   assign  _net_448 = (_reg_1&_net_4);
   assign  _net_449 = (_reg_1&_net_4);
   assign  _net_450 = (_reg_1&_net_4);
   assign  _net_451 = (_reg_1&_net_4);
   assign  _net_452 = (_reg_1&_net_4);
   assign  _net_453 = (_reg_1&_net_4);
   assign  _net_454 = (_reg_1&_net_4);
   assign  _net_455 = (_reg_1&_net_4);
   assign  _net_456 = (_reg_1&_net_4);
   assign  _net_457 = (_reg_1&_net_4);
   assign  _net_458 = (_reg_1&_net_4);
   assign  _net_459 = (_reg_1&_net_4);
   assign  _net_460 = (_reg_1&_net_4);
   assign  _net_461 = (_reg_1&_net_4);
   assign  _net_462 = (_reg_1&_net_4);
   assign  _net_463 = (_reg_1&_net_4);
   assign  _net_464 = (_reg_1&_net_4);
   assign  _net_465 = (_reg_1&_net_4);
   assign  _net_466 = (_reg_1&_net_4);
   assign  _net_467 = (_reg_1&_net_4);
   assign  _net_468 = (_reg_1&_net_4);
   assign  _net_469 = (_reg_1&_net_4);
   assign  _net_470 = (_reg_1&_net_4);
   assign  _net_471 = (_reg_1&_net_4);
   assign  _net_472 = (_reg_1&_net_4);
   assign  _net_473 = (_reg_1&_net_4);
   assign  _net_474 = (_reg_1&_net_4);
   assign  _net_475 = (_reg_1&_net_4);
   assign  _net_476 = (_reg_1&_net_4);
   assign  _net_477 = (_reg_1&_net_4);
   assign  _net_478 = (_reg_1&_net_4);
   assign  _net_479 = (_reg_1&_net_4);
   assign  _net_480 = (_reg_1&_net_4);
   assign  _net_481 = (_reg_1&_net_4);
   assign  _net_482 = (_reg_1&_net_4);
   assign  _net_483 = (_reg_1&_net_4);
   assign  _net_484 = (_reg_1&_net_4);
   assign  _net_485 = (_reg_1&_net_4);
   assign  _net_486 = (_reg_1&_net_4);
   assign  _net_487 = (_reg_1&_net_4);
   assign  _net_488 = (_reg_1&_net_4);
   assign  _net_489 = (_reg_1&_net_4);
   assign  _net_490 = (_reg_1&_net_4);
   assign  _net_491 = (_reg_1&_net_4);
   assign  _net_492 = (_reg_1&_net_4);
   assign  _net_493 = (_reg_1&_net_4);
   assign  _net_494 = (_reg_1&_net_4);
   assign  _net_495 = (_reg_1&_net_4);
   assign  _net_496 = (_reg_1&_net_4);
   assign  _net_497 = (_reg_1&_net_4);
   assign  _net_498 = (_reg_1&_net_4);
   assign  _net_499 = (_reg_1&_net_4);
   assign  _net_500 = (_reg_1&_net_4);
   assign  _net_501 = (_reg_1&_net_4);
   assign  _net_502 = (_reg_1&_net_4);
   assign  _net_503 = (_reg_1&_net_4);
   assign  _net_504 = (_reg_1&_net_4);
   assign  _net_505 = (_reg_1&_net_4);
   assign  _net_506 = (_reg_1&_net_4);
   assign  _net_507 = (_reg_1&_net_4);
   assign  _net_508 = (_reg_1&_net_4);
   assign  _net_509 = (_reg_1&_net_4);
   assign  _net_510 = (_reg_1&_net_4);
   assign  _net_511 = (_reg_1&_net_4);
   assign  _net_512 = (_reg_1&_net_4);
   assign  _net_513 = (_reg_1&_net_4);
   assign  _net_514 = (_reg_1&_net_4);
   assign  _net_515 = (_reg_1&_net_4);
   assign  _net_516 = (_reg_1&_net_4);
   assign  _net_517 = (_reg_1&_net_4);
   assign  _net_518 = (_reg_1&_net_4);
   assign  _net_519 = (_reg_1&_net_4);
   assign  _net_520 = (_reg_1&_net_4);
   assign  _net_521 = (_reg_1&_net_4);
   assign  _net_522 = (_reg_1&_net_4);
   assign  _net_523 = (_reg_1&_net_4);
   assign  _net_524 = (_reg_1&_net_4);
   assign  _net_525 = (_reg_1&_net_4);
   assign  _net_526 = (_reg_1&_net_4);
   assign  _net_527 = (_reg_1&_net_4);
   assign  _net_528 = (_reg_1&_net_4);
   assign  _net_529 = (_reg_1&_net_4);
   assign  _net_530 = (_reg_1&_net_4);
   assign  _net_531 = (_reg_1&_net_4);
   assign  _net_532 = (_reg_1&_net_4);
   assign  _net_533 = (_reg_1&_net_4);
   assign  _net_534 = (_reg_1&_net_4);
   assign  _net_535 = (_reg_1&_net_4);
   assign  _net_536 = (_reg_1&_net_4);
   assign  _net_537 = (_reg_1&_net_4);
   assign  _net_538 = (_reg_1&_net_4);
   assign  _net_539 = (_reg_1&_net_4);
   assign  _net_540 = (_reg_1&_net_4);
   assign  _net_541 = (_reg_1&_net_4);
   assign  _net_542 = (_reg_1&_net_4);
   assign  _net_543 = (_reg_1&_net_4);
   assign  _net_544 = (_reg_1&_net_4);
   assign  _net_545 = (_reg_1&_net_4);
   assign  _net_546 = (_reg_1&_net_4);
   assign  _net_547 = (_reg_1&_net_4);
   assign  _net_548 = (_reg_1&_net_4);
   assign  _net_549 = (_reg_1&_net_4);
   assign  _net_550 = (_reg_1&_net_4);
   assign  _net_551 = (_reg_1&_net_4);
   assign  _net_552 = (_reg_1&_net_4);
   assign  _net_553 = (_reg_1&_net_4);
   assign  _net_554 = (_reg_1&_net_4);
   assign  _net_555 = (_reg_1&_net_4);
   assign  _net_556 = (_reg_1&_net_4);
   assign  _net_557 = (_reg_1&_net_4);
   assign  _net_558 = (_reg_1&_net_4);
   assign  _net_559 = (_reg_1&_net_4);
   assign  _net_560 = (_reg_1&_net_4);
   assign  _net_561 = (_reg_1&_net_4);
   assign  _net_562 = (_reg_1&_net_4);
   assign  _net_563 = (_reg_1&_net_4);
   assign  _net_564 = (_reg_1&_net_4);
   assign  _net_565 = (_reg_1&_net_4);
   assign  _net_566 = (_reg_1&_net_4);
   assign  _net_567 = (_reg_1&_net_4);
   assign  _net_568 = (_reg_1&_net_4);
   assign  _net_569 = (_reg_1&_net_4);
   assign  _net_570 = (_reg_1&_net_4);
   assign  _net_571 = (_reg_1&_net_4);
   assign  _net_572 = (_reg_1&_net_4);
   assign  _net_573 = (_reg_1&_net_4);
   assign  _net_574 = (_reg_1&_net_4);
   assign  _net_575 = (_reg_1&_net_4);
   assign  _net_576 = (_reg_1&_net_4);
   assign  _net_577 = (_reg_1&_net_4);
   assign  _net_578 = (_reg_1&_net_4);
   assign  _net_579 = (_reg_1&_net_4);
   assign  _net_580 = (_reg_1&_net_4);
   assign  _net_581 = (_reg_1&_net_4);
   assign  _net_582 = (_reg_1&_net_4);
   assign  _net_583 = (_reg_1&_net_4);
   assign  _net_584 = (_reg_1&_net_4);
   assign  _net_585 = (_reg_1&_net_4);
   assign  _net_586 = (_reg_1&_net_4);
   assign  _net_587 = (_reg_1&_net_4);
   assign  _net_588 = (_reg_1&_net_4);
   assign  _net_589 = (_reg_1&_net_4);
   assign  _net_590 = (_reg_1&_net_4);
   assign  _net_591 = (_reg_1&_net_4);
   assign  _net_592 = (_reg_1&_net_4);
   assign  _net_593 = (_reg_1&_net_4);
   assign  _net_594 = (_reg_1&_net_4);
   assign  _net_595 = (_reg_1&_net_4);
   assign  _net_596 = (_reg_1&_net_4);
   assign  _net_597 = (_reg_1&_net_4);
   assign  _net_598 = (_reg_1&_net_4);
   assign  _net_599 = (_reg_1&_net_4);
   assign  _net_600 = (_reg_1&_net_4);
   assign  _net_601 = (_reg_1&_net_4);
   assign  _net_602 = (_reg_1&_net_4);
   assign  _net_603 = (_reg_1&_net_4);
   assign  _net_604 = (_reg_1&_net_4);
   assign  _net_605 = (_reg_1&_net_4);
   assign  _net_606 = (_reg_1&_net_4);
   assign  _net_607 = (_reg_1&_net_4);
   assign  _net_608 = (_reg_1&_net_4);
   assign  _net_609 = (_reg_1&_net_4);
   assign  _net_610 = (_reg_1&_net_4);
   assign  _net_611 = (_reg_1&_net_4);
   assign  _net_612 = (_reg_1&_net_4);
   assign  _net_613 = (_reg_1&_net_4);
   assign  _net_614 = (_reg_1&_net_4);
   assign  _net_615 = (_reg_1&_net_4);
   assign  _net_616 = (_reg_1&_net_4);
   assign  _net_617 = (_reg_1&_net_4);
   assign  _net_618 = (_reg_1&_net_4);
   assign  _net_619 = (_reg_1&_net_4);
   assign  _net_620 = (_reg_1&_net_4);
   assign  _net_621 = (_reg_1&_net_4);
   assign  _net_622 = (_reg_1&_net_4);
   assign  _net_623 = (_reg_1&_net_4);
   assign  _net_624 = (_reg_1&_net_4);
   assign  _net_625 = (_reg_1&_net_4);
   assign  _net_626 = (_reg_1&_net_4);
   assign  _net_627 = (_reg_1&_net_4);
   assign  _net_628 = (_reg_1&_net_4);
   assign  _net_629 = (_reg_1&_net_4);
   assign  _net_630 = (_reg_1&_net_4);
   assign  _net_631 = (_reg_1&_net_4);
   assign  _net_632 = (_reg_1&_net_4);
   assign  _net_633 = (_reg_1&_net_4);
   assign  _net_634 = (_reg_1&_net_4);
   assign  _net_635 = (_reg_1&_net_4);
   assign  _net_636 = (_reg_1&_net_4);
   assign  _net_637 = (_reg_1&_net_4);
   assign  _net_638 = (_reg_1&_net_4);
   assign  _net_639 = (_reg_1&_net_4);
   assign  _net_640 = (_reg_1&_net_4);
   assign  _net_641 = (_reg_1&_net_4);
   assign  _net_642 = (_reg_1&_net_4);
   assign  _net_643 = (_reg_1&_net_4);
   assign  _net_644 = (_reg_1&_net_4);
   assign  _net_645 = (_reg_1&_net_4);
   assign  _net_646 = (_reg_1&_net_4);
   assign  _net_647 = (_reg_1&_net_4);
   assign  _net_648 = (_reg_1&_net_4);
   assign  _net_649 = (_reg_1&_net_4);
   assign  _net_650 = (_reg_1&_net_4);
   assign  _net_651 = (_reg_1&_net_4);
   assign  _net_652 = (_reg_1&_net_4);
   assign  _net_653 = (_reg_1&_net_4);
   assign  _net_654 = (_reg_1&_net_4);
   assign  _net_655 = (_reg_1&_net_4);
   assign  _net_656 = (_reg_1&_net_4);
   assign  _net_657 = (_reg_1&_net_4);
   assign  _net_658 = (_reg_1&_net_4);
   assign  _net_659 = (_reg_1&_net_4);
   assign  _net_660 = (_reg_1&_net_4);
   assign  _net_661 = (_reg_1&_net_4);
   assign  _net_662 = (_reg_1&_net_4);
   assign  _net_663 = (_reg_1&_net_4);
   assign  _net_664 = (_reg_1&_net_4);
   assign  _net_665 = (_reg_1&_net_4);
   assign  _net_666 = (_reg_1&_net_4);
   assign  _net_667 = (_reg_1&_net_4);
   assign  _net_668 = (_reg_1&_net_4);
   assign  _net_669 = (_reg_1&_net_4);
   assign  _net_670 = (_reg_1&_net_4);
   assign  _net_671 = (_reg_1&_net_4);
   assign  _net_672 = (_reg_1&_net_4);
   assign  _net_673 = (_reg_1&_net_4);
   assign  _net_674 = (_reg_1&_net_4);
   assign  _net_675 = (_reg_1&_net_4);
   assign  _net_676 = (_reg_1&_net_4);
   assign  _net_677 = (_reg_1&_net_4);
   assign  _net_678 = (_reg_1&_net_4);
   assign  _net_679 = (_reg_1&_net_4);
   assign  _net_680 = (_reg_1&_net_4);
   assign  _net_681 = (_reg_1&_net_4);
   assign  _net_682 = (_reg_1&_net_4);
   assign  _net_683 = (_reg_1&_net_4);
   assign  _net_684 = (_reg_1&_net_4);
   assign  _net_685 = (_reg_1&_net_4);
   assign  _net_686 = (_reg_1&_net_4);
   assign  _net_687 = (_reg_1&_net_4);
   assign  _net_688 = (_reg_1&_net_4);
   assign  _net_689 = (_reg_1&_net_4);
   assign  _net_690 = (_reg_1&_net_4);
   assign  _net_691 = (_reg_1&_net_4);
   assign  _net_692 = (_reg_1&_net_4);
   assign  _net_693 = (_reg_1&_net_4);
   assign  _net_694 = (_reg_1&_net_4);
   assign  _net_695 = (_reg_1&_net_4);
   assign  _net_696 = (_reg_1&_net_4);
   assign  _net_697 = (_reg_1&_net_4);
   assign  _net_698 = (_reg_1&_net_4);
   assign  _net_699 = (_reg_1&_net_4);
   assign  _net_700 = (_reg_1&_net_4);
   assign  _net_701 = (_reg_1&_net_4);
   assign  _net_702 = (_reg_1&_net_4);
   assign  _net_703 = (_reg_1&_net_4);
   assign  _net_704 = (_reg_1&_net_4);
   assign  _net_705 = (_reg_1&_net_4);
   assign  _net_706 = (_reg_1&_net_4);
   assign  _net_707 = (_reg_1&_net_4);
   assign  _net_708 = (_reg_1&_net_4);
   assign  _net_709 = (_reg_1&_net_4);
   assign  _net_710 = (_reg_1&_net_4);
   assign  _net_711 = (_reg_1&_net_4);
   assign  _net_712 = (_reg_1&_net_4);
   assign  _net_713 = (_reg_1&_net_4);
   assign  _net_714 = (_reg_1&_net_4);
   assign  _net_715 = (_reg_1&_net_4);
   assign  _net_716 = (_reg_1&_net_4);
   assign  _net_717 = (_reg_1&_net_4);
   assign  _net_718 = (_reg_1&_net_4);
   assign  _net_719 = (_reg_1&_net_4);
   assign  _net_720 = (_reg_1&_net_4);
   assign  _net_721 = (_reg_1&_net_4);
   assign  _net_722 = (_reg_1&_net_4);
   assign  _net_723 = (_reg_1&_net_4);
   assign  _net_724 = (_reg_1&_net_4);
   assign  _net_725 = (_reg_1&_net_4);
   assign  _net_726 = (_reg_1&_net_4);
   assign  _net_727 = (_reg_1&_net_4);
   assign  _net_728 = (_reg_1&_net_4);
   assign  _net_729 = (_reg_1&_net_4);
   assign  _net_730 = (_reg_1&_net_4);
   assign  _net_731 = (_reg_1&_net_4);
   assign  _net_732 = (_reg_1&_net_4);
   assign  _net_733 = (_reg_1&_net_4);
   assign  _net_734 = (_reg_1&_net_4);
   assign  _net_735 = (_reg_1&_net_4);
   assign  _net_736 = (_reg_1&_net_4);
   assign  _net_737 = (_reg_1&_net_4);
   assign  _net_738 = (_reg_1&_net_4);
   assign  _net_739 = (_reg_1&_net_4);
   assign  _net_740 = (_reg_1&_net_4);
   assign  _net_741 = (_reg_1&_net_4);
   assign  _net_742 = (_reg_1&_net_4);
   assign  _net_743 = (_reg_1&_net_4);
   assign  _net_744 = (_reg_1&_net_4);
   assign  _net_745 = (_reg_1&_net_4);
   assign  _net_746 = (_reg_1&_net_4);
   assign  _net_747 = (_reg_1&_net_4);
   assign  _net_748 = (_reg_1&_net_4);
   assign  _net_749 = (_reg_1&_net_4);
   assign  _net_750 = (_reg_1&_net_4);
   assign  _net_751 = (_reg_1&_net_4);
   assign  _net_752 = (_reg_1&_net_4);
   assign  _net_753 = (_reg_1&_net_4);
   assign  _net_754 = (_reg_1&_net_4);
   assign  _net_755 = (_reg_1&_net_4);
   assign  _net_756 = (_reg_1&_net_4);
   assign  _net_757 = (_reg_1&_net_4);
   assign  _net_758 = (_reg_1&_net_4);
   assign  _net_759 = (_reg_1&_net_4);
   assign  _net_760 = (_reg_1&_net_4);
   assign  _net_761 = (_reg_1&_net_4);
   assign  _net_762 = (_reg_1&_net_4);
   assign  _net_763 = (_reg_1&_net_4);
   assign  _net_764 = (_reg_1&_net_4);
   assign  _net_765 = (_reg_1&_net_4);
   assign  _net_766 = (_reg_1&_net_4);
   assign  _net_767 = (_reg_1&_net_4);
   assign  _net_768 = (_reg_1&_net_4);
   assign  _net_769 = (_reg_1&_net_4);
   assign  _net_770 = (_reg_1&_net_4);
   assign  _net_771 = (_reg_1&_net_4);
   assign  _net_772 = (_reg_1&_net_4);
   assign  _net_773 = (_reg_1&_net_4);
   assign  _net_774 = (_reg_1&_net_4);
   assign  _net_775 = (_reg_1&_net_4);
   assign  _net_776 = (_reg_1&_net_4);
   assign  _net_777 = (_reg_1&_net_4);
   assign  _net_778 = (_reg_1&_net_4);
   assign  _net_779 = (_reg_1&_net_4);
   assign  _net_780 = (_reg_1&_net_4);
   assign  _net_781 = (_reg_1&_net_4);
   assign  _net_782 = (_reg_1&_net_4);
   assign  _net_783 = (_reg_1&_net_4);
   assign  _net_784 = (_reg_1&_net_4);
   assign  _net_785 = (_reg_1&_net_4);
   assign  _net_786 = (_reg_1&_net_4);
   assign  _net_787 = (_reg_1&_net_4);
   assign  _net_788 = (_reg_1&_net_4);
   assign  _net_789 = (_reg_1&_net_4);
   assign  _net_790 = (_reg_1&_net_4);
   assign  _net_791 = (_reg_1&_net_4);
   assign  _net_792 = (_reg_1&_net_4);
   assign  _net_793 = (_reg_1&_net_4);
   assign  _net_794 = (_reg_1&_net_4);
   assign  _net_795 = (_reg_1&_net_4);
   assign  _net_796 = (_reg_1&_net_4);
   assign  _net_797 = (_reg_1&_net_4);
   assign  _net_798 = (_reg_1&_net_4);
   assign  _net_799 = (_reg_1&_net_4);
   assign  _net_800 = (_reg_1&_net_4);
   assign  _net_801 = (_reg_1&_net_4);
   assign  _net_802 = (_reg_1&_net_4);
   assign  _net_803 = (_reg_1&_net_4);
   assign  _net_804 = (_reg_1&_net_4);
   assign  _net_805 = (_reg_1&_net_4);
   assign  _net_806 = (_reg_1&_net_4);
   assign  _net_807 = (_reg_1&_net_4);
   assign  _net_808 = (_reg_1&_net_4);
   assign  _net_809 = (_reg_1&_net_4);
   assign  _net_810 = (_reg_1&_net_4);
   assign  _net_811 = (_reg_1&_net_4);
   assign  _net_812 = (_reg_1&_net_4);
   assign  _net_813 = (_reg_1&_net_4);
   assign  _net_814 = (_reg_1&_net_4);
   assign  _net_815 = (_reg_1&_net_4);
   assign  _net_816 = (_reg_1&_net_4);
   assign  _net_817 = (_reg_1&_net_4);
   assign  _net_818 = (_reg_1&_net_4);
   assign  _net_819 = (_reg_1&_net_4);
   assign  _net_820 = (_reg_1&_net_4);
   assign  _net_821 = (_reg_1&_net_4);
   assign  _net_822 = (_reg_1&_net_4);
   assign  _net_823 = (_reg_1&_net_4);
   assign  _net_824 = (_reg_1&_net_4);
   assign  _net_825 = (_reg_1&_net_4);
   assign  _net_826 = (_reg_1&_net_4);
   assign  _net_827 = (_reg_1&_net_4);
   assign  _net_828 = (_reg_1&_net_4);
   assign  _net_829 = (_reg_1&_net_4);
   assign  _net_830 = (_reg_1&_net_4);
   assign  _net_831 = (_reg_1&_net_4);
   assign  _net_832 = (_reg_1&_net_4);
   assign  _net_833 = (_reg_1&_net_4);
   assign  _net_834 = (_reg_1&_net_4);
   assign  _net_835 = (_reg_1&_net_4);
   assign  _net_836 = (_reg_1&_net_4);
   assign  _net_837 = (_reg_1&_net_4);
   assign  _net_838 = (_reg_1&_net_4);
   assign  _net_839 = (_reg_1&_net_4);
   assign  _net_840 = (_reg_1&_net_4);
   assign  _net_841 = (_reg_1&_net_4);
   assign  _net_842 = (_reg_1&_net_4);
   assign  _net_843 = (_reg_1&_net_4);
   assign  _net_844 = (_reg_1&_net_4);
   assign  _net_845 = (_reg_1&_net_4);
   assign  _net_846 = (_reg_1&_net_4);
   assign  _net_847 = (_reg_1&_net_4);
   assign  _net_848 = (_reg_1&_net_4);
   assign  _net_849 = (_reg_1&_net_4);
   assign  _net_850 = (_reg_1&_net_4);
   assign  _net_851 = (_reg_1&_net_4);
   assign  _net_852 = (_reg_1&_net_4);
   assign  _net_853 = (_reg_1&_net_4);
   assign  _net_854 = (_reg_1&_net_4);
   assign  _net_855 = (_reg_1&_net_4);
   assign  _net_856 = (_reg_1&_net_4);
   assign  _net_857 = (_reg_1&_net_4);
   assign  _net_858 = (_reg_1&_net_4);
   assign  _net_859 = (_reg_1&_net_4);
   assign  _net_860 = (_reg_1&_net_4);
   assign  _net_861 = (_reg_1&_net_4);
   assign  _net_862 = (_reg_1&_net_4);
   assign  _net_863 = (_reg_1&_net_4);
   assign  _net_864 = (_reg_1&_net_4);
   assign  _net_865 = (_reg_1&_net_4);
   assign  _net_866 = (_reg_1&_net_4);
   assign  _net_867 = (_reg_1&_net_4);
   assign  _net_868 = (_reg_1&_net_4);
   assign  _net_869 = (_reg_1&_net_4);
   assign  _net_870 = (_reg_1&_net_4);
   assign  _net_871 = (_reg_1&_net_4);
   assign  _net_872 = (_reg_1&_net_4);
   assign  _net_873 = (_reg_1&_net_4);
   assign  _net_874 = (_reg_1&_net_4);
   assign  _net_875 = (_reg_1&_net_4);
   assign  _net_876 = (_reg_1&_net_4);
   assign  _net_877 = (_reg_1&_net_4);
   assign  _net_878 = (_reg_1&_net_4);
   assign  _net_879 = (_reg_1&_net_4);
   assign  _net_880 = (_reg_1&_net_4);
   assign  _net_881 = (_reg_1&_net_4);
   assign  _net_882 = (_reg_1&_net_4);
   assign  _net_883 = (_reg_1&_net_4);
   assign  _net_884 = (_reg_1&_net_4);
   assign  _net_885 = (_reg_1&_net_4);
   assign  _net_886 = (_reg_1&_net_4);
   assign  _net_887 = (_reg_1&_net_4);
   assign  _net_888 = (_reg_1&_net_4);
   assign  _net_889 = (_reg_1&_net_4);
   assign  _net_890 = (_reg_1&_net_4);
   assign  _net_891 = (_reg_1&_net_4);
   assign  _net_892 = (_reg_1&_net_4);
   assign  _net_893 = (_reg_1&_net_4);
   assign  _net_894 = (_reg_1&_net_4);
   assign  _net_895 = (_reg_1&_net_4);
   assign  _net_896 = (_reg_1&_net_4);
   assign  _net_897 = (_reg_1&_net_4);
   assign  _net_898 = (_reg_1&_net_4);
   assign  _net_899 = (_reg_1&_net_4);
   assign  _net_900 = (_reg_1&_net_4);
   assign  _net_901 = (_reg_1&_net_4);
   assign  _net_902 = (_reg_1&_net_4);
   assign  _net_903 = (_reg_1&_net_4);
   assign  _net_904 = (_reg_1&_net_4);
   assign  _net_905 = (_reg_1&_net_4);
   assign  _net_906 = (_reg_1&_net_4);
   assign  _net_907 = (_reg_1&_net_4);
   assign  _net_908 = (_reg_1&_net_4);
   assign  _net_909 = (_reg_1&_net_4);
   assign  _net_910 = (_reg_1&_net_4);
   assign  _net_911 = (_reg_1&_net_4);
   assign  _net_912 = (_reg_1&_net_4);
   assign  _net_913 = (_reg_1&_net_4);
   assign  _net_914 = (_reg_1&_net_4);
   assign  _net_915 = (_reg_1&_net_4);
   assign  _net_916 = (_reg_1&_net_4);
   assign  _net_917 = (_reg_1&_net_4);
   assign  _net_918 = (_reg_1&_net_4);
   assign  _net_919 = (_reg_1&_net_4);
   assign  _net_920 = (_reg_1&_net_4);
   assign  _net_921 = (_reg_1&_net_4);
   assign  _net_922 = (_reg_1&_net_4);
   assign  _net_923 = (_reg_1&_net_4);
   assign  _net_924 = (_reg_1&_net_4);
   assign  _net_925 = (_reg_1&_net_4);
   assign  _net_926 = (_reg_1&_net_4);
   assign  _net_927 = (_reg_1&_net_4);
   assign  _net_928 = (_reg_1&_net_4);
   assign  _net_929 = (_reg_1&_net_4);
   assign  _net_930 = (_reg_1&_net_4);
   assign  _net_931 = (_reg_1&_net_4);
   assign  _net_932 = (_reg_1&_net_4);
   assign  _net_933 = (_reg_1&_net_4);
   assign  _net_934 = (_reg_1&_net_4);
   assign  _net_935 = (_reg_1&_net_4);
   assign  _net_936 = (_reg_1&_net_4);
   assign  _net_937 = (_reg_1&_net_4);
   assign  _net_938 = (_reg_1&_net_4);
   assign  _net_939 = (_reg_1&_net_4);
   assign  _net_940 = (_reg_1&_net_4);
   assign  _net_941 = (_reg_1&_net_4);
   assign  _net_942 = (_reg_1&_net_4);
   assign  _net_943 = (_reg_1&_net_4);
   assign  _net_944 = (_reg_1&_net_4);
   assign  _net_945 = (_reg_1&_net_4);
   assign  _net_946 = (_reg_1&_net_4);
   assign  _net_947 = (_reg_1&_net_4);
   assign  _net_948 = (_reg_1&_net_4);
   assign  _net_949 = (_reg_1&_net_4);
   assign  _net_950 = (_reg_1&_net_4);
   assign  _net_951 = (_reg_1&_net_4);
   assign  _net_952 = (_reg_1&_net_4);
   assign  _net_953 = (_reg_1&_net_4);
   assign  _net_954 = (_reg_1&_net_4);
   assign  _net_955 = (_reg_1&_net_4);
   assign  _net_956 = (_reg_1&_net_4);
   assign  _net_957 = (_reg_1&_net_4);
   assign  _net_958 = (_reg_1&_net_4);
   assign  _net_959 = (_reg_1&_net_4);
   assign  _net_960 = (_reg_1&_net_4);
   assign  _net_961 = (_reg_1&_net_4);
   assign  _net_962 = (_reg_1&_net_4);
   assign  _net_963 = (_reg_1&_net_4);
   assign  _net_964 = (_reg_1&_net_4);
   assign  _net_965 = (_reg_1&_net_4);
   assign  _net_966 = (_reg_1&_net_4);
   assign  _net_967 = (_reg_1&_net_4);
   assign  _net_968 = (_reg_1&_net_4);
   assign  _net_969 = (_reg_1&_net_4);
   assign  _net_970 = (_reg_1&_net_4);
   assign  _net_971 = (_reg_1&_net_4);
   assign  _net_972 = (_reg_1&_net_4);
   assign  _net_973 = (_reg_1&_net_4);
   assign  _net_974 = (_reg_1&_net_4);
   assign  _net_975 = (_reg_1&_net_4);
   assign  _net_976 = (_reg_1&_net_4);
   assign  _net_977 = (_reg_1&_net_4);
   assign  _net_978 = (_reg_1&_net_4);
   assign  _net_979 = (_reg_1&_net_4);
   assign  _net_980 = (_reg_1&_net_4);
   assign  _net_981 = (_reg_1&_net_4);
   assign  _net_982 = (_reg_1&_net_4);
   assign  _net_983 = (_reg_1&_net_4);
   assign  _net_984 = (_reg_1&_net_4);
   assign  _net_985 = (_reg_1&_net_4);
   assign  _net_986 = (_reg_1&_net_4);
   assign  _net_987 = (_reg_1&_net_4);
   assign  _net_988 = (_reg_1&_net_4);
   assign  _net_989 = (_reg_1&_net_4);
   assign  _net_990 = (_reg_1&_net_4);
   assign  _net_991 = (_reg_1&_net_4);
   assign  _net_992 = (_reg_1&_net_4);
   assign  _net_993 = (_reg_1&_net_4);
   assign  _net_994 = (_reg_1&_net_4);
   assign  _net_995 = (_reg_1&_net_4);
   assign  _net_996 = (_reg_1&_net_4);
   assign  _net_997 = (_reg_1&_net_4);
   assign  _net_998 = (_reg_1&_net_4);
   assign  _net_999 = (_reg_1&_net_4);
   assign  _net_1000 = (_reg_1&_net_4);
   assign  _net_1001 = (_reg_1&_net_4);
   assign  _net_1002 = (_reg_1&_net_4);
   assign  _net_1003 = (_reg_1&_net_4);
   assign  _net_1004 = (_reg_1&_net_4);
   assign  _net_1005 = (_reg_1&_net_4);
   assign  _net_1006 = (_reg_1&_net_4);
   assign  _net_1007 = (_reg_1&_net_4);
   assign  _net_1008 = (_reg_1&_net_4);
   assign  _net_1009 = (_reg_1&_net_4);
   assign  _net_1010 = (_reg_1&_net_4);
   assign  _net_1011 = (_reg_1&_net_4);
   assign  _net_1012 = (_reg_1&_net_4);
   assign  _net_1013 = (_reg_1&_net_4);
   assign  _net_1014 = (_reg_1&_net_4);
   assign  _net_1015 = (_reg_1&_net_4);
   assign  _net_1016 = (_reg_1&_net_4);
   assign  _net_1017 = (_reg_1&_net_4);
   assign  _net_1018 = (_reg_1&_net_4);
   assign  _net_1019 = (_reg_1&_net_4);
   assign  _net_1020 = (_reg_1&_net_4);
   assign  _net_1021 = (_reg_1&_net_4);
   assign  _net_1022 = (_reg_1&_net_4);
   assign  _net_1023 = (_reg_1&_net_4);
   assign  _net_1024 = (_reg_1&_net_4);
   assign  _net_1025 = (_reg_1&_net_4);
   assign  _net_1026 = (_reg_1&_net_4);
   assign  _net_1027 = (_reg_1&_net_4);
   assign  _net_1028 = (_reg_1&_net_4);
   assign  _net_1029 = (_reg_1&_net_4);
   assign  _net_1030 = (_reg_1&_net_4);
   assign  _net_1031 = (_reg_1&_net_4);
   assign  _net_1032 = (_reg_1&_net_4);
   assign  _net_1033 = (_reg_1&_net_4);
   assign  _net_1034 = (_reg_1&_net_4);
   assign  _net_1035 = (_reg_1&_net_4);
   assign  _net_1036 = (_reg_1&_net_4);
   assign  _net_1037 = (_reg_1&_net_4);
   assign  _net_1038 = (_reg_1&_net_4);
   assign  _net_1039 = (_reg_1&_net_4);
   assign  _net_1040 = (_reg_1&_net_4);
   assign  _net_1041 = (_reg_1&_net_4);
   assign  _net_1042 = (_reg_1&_net_4);
   assign  _net_1043 = (_reg_1&_net_4);
   assign  _net_1044 = (_reg_1&_net_4);
   assign  _net_1045 = (_reg_1&_net_4);
   assign  _net_1046 = (_reg_1&_net_4);
   assign  _net_1047 = (_reg_1&_net_4);
   assign  _net_1048 = (_reg_1&_net_4);
   assign  _net_1049 = (_reg_1&_net_4);
   assign  _net_1050 = (_reg_1&_net_4);
   assign  _net_1051 = (_reg_1&_net_4);
   assign  _net_1052 = (_reg_1&_net_4);
   assign  _net_1053 = (_reg_1&_net_4);
   assign  _net_1054 = (_reg_1&_net_4);
   assign  _net_1055 = (_reg_1&_net_4);
   assign  _net_1056 = (_reg_1&_net_4);
   assign  _net_1057 = (_reg_1&_net_4);
   assign  _net_1058 = (_reg_1&_net_4);
   assign  _net_1059 = (_reg_1&_net_4);
   assign  _net_1060 = (_reg_1&_net_4);
   assign  _net_1061 = (_reg_1&_net_4);
   assign  _net_1062 = (_reg_1&_net_4);
   assign  _net_1063 = (_reg_1&_net_4);
   assign  _net_1064 = (_reg_1&_net_4);
   assign  _net_1065 = (_reg_1&_net_4);
   assign  _net_1066 = (_reg_1&_net_4);
   assign  _net_1067 = (_reg_1&_net_4);
   assign  _net_1068 = (_reg_1&_net_4);
   assign  _net_1069 = (_reg_1&_net_4);
   assign  _net_1070 = (_reg_1&_net_4);
   assign  _net_1071 = (_reg_1&_net_4);
   assign  _net_1072 = (_reg_1&_net_4);
   assign  _net_1073 = (_reg_1&_net_4);
   assign  _net_1074 = (_reg_1&_net_4);
   assign  _net_1075 = (_reg_1&_net_4);
   assign  _net_1076 = (_reg_1&_net_4);
   assign  _net_1077 = (_reg_1&_net_4);
   assign  _net_1078 = (_reg_1&_net_4);
   assign  _net_1079 = (_reg_1&_net_4);
   assign  _net_1080 = (_reg_1&_net_4);
   assign  _net_1081 = (_reg_1&_net_4);
   assign  _net_1082 = (_reg_1&_net_4);
   assign  _net_1083 = (_reg_1&_net_4);
   assign  _net_1084 = (_reg_1&_net_4);
   assign  _net_1085 = (_reg_1&_net_4);
   assign  _net_1086 = (_reg_1&_net_4);
   assign  _net_1087 = (_reg_1&_net_4);
   assign  _net_1088 = (_reg_1&_net_4);
   assign  _net_1089 = (_reg_1&_net_4);
   assign  _net_1090 = (_reg_1&_net_4);
   assign  _net_1091 = (_reg_1&_net_4);
   assign  _net_1092 = (_reg_1&_net_4);
   assign  _net_1093 = (_reg_1&_net_4);
   assign  _net_1094 = (_reg_1&_net_4);
   assign  _net_1095 = (_reg_1&_net_4);
   assign  _net_1096 = (_reg_1&_net_4);
   assign  _net_1097 = (_reg_1&_net_4);
   assign  _net_1098 = (_reg_1&_net_4);
   assign  _net_1099 = (_reg_1&_net_4);
   assign  _net_1100 = (_reg_1&_net_4);
   assign  _net_1101 = (_reg_1&_net_4);
   assign  _net_1102 = (_reg_1&_net_4);
   assign  _net_1103 = (_reg_1&_net_4);
   assign  _net_1104 = (_reg_1&_net_4);
   assign  _net_1105 = (_reg_1&_net_4);
   assign  _net_1106 = (_reg_1&_net_4);
   assign  _net_1107 = (_reg_1&_net_4);
   assign  _net_1108 = (_reg_1&_net_4);
   assign  _net_1109 = (_reg_1&_net_4);
   assign  _net_1110 = (_reg_1&_net_4);
   assign  _net_1111 = (_reg_1&_net_4);
   assign  _net_1112 = (_reg_1&_net_4);
   assign  _net_1113 = (_reg_1&_net_4);
   assign  _net_1114 = (_reg_1&_net_4);
   assign  _net_1115 = (_reg_1&_net_4);
   assign  _net_1116 = (_reg_1&_net_4);
   assign  _net_1117 = (_reg_1&_net_4);
   assign  _net_1118 = (_reg_1&_net_4);
   assign  _net_1119 = (_reg_1&_net_4);
   assign  _net_1120 = (_reg_1&_net_4);
   assign  _net_1121 = (_reg_1&_net_4);
   assign  _net_1122 = (_reg_1&_net_4);
   assign  _net_1123 = (_reg_1&_net_4);
   assign  _net_1124 = (_reg_1&_net_4);
   assign  _net_1125 = (_reg_1&_net_4);
   assign  _net_1126 = (_reg_1&_net_4);
   assign  _net_1127 = (_reg_1&_net_4);
   assign  _net_1128 = (_reg_1&_net_4);
   assign  _net_1129 = (_reg_1&_net_4);
   assign  _net_1130 = (_reg_1&_net_4);
   assign  _net_1131 = (_reg_1&_net_4);
   assign  _net_1132 = (_reg_1&_net_4);
   assign  _net_1133 = (_reg_1&_net_4);
   assign  _net_1134 = (_reg_1&_net_4);
   assign  _net_1135 = (_reg_1&_net_4);
   assign  _net_1136 = (_reg_1&_net_4);
   assign  _net_1137 = (_reg_1&_net_4);
   assign  _net_1138 = (_reg_1&_net_4);
   assign  _net_1139 = (_reg_1&_net_4);
   assign  _net_1140 = (_reg_1&_net_4);
   assign  _net_1141 = (_reg_1&_net_4);
   assign  _net_1142 = (_reg_1&_net_4);
   assign  _net_1143 = (_reg_1&_net_4);
   assign  _net_1144 = (_reg_1&_net_4);
   assign  _net_1145 = (_reg_1&_net_4);
   assign  _net_1146 = (_reg_1&_net_4);
   assign  _net_1147 = (_reg_1&_net_4);
   assign  _net_1148 = (_reg_1&_net_4);
   assign  _net_1149 = (_reg_1&_net_4);
   assign  _net_1150 = (_reg_1&_net_4);
   assign  _net_1151 = (_reg_1&_net_4);
   assign  _net_1152 = (_reg_1&_net_4);
   assign  _net_1153 = (_reg_1&_net_4);
   assign  _net_1154 = (_reg_1&_net_4);
   assign  _net_1155 = (_reg_1&_net_4);
   assign  _net_1156 = (_reg_1&_net_4);
   assign  _net_1157 = (_reg_1&_net_4);
   assign  _net_1158 = (_reg_1&_net_4);
   assign  _net_1159 = (_reg_1&_net_4);
   assign  _net_1160 = (_reg_1&_net_4);
   assign  _net_1161 = (_reg_1&_net_4);
   assign  _net_1162 = (_reg_1&_net_4);
   assign  _net_1163 = (_reg_1&_net_4);
   assign  _net_1164 = (_reg_1&_net_4);
   assign  _net_1165 = (_reg_1&_net_4);
   assign  _net_1166 = (_reg_1&_net_4);
   assign  _net_1167 = (_reg_1&_net_4);
   assign  _net_1168 = (_reg_1&_net_4);
   assign  _net_1169 = (_reg_1&_net_4);
   assign  _net_1170 = (_reg_1&_net_4);
   assign  _net_1171 = (_reg_1&_net_4);
   assign  _net_1172 = (_reg_1&_net_4);
   assign  _net_1173 = (_reg_1&_net_4);
   assign  _net_1174 = (_reg_1&_net_4);
   assign  _net_1175 = (_reg_1&_net_4);
   assign  _net_1176 = (_reg_1&_net_4);
   assign  _net_1177 = (_reg_1&_net_4);
   assign  _net_1178 = (_reg_1&_net_4);
   assign  _net_1179 = (_reg_1&_net_4);
   assign  _net_1180 = (_reg_1&_net_4);
   assign  _net_1181 = (_reg_1&_net_4);
   assign  _net_1182 = (_reg_1&_net_4);
   assign  _net_1183 = (_reg_1&_net_4);
   assign  _net_1184 = (_reg_1&_net_4);
   assign  _net_1185 = (_reg_1&_net_4);
   assign  _net_1186 = (_reg_1&_net_4);
   assign  _net_1187 = (_reg_1&_net_4);
   assign  _net_1188 = (_reg_1&_net_4);
   assign  _net_1189 = (_reg_1&_net_4);
   assign  _net_1190 = (_reg_1&_net_4);
   assign  _net_1191 = (_reg_1&_net_4);
   assign  _net_1192 = (_reg_1&_net_4);
   assign  _net_1193 = (_reg_1&_net_4);
   assign  _net_1194 = (_reg_1&_net_4);
   assign  _net_1195 = (_reg_1&_net_4);
   assign  _net_1196 = (_reg_1&_net_4);
   assign  _net_1197 = (_reg_1&_net_4);
   assign  _net_1198 = (_reg_1&_net_4);
   assign  _net_1199 = (_reg_1&_net_4);
   assign  _net_1200 = (_reg_1&_net_4);
   assign  _net_1201 = (_reg_1&_net_4);
   assign  _net_1202 = (_reg_1&_net_4);
   assign  _net_1203 = (_reg_1&_net_4);
   assign  _net_1204 = (_reg_1&_net_4);
   assign  _net_1205 = (_reg_1&_net_4);
   assign  _net_1206 = (_reg_1&_net_4);
   assign  _net_1207 = (_reg_1&_net_4);
   assign  _net_1208 = (_reg_1&_net_4);
   assign  _net_1209 = (_reg_1&_net_4);
   assign  _net_1210 = (_reg_1&_net_4);
   assign  _net_1211 = (_reg_1&_net_4);
   assign  _net_1212 = (_reg_1&_net_4);
   assign  _net_1213 = (_reg_1&_net_4);
   assign  _net_1214 = (_reg_1&_net_4);
   assign  _net_1215 = (_reg_1&_net_4);
   assign  _net_1216 = (_reg_1&_net_4);
   assign  _net_1217 = (_reg_1&_net_4);
   assign  _net_1218 = (_reg_1&_net_4);
   assign  _net_1219 = (_reg_1&_net_4);
   assign  _net_1220 = (_reg_1&_net_4);
   assign  _net_1221 = (_reg_1&_net_4);
   assign  _net_1222 = (_reg_1&_net_4);
   assign  _net_1223 = (_reg_1&_net_4);
   assign  _net_1224 = (_reg_1&_net_4);
   assign  _net_1225 = (_reg_1&_net_4);
   assign  _net_1226 = (_reg_1&_net_4);
   assign  _net_1227 = (_reg_1&_net_4);
   assign  _net_1228 = (_reg_1&_net_4);
   assign  _net_1229 = (_reg_1&_net_4);
   assign  _net_1230 = (_reg_1&_net_4);
   assign  _net_1231 = (_reg_1&_net_4);
   assign  _net_1232 = (_reg_1&_net_4);
   assign  _net_1233 = (_reg_1&_net_4);
   assign  _net_1234 = (_reg_1&_net_4);
   assign  _net_1235 = (_reg_1&_net_4);
   assign  _net_1236 = (_reg_1&_net_4);
   assign  _net_1237 = (_reg_1&_net_4);
   assign  _net_1238 = (_reg_1&_net_4);
   assign  _net_1239 = (_reg_1&_net_4);
   assign  _net_1240 = (_reg_1&_net_4);
   assign  _net_1241 = (_reg_1&_net_4);
   assign  _net_1242 = (_reg_1&_net_4);
   assign  _net_1243 = (_reg_1&_net_4);
   assign  _net_1244 = (_reg_1&_net_4);
   assign  _net_1245 = (_reg_1&_net_4);
   assign  _net_1246 = (_reg_1&_net_4);
   assign  _net_1247 = (_reg_1&_net_4);
   assign  _net_1248 = (_reg_1&_net_4);
   assign  _net_1249 = (_reg_1&_net_4);
   assign  _net_1250 = (_reg_1&_net_4);
   assign  _net_1251 = (_reg_1&_net_4);
   assign  _net_1252 = (_reg_1&_net_4);
   assign  _net_1253 = (_reg_1&_net_4);
   assign  _net_1254 = (_reg_1&_net_4);
   assign  _net_1255 = (_reg_1&_net_4);
   assign  _net_1256 = (_reg_1&_net_4);
   assign  _net_1257 = (_reg_1&_net_4);
   assign  _net_1258 = (_reg_1&_net_4);
   assign  _net_1259 = (_reg_1&_net_4);
   assign  _net_1260 = (_reg_1&_net_4);
   assign  _net_1261 = (_reg_1&_net_4);
   assign  _net_1262 = (_reg_1&_net_4);
   assign  _net_1263 = (_reg_1&_net_4);
   assign  _net_1264 = (_reg_1&_net_4);
   assign  _net_1265 = (_reg_1&_net_4);
   assign  _net_1266 = (_reg_1&_net_4);
   assign  _net_1267 = (_reg_1&_net_4);
   assign  _net_1268 = (_reg_1&_net_4);
   assign  _net_1269 = (_reg_1&_net_4);

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_net_1271)
    begin
    $display("exit %b",kanwa_exit);
    end
  end

// synthesis translate_on
// synopsys translate_on
   assign  _net_1271 = (_reg_1&_net_4);
   assign  _reg_1_goto = _net_1272;
   assign  _net_1272 = (_reg_1&_net_4);
   assign  _reg_2_goin = _net_1273;
   assign  _net_1273 = (_reg_1&_net_4);

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_reg_2)
    begin
    $display("exit %b,dig_exit%d",kanwa_exit,dig_exit);
    end
  end

// synthesis translate_on
// synopsys translate_on
   assign  _net_1275 = (in_do|_reg_3);
   assign  _net_1276 = (in_do|_reg_3);
   assign  _net_1277 = (in_do|_reg_3);
   assign  _net_1278 = (in_do|_reg_3);
   assign  _net_1279 = (in_do|_reg_3);
   assign  _net_1280 = (in_do|_reg_3);
   assign  _net_1281 = (in_do|_reg_3);
   assign  _net_1282 = (in_do|_reg_3);
   assign  _net_1283 = (in_do|_reg_3);
   assign  _net_1284 = (in_do|_reg_3);
   assign  _net_1285 = (in_do|_reg_3);
   assign  _net_1286 = (in_do|_reg_3);
   assign  _net_1287 = (in_do|_reg_3);
   assign  _net_1288 = (in_do|_reg_3);
   assign  _net_1289 = (in_do|_reg_3);
   assign  _net_1290 = (in_do|_reg_3);
   assign  _net_1291 = (in_do|_reg_3);
   assign  _net_1292 = (in_do|_reg_3);
   assign  _net_1293 = (in_do|_reg_3);
   assign  _net_1294 = (in_do|_reg_3);
   assign  _net_1295 = (in_do|_reg_3);
   assign  _net_1296 = (in_do|_reg_3);
   assign  _net_1297 = (in_do|_reg_3);
   assign  _net_1298 = (in_do|_reg_3);
   assign  _net_1299 = (in_do|_reg_3);
   assign  _net_1300 = (in_do|_reg_3);
   assign  _net_1301 = (in_do|_reg_3);
   assign  _net_1302 = (in_do|_reg_3);
   assign  _net_1303 = (in_do|_reg_3);
   assign  _net_1304 = (in_do|_reg_3);
   assign  _net_1305 = (in_do|_reg_3);
   assign  _net_1306 = (in_do|_reg_3);
   assign  _net_1307 = (in_do|_reg_3);
   assign  _net_1308 = (in_do|_reg_3);
   assign  _net_1309 = (in_do|_reg_3);
   assign  _net_1310 = (in_do|_reg_3);
   assign  _net_1311 = (in_do|_reg_3);
   assign  _net_1312 = (in_do|_reg_3);
   assign  _net_1313 = (in_do|_reg_3);
   assign  _net_1314 = (in_do|_reg_3);
   assign  _net_1315 = (in_do|_reg_3);
   assign  _net_1316 = (in_do|_reg_3);
   assign  _net_1317 = (in_do|_reg_3);
   assign  _net_1318 = (in_do|_reg_3);
   assign  _net_1319 = (in_do|_reg_3);
   assign  _net_1320 = (in_do|_reg_3);
   assign  _net_1321 = (in_do|_reg_3);
   assign  _net_1322 = (in_do|_reg_3);
   assign  _net_1323 = (in_do|_reg_3);
   assign  _net_1324 = (in_do|_reg_3);
   assign  _net_1325 = (in_do|_reg_3);
   assign  _net_1326 = (in_do|_reg_3);
   assign  _net_1327 = (in_do|_reg_3);
   assign  _net_1328 = (in_do|_reg_3);
   assign  _net_1329 = (in_do|_reg_3);
   assign  _net_1330 = (in_do|_reg_3);
   assign  _net_1331 = (in_do|_reg_3);
   assign  _net_1332 = (in_do|_reg_3);
   assign  _net_1333 = (in_do|_reg_3);
   assign  _net_1334 = (in_do|_reg_3);
   assign  _net_1335 = (in_do|_reg_3);
   assign  _net_1336 = (in_do|_reg_3);
   assign  _net_1337 = (in_do|_reg_3);
   assign  _net_1338 = (in_do|_reg_3);
   assign  _net_1339 = (in_do|_reg_3);
   assign  _net_1340 = (in_do|_reg_3);
   assign  _net_1341 = (in_do|_reg_3);
   assign  _net_1342 = (in_do|_reg_3);
   assign  _net_1343 = (in_do|_reg_3);
   assign  _net_1344 = (in_do|_reg_3);
   assign  _net_1345 = (in_do|_reg_3);
   assign  _net_1346 = (in_do|_reg_3);
   assign  _net_1347 = (in_do|_reg_3);
   assign  _net_1348 = (in_do|_reg_3);
   assign  _net_1349 = (in_do|_reg_3);
   assign  _net_1350 = (in_do|_reg_3);
   assign  _net_1351 = (in_do|_reg_3);
   assign  _net_1352 = (in_do|_reg_3);
   assign  _net_1353 = (in_do|_reg_3);
   assign  _net_1354 = (in_do|_reg_3);
   assign  _net_1355 = (in_do|_reg_3);
   assign  _net_1356 = (in_do|_reg_3);
   assign  _net_1357 = (in_do|_reg_3);
   assign  _net_1358 = (in_do|_reg_3);
   assign  _net_1359 = (in_do|_reg_3);
   assign  _net_1360 = (in_do|_reg_3);
   assign  _net_1361 = (in_do|_reg_3);
   assign  _net_1362 = (in_do|_reg_3);
   assign  _net_1363 = (in_do|_reg_3);
   assign  _net_1364 = (in_do|_reg_3);
   assign  _net_1365 = (in_do|_reg_3);
   assign  _net_1366 = (in_do|_reg_3);
   assign  _net_1367 = (in_do|_reg_3);
   assign  _net_1368 = (in_do|_reg_3);
   assign  _net_1369 = (in_do|_reg_3);
   assign  _net_1370 = (in_do|_reg_3);
   assign  _net_1371 = (in_do|_reg_3);
   assign  _net_1372 = (in_do|_reg_3);
   assign  _net_1373 = (in_do|_reg_3);
   assign  _net_1374 = (in_do|_reg_3);
   assign  _net_1375 = (in_do|_reg_3);
   assign  _net_1376 = (in_do|_reg_3);
   assign  _net_1377 = (in_do|_reg_3);
   assign  _net_1378 = (in_do|_reg_3);
   assign  _net_1379 = (in_do|_reg_3);
   assign  _net_1380 = (in_do|_reg_3);
   assign  _net_1381 = (in_do|_reg_3);
   assign  _net_1382 = (in_do|_reg_3);
   assign  _net_1383 = (in_do|_reg_3);
   assign  _net_1384 = (in_do|_reg_3);
   assign  _net_1385 = (in_do|_reg_3);
   assign  _net_1386 = (in_do|_reg_3);
   assign  _net_1387 = (in_do|_reg_3);
   assign  _net_1388 = (in_do|_reg_3);
   assign  _net_1389 = (in_do|_reg_3);
   assign  _net_1390 = (in_do|_reg_3);
   assign  _net_1391 = (in_do|_reg_3);
   assign  _net_1392 = (in_do|_reg_3);
   assign  _net_1393 = (in_do|_reg_3);
   assign  _net_1394 = (in_do|_reg_3);
   assign  _net_1395 = (in_do|_reg_3);
   assign  _net_1396 = (in_do|_reg_3);
   assign  _net_1397 = (in_do|_reg_3);
   assign  _net_1398 = (in_do|_reg_3);
   assign  _net_1399 = (in_do|_reg_3);
   assign  _net_1400 = (in_do|_reg_3);
   assign  _net_1401 = (in_do|_reg_3);
   assign  _net_1402 = (in_do|_reg_3);
   assign  _net_1403 = (in_do|_reg_3);
   assign  _net_1404 = (in_do|_reg_3);
   assign  _net_1405 = (in_do|_reg_3);
   assign  _net_1406 = (in_do|_reg_3);
   assign  _net_1407 = (in_do|_reg_3);
   assign  _net_1408 = (in_do|_reg_3);
   assign  _net_1409 = (in_do|_reg_3);
   assign  _net_1410 = (in_do|_reg_3);
   assign  _net_1411 = (in_do|_reg_3);
   assign  _net_1412 = (in_do|_reg_3);
   assign  _net_1413 = (in_do|_reg_3);
   assign  _net_1414 = (in_do|_reg_3);
   assign  _net_1415 = (in_do|_reg_3);
   assign  _net_1416 = (in_do|_reg_3);
   assign  _net_1417 = (in_do|_reg_3);
   assign  _net_1418 = (in_do|_reg_3);
   assign  _net_1419 = (in_do|_reg_3);
   assign  _net_1420 = (in_do|_reg_3);
   assign  _net_1421 = (in_do|_reg_3);
   assign  _net_1422 = (in_do|_reg_3);
   assign  _net_1423 = (in_do|_reg_3);
   assign  _net_1424 = (in_do|_reg_3);
   assign  _net_1425 = (in_do|_reg_3);
   assign  _net_1426 = (in_do|_reg_3);
   assign  _net_1427 = (in_do|_reg_3);
   assign  _net_1428 = (in_do|_reg_3);
   assign  _net_1429 = (in_do|_reg_3);
   assign  _net_1430 = (in_do|_reg_3);
   assign  _net_1431 = (in_do|_reg_3);
   assign  _net_1432 = (in_do|_reg_3);
   assign  _net_1433 = (in_do|_reg_3);
   assign  _net_1434 = (in_do|_reg_3);
   assign  _net_1435 = (in_do|_reg_3);
   assign  _net_1436 = (in_do|_reg_3);
   assign  _net_1437 = (in_do|_reg_3);
   assign  _net_1438 = (in_do|_reg_3);
   assign  _net_1439 = (in_do|_reg_3);
   assign  _net_1440 = (in_do|_reg_3);
   assign  _net_1441 = (in_do|_reg_3);
   assign  _net_1442 = (in_do|_reg_3);
   assign  _net_1443 = (in_do|_reg_3);
   assign  _net_1444 = (in_do|_reg_3);
   assign  _net_1445 = (in_do|_reg_3);
   assign  _net_1446 = (in_do|_reg_3);
   assign  _net_1447 = (in_do|_reg_3);
   assign  _net_1448 = (in_do|_reg_3);
   assign  _net_1449 = (in_do|_reg_3);
   assign  _net_1450 = (in_do|_reg_3);
   assign  _net_1451 = (in_do|_reg_3);
   assign  _net_1452 = (in_do|_reg_3);
   assign  _net_1453 = (in_do|_reg_3);
   assign  _net_1454 = (in_do|_reg_3);
   assign  _net_1455 = (in_do|_reg_3);
   assign  _net_1456 = (in_do|_reg_3);
   assign  _net_1457 = (in_do|_reg_3);
   assign  _net_1458 = (in_do|_reg_3);
   assign  _net_1459 = (in_do|_reg_3);
   assign  _net_1460 = (in_do|_reg_3);
   assign  _net_1461 = (in_do|_reg_3);
   assign  _net_1462 = (in_do|_reg_3);
   assign  _net_1463 = (in_do|_reg_3);
   assign  _net_1464 = (in_do|_reg_3);
   assign  _net_1465 = (in_do|_reg_3);
   assign  _net_1466 = (in_do|_reg_3);
   assign  _net_1467 = (in_do|_reg_3);
   assign  _net_1468 = (in_do|_reg_3);
   assign  _net_1469 = (in_do|_reg_3);
   assign  _net_1470 = (in_do|_reg_3);
   assign  _net_1471 = (in_do|_reg_3);
   assign  _net_1472 = (in_do|_reg_3);
   assign  _net_1473 = (in_do|_reg_3);
   assign  _net_1474 = (in_do|_reg_3);
   assign  _net_1475 = (in_do|_reg_3);
   assign  _net_1476 = (in_do|_reg_3);
   assign  _net_1477 = (in_do|_reg_3);
   assign  _net_1478 = (in_do|_reg_3);
   assign  _net_1479 = (in_do|_reg_3);
   assign  _net_1480 = (in_do|_reg_3);
   assign  _net_1481 = (in_do|_reg_3);
   assign  _net_1482 = (in_do|_reg_3);
   assign  _net_1483 = (in_do|_reg_3);
   assign  _net_1484 = (in_do|_reg_3);
   assign  _net_1485 = (in_do|_reg_3);
   assign  _net_1486 = (in_do|_reg_3);
   assign  _net_1487 = (in_do|_reg_3);
   assign  _net_1488 = (in_do|_reg_3);
   assign  _net_1489 = (in_do|_reg_3);
   assign  _net_1490 = (in_do|_reg_3);
   assign  _net_1491 = (in_do|_reg_3);
   assign  _net_1492 = (in_do|_reg_3);
   assign  _net_1493 = (in_do|_reg_3);
   assign  _net_1494 = (in_do|_reg_3);
   assign  _net_1495 = (in_do|_reg_3);
   assign  _net_1496 = (in_do|_reg_3);
   assign  _net_1497 = (in_do|_reg_3);
   assign  _net_1498 = (in_do|_reg_3);
   assign  _net_1499 = (in_do|_reg_3);
   assign  _net_1500 = (in_do|_reg_3);
   assign  _net_1501 = (in_do|_reg_3);
   assign  _net_1502 = (in_do|_reg_3);
   assign  _net_1503 = (in_do|_reg_3);
   assign  _net_1504 = (in_do|_reg_3);
   assign  _net_1505 = (in_do|_reg_3);
   assign  _net_1506 = (in_do|_reg_3);
   assign  _net_1507 = (in_do|_reg_3);
   assign  _net_1508 = (in_do|_reg_3);
   assign  _net_1509 = (in_do|_reg_3);
   assign  _net_1510 = (in_do|_reg_3);
   assign  _net_1511 = (in_do|_reg_3);
   assign  _net_1512 = (in_do|_reg_3);
   assign  _net_1513 = (in_do|_reg_3);
   assign  _net_1514 = (in_do|_reg_3);
   assign  _net_1515 = (in_do|_reg_3);
   assign  _net_1516 = (in_do|_reg_3);
   assign  _net_1517 = (in_do|_reg_3);
   assign  _net_1518 = (in_do|_reg_3);
   assign  _net_1519 = (in_do|_reg_3);
   assign  _net_1520 = (in_do|_reg_3);
   assign  _net_1521 = (in_do|_reg_3);
   assign  _net_1522 = (in_do|_reg_3);
   assign  _net_1523 = (in_do|_reg_3);
   assign  _net_1524 = (in_do|_reg_3);
   assign  _net_1525 = (in_do|_reg_3);
   assign  _net_1526 = (in_do|_reg_3);
   assign  _net_1527 = (in_do|_reg_3);
   assign  _net_1528 = (in_do|_reg_3);
   assign  _net_1529 = (in_do|_reg_3);
   assign  _net_1530 = (in_do|_reg_3);
   assign  _net_1531 = (in_do|_reg_3);
   assign  _net_1532 = (in_do|_reg_3);
   assign  _net_1533 = (in_do|_reg_3);
   assign  _net_1534 = (in_do|_reg_3);
   assign  _net_1535 = (in_do|_reg_3);
   assign  _net_1536 = (in_do|_reg_3);
   assign  _net_1537 = (in_do|_reg_3);
   assign  _net_1538 = (in_do|_reg_3);
   assign  _net_1539 = (in_do|_reg_3);
   assign  _net_1540 = (in_do|_reg_3);
   assign  _net_1541 = (in_do|_reg_3);
   assign  _net_1542 = (in_do|_reg_3);
   assign  _net_1543 = (in_do|_reg_3);
   assign  _net_1544 = (in_do|_reg_3);
   assign  _net_1545 = (in_do|_reg_3);
   assign  _net_1546 = (in_do|_reg_3);
   assign  _net_1547 = (in_do|_reg_3);
   assign  _net_1548 = (in_do|_reg_3);
   assign  _net_1549 = (in_do|_reg_3);
   assign  _net_1550 = (in_do|_reg_3);
   assign  _net_1551 = (in_do|_reg_3);
   assign  _net_1552 = (in_do|_reg_3);
   assign  _net_1553 = (in_do|_reg_3);
   assign  _net_1554 = (in_do|_reg_3);
   assign  _net_1555 = (in_do|_reg_3);
   assign  _net_1556 = (in_do|_reg_3);
   assign  _net_1557 = (in_do|_reg_3);
   assign  _net_1558 = (in_do|_reg_3);
   assign  _net_1559 = (in_do|_reg_3);
   assign  _net_1560 = (in_do|_reg_3);
   assign  _net_1561 = (in_do|_reg_3);
   assign  _net_1562 = (in_do|_reg_3);
   assign  _net_1563 = (in_do|_reg_3);
   assign  _net_1564 = (in_do|_reg_3);
   assign  _net_1565 = (in_do|_reg_3);
   assign  _net_1566 = (in_do|_reg_3);
   assign  _net_1567 = (in_do|_reg_3);
   assign  _net_1568 = (in_do|_reg_3);
   assign  _net_1569 = (in_do|_reg_3);
   assign  _net_1570 = (in_do|_reg_3);
   assign  _net_1571 = (in_do|_reg_3);
   assign  _net_1572 = (in_do|_reg_3);
   assign  _net_1573 = (in_do|_reg_3);
   assign  _net_1574 = (in_do|_reg_3);
   assign  _net_1575 = (in_do|_reg_3);
   assign  _net_1576 = (in_do|_reg_3);
   assign  _net_1577 = (in_do|_reg_3);
   assign  _net_1578 = (in_do|_reg_3);
   assign  _net_1579 = (in_do|_reg_3);
   assign  _net_1580 = (in_do|_reg_3);
   assign  _net_1581 = (in_do|_reg_3);
   assign  _net_1582 = (in_do|_reg_3);
   assign  _net_1583 = (in_do|_reg_3);
   assign  _net_1584 = (in_do|_reg_3);
   assign  _net_1585 = (in_do|_reg_3);
   assign  _net_1586 = (in_do|_reg_3);
   assign  _net_1587 = (in_do|_reg_3);
   assign  _net_1588 = (in_do|_reg_3);
   assign  _net_1589 = (in_do|_reg_3);
   assign  _net_1590 = (in_do|_reg_3);
   assign  _net_1591 = (in_do|_reg_3);
   assign  _net_1592 = (in_do|_reg_3);
   assign  _net_1593 = (in_do|_reg_3);
   assign  _net_1594 = (in_do|_reg_3);
   assign  _net_1595 = (in_do|_reg_3);
   assign  _net_1596 = (in_do|_reg_3);
   assign  _net_1597 = (in_do|_reg_3);
   assign  _net_1598 = (in_do|_reg_3);
   assign  _net_1599 = (in_do|_reg_3);
   assign  _net_1600 = (in_do|_reg_3);
   assign  _net_1601 = (in_do|_reg_3);
   assign  _net_1602 = (in_do|_reg_3);
   assign  _net_1603 = (in_do|_reg_3);
   assign  _net_1604 = (in_do|_reg_3);
   assign  _net_1605 = (in_do|_reg_3);
   assign  _net_1606 = (in_do|_reg_3);
   assign  _net_1607 = (in_do|_reg_3);
   assign  _net_1608 = (in_do|_reg_3);
   assign  _net_1609 = (in_do|_reg_3);
   assign  _net_1610 = (in_do|_reg_3);
   assign  _net_1611 = (in_do|_reg_3);
   assign  _net_1612 = (in_do|_reg_3);
   assign  _net_1613 = (in_do|_reg_3);
   assign  _net_1614 = (in_do|_reg_3);
   assign  _net_1615 = (in_do|_reg_3);
   assign  _net_1616 = (in_do|_reg_3);
   assign  _net_1617 = (in_do|_reg_3);
   assign  _net_1618 = (in_do|_reg_3);
   assign  _net_1619 = (in_do|_reg_3);
   assign  _net_1620 = (in_do|_reg_3);
   assign  _net_1621 = (in_do|_reg_3);
   assign  _net_1622 = (in_do|_reg_3);
   assign  _net_1623 = (in_do|_reg_3);
   assign  _net_1624 = (in_do|_reg_3);
   assign  _net_1625 = (in_do|_reg_3);
   assign  _net_1626 = (in_do|_reg_3);
   assign  _net_1627 = (in_do|_reg_3);
   assign  _net_1628 = (in_do|_reg_3);
   assign  _net_1629 = (in_do|_reg_3);
   assign  _net_1630 = (in_do|_reg_3);
   assign  _net_1631 = (in_do|_reg_3);
   assign  _net_1632 = (in_do|_reg_3);
   assign  _net_1633 = (in_do|_reg_3);
   assign  _net_1634 = (in_do|_reg_3);
   assign  _net_1635 = (in_do|_reg_3);
   assign  _net_1636 = (in_do|_reg_3);
   assign  _net_1637 = (in_do|_reg_3);
   assign  _net_1638 = (in_do|_reg_3);
   assign  _net_1639 = (in_do|_reg_3);
   assign  _net_1640 = (in_do|_reg_3);
   assign  _net_1641 = (in_do|_reg_3);
   assign  _net_1642 = (in_do|_reg_3);
   assign  _net_1643 = (in_do|_reg_3);
   assign  _net_1644 = (in_do|_reg_3);
   assign  _net_1645 = (in_do|_reg_3);
   assign  _net_1646 = (in_do|_reg_3);
   assign  _net_1647 = (in_do|_reg_3);
   assign  _net_1648 = (in_do|_reg_3);
   assign  _net_1649 = (in_do|_reg_3);
   assign  _net_1650 = (in_do|_reg_3);
   assign  _net_1651 = (in_do|_reg_3);
   assign  _net_1652 = (in_do|_reg_3);
   assign  _net_1653 = (in_do|_reg_3);
   assign  _net_1654 = (in_do|_reg_3);
   assign  _net_1655 = (in_do|_reg_3);
   assign  _net_1656 = (in_do|_reg_3);
   assign  _net_1657 = (in_do|_reg_3);
   assign  _net_1658 = (in_do|_reg_3);
   assign  _net_1659 = (in_do|_reg_3);
   assign  _net_1660 = (in_do|_reg_3);
   assign  _net_1661 = (in_do|_reg_3);
   assign  _net_1662 = (in_do|_reg_3);
   assign  _net_1663 = (in_do|_reg_3);
   assign  _net_1664 = (in_do|_reg_3);
   assign  _net_1665 = (in_do|_reg_3);
   assign  _net_1666 = (in_do|_reg_3);
   assign  _net_1667 = (in_do|_reg_3);
   assign  _net_1668 = (in_do|_reg_3);
   assign  _net_1669 = (in_do|_reg_3);
   assign  _net_1670 = (in_do|_reg_3);
   assign  _net_1671 = (in_do|_reg_3);
   assign  _net_1672 = (in_do|_reg_3);
   assign  _net_1673 = (in_do|_reg_3);
   assign  _net_1674 = (in_do|_reg_3);
   assign  _net_1675 = (in_do|_reg_3);
   assign  _net_1676 = (in_do|_reg_3);
   assign  _net_1677 = (in_do|_reg_3);
   assign  _net_1678 = (in_do|_reg_3);
   assign  _net_1679 = (in_do|_reg_3);
   assign  _net_1680 = (in_do|_reg_3);
   assign  _net_1681 = (in_do|_reg_3);
   assign  _net_1682 = (in_do|_reg_3);
   assign  _net_1683 = (in_do|_reg_3);
   assign  _net_1684 = (in_do|_reg_3);
   assign  _net_1685 = (in_do|_reg_3);
   assign  _net_1686 = (in_do|_reg_3);
   assign  _net_1687 = (in_do|_reg_3);
   assign  _net_1688 = (in_do|_reg_3);
   assign  _net_1689 = (in_do|_reg_3);
   assign  _net_1690 = (in_do|_reg_3);
   assign  _net_1691 = (in_do|_reg_3);
   assign  _net_1692 = (in_do|_reg_3);
   assign  _net_1693 = (in_do|_reg_3);
   assign  _net_1694 = (in_do|_reg_3);
   assign  _net_1695 = (in_do|_reg_3);
   assign  _net_1696 = (in_do|_reg_3);
   assign  _net_1697 = (in_do|_reg_3);
   assign  _net_1698 = (in_do|_reg_3);
   assign  _net_1699 = (in_do|_reg_3);
   assign  _net_1700 = (in_do|_reg_3);
   assign  _net_1701 = (in_do|_reg_3);
   assign  _net_1702 = (in_do|_reg_3);
   assign  _net_1703 = (in_do|_reg_3);
   assign  _net_1704 = (in_do|_reg_3);
   assign  _net_1705 = (in_do|_reg_3);
   assign  _net_1706 = (in_do|_reg_3);
   assign  _net_1707 = (in_do|_reg_3);
   assign  _net_1708 = (in_do|_reg_3);
   assign  _net_1709 = (in_do|_reg_3);
   assign  _net_1710 = (in_do|_reg_3);
   assign  _net_1711 = (in_do|_reg_3);
   assign  _net_1712 = (in_do|_reg_3);
   assign  _net_1713 = (in_do|_reg_3);
   assign  _net_1714 = (in_do|_reg_3);
   assign  _net_1715 = (in_do|_reg_3);
   assign  _net_1716 = (in_do|_reg_3);
   assign  _net_1717 = (in_do|_reg_3);
   assign  _net_1718 = (in_do|_reg_3);
   assign  _net_1719 = (in_do|_reg_3);
   assign  _net_1720 = (in_do|_reg_3);
   assign  _net_1721 = (in_do|_reg_3);
   assign  _net_1722 = (in_do|_reg_3);
   assign  _net_1723 = (in_do|_reg_3);
   assign  _net_1724 = (in_do|_reg_3);
   assign  _net_1725 = (in_do|_reg_3);
   assign  _net_1726 = (in_do|_reg_3);
   assign  _net_1727 = (in_do|_reg_3);
   assign  _net_1728 = (in_do|_reg_3);
   assign  _net_1729 = (in_do|_reg_3);
   assign  _net_1730 = (in_do|_reg_3);
   assign  _net_1731 = (in_do|_reg_3);
   assign  _net_1732 = (in_do|_reg_3);
   assign  _net_1733 = (in_do|_reg_3);
   assign  _net_1734 = (in_do|_reg_3);
   assign  _net_1735 = (in_do|_reg_3);
   assign  _net_1736 = (in_do|_reg_3);
   assign  _net_1737 = (in_do|_reg_3);
   assign  _net_1738 = (in_do|_reg_3);
   assign  _net_1739 = (in_do|_reg_3);
   assign  _net_1740 = (in_do|_reg_3);
   assign  _net_1741 = (in_do|_reg_3);
   assign  _net_1742 = (in_do|_reg_3);
   assign  _net_1743 = (in_do|_reg_3);
   assign  _net_1744 = (in_do|_reg_3);
   assign  _net_1745 = (in_do|_reg_3);
   assign  _net_1746 = (in_do|_reg_3);
   assign  _net_1747 = (in_do|_reg_3);
   assign  _net_1748 = (in_do|_reg_3);
   assign  _net_1749 = (in_do|_reg_3);
   assign  _net_1750 = (in_do|_reg_3);
   assign  _net_1751 = (in_do|_reg_3);
   assign  _net_1752 = (in_do|_reg_3);
   assign  _net_1753 = (in_do|_reg_3);
   assign  _net_1754 = (in_do|_reg_3);
   assign  _net_1755 = (in_do|_reg_3);
   assign  _net_1756 = (in_do|_reg_3);
   assign  _net_1757 = (in_do|_reg_3);
   assign  _net_1758 = (in_do|_reg_3);
   assign  _net_1759 = (in_do|_reg_3);
   assign  _net_1760 = (in_do|_reg_3);
   assign  _net_1761 = (in_do|_reg_3);
   assign  _net_1762 = (in_do|_reg_3);
   assign  _net_1763 = (in_do|_reg_3);
   assign  _net_1764 = (in_do|_reg_3);
   assign  _net_1765 = (in_do|_reg_3);
   assign  _net_1766 = (in_do|_reg_3);
   assign  _net_1767 = (in_do|_reg_3);
   assign  _net_1768 = (in_do|_reg_3);
   assign  _net_1769 = (in_do|_reg_3);
   assign  _net_1770 = (in_do|_reg_3);
   assign  _net_1771 = (in_do|_reg_3);
   assign  _net_1772 = (in_do|_reg_3);
   assign  _net_1773 = (in_do|_reg_3);
   assign  _net_1774 = (in_do|_reg_3);
   assign  _net_1775 = (in_do|_reg_3);
   assign  _net_1776 = (in_do|_reg_3);
   assign  _net_1777 = (in_do|_reg_3);
   assign  _net_1778 = (in_do|_reg_3);
   assign  _net_1779 = (in_do|_reg_3);
   assign  _net_1780 = (in_do|_reg_3);
   assign  _net_1781 = (in_do|_reg_3);
   assign  _net_1782 = (in_do|_reg_3);
   assign  _net_1783 = (in_do|_reg_3);
   assign  _net_1784 = (in_do|_reg_3);
   assign  _net_1785 = (in_do|_reg_3);
   assign  _net_1786 = (in_do|_reg_3);
   assign  _net_1787 = (in_do|_reg_3);
   assign  _net_1788 = (in_do|_reg_3);
   assign  _net_1789 = (in_do|_reg_3);
   assign  _net_1790 = (in_do|_reg_3);
   assign  _net_1791 = (in_do|_reg_3);
   assign  _net_1792 = (in_do|_reg_3);
   assign  _net_1793 = (in_do|_reg_3);
   assign  _net_1794 = (in_do|_reg_3);
   assign  _net_1795 = (in_do|_reg_3);
   assign  _net_1796 = (in_do|_reg_3);
   assign  _net_1797 = (in_do|_reg_3);
   assign  _net_1798 = (in_do|_reg_3);
   assign  _net_1799 = (in_do|_reg_3);
   assign  _net_1800 = (in_do|_reg_3);
   assign  _net_1801 = (in_do|_reg_3);
   assign  _net_1802 = (in_do|_reg_3);
   assign  _net_1803 = (in_do|_reg_3);
   assign  _net_1804 = (in_do|_reg_3);
   assign  _net_1805 = (in_do|_reg_3);
   assign  _net_1806 = (in_do|_reg_3);
   assign  _net_1807 = (in_do|_reg_3);
   assign  _net_1808 = (in_do|_reg_3);
   assign  _net_1809 = (in_do|_reg_3);
   assign  _net_1810 = (in_do|_reg_3);
   assign  _net_1811 = (in_do|_reg_3);
   assign  _net_1812 = (in_do|_reg_3);
   assign  _net_1813 = (in_do|_reg_3);
   assign  _net_1814 = (in_do|_reg_3);
   assign  _net_1815 = (in_do|_reg_3);
   assign  _net_1816 = (in_do|_reg_3);
   assign  _net_1817 = (in_do|_reg_3);
   assign  _net_1818 = (in_do|_reg_3);
   assign  _net_1819 = (in_do|_reg_3);
   assign  _net_1820 = (in_do|_reg_3);
   assign  _net_1821 = (in_do|_reg_3);
   assign  _net_1822 = (in_do|_reg_3);
   assign  _net_1823 = (in_do|_reg_3);
   assign  _net_1824 = (in_do|_reg_3);
   assign  _net_1825 = (in_do|_reg_3);
   assign  _net_1826 = (in_do|_reg_3);
   assign  _net_1827 = (in_do|_reg_3);
   assign  _net_1828 = (in_do|_reg_3);
   assign  _net_1829 = (in_do|_reg_3);
   assign  _net_1830 = (in_do|_reg_3);
   assign  _net_1831 = (in_do|_reg_3);
   assign  _net_1832 = (in_do|_reg_3);
   assign  _net_1833 = (in_do|_reg_3);
   assign  _net_1834 = (in_do|_reg_3);
   assign  _net_1835 = (in_do|_reg_3);
   assign  _net_1836 = (in_do|_reg_3);
   assign  _net_1837 = (in_do|_reg_3);
   assign  _net_1838 = (in_do|_reg_3);
   assign  _net_1839 = (in_do|_reg_3);
   assign  _net_1840 = (in_do|_reg_3);
   assign  _net_1841 = (in_do|_reg_3);
   assign  _net_1842 = (in_do|_reg_3);
   assign  _net_1843 = (in_do|_reg_3);
   assign  _net_1844 = (in_do|_reg_3);
   assign  _net_1845 = (in_do|_reg_3);
   assign  _net_1846 = (in_do|_reg_3);
   assign  _net_1847 = (in_do|_reg_3);
   assign  _net_1848 = (in_do|_reg_3);
   assign  _net_1849 = (in_do|_reg_3);
   assign  _net_1850 = (in_do|_reg_3);
   assign  _net_1851 = (in_do|_reg_3);
   assign  _net_1852 = (in_do|_reg_3);
   assign  _net_1853 = (in_do|_reg_3);
   assign  _net_1854 = (in_do|_reg_3);
   assign  _net_1855 = (in_do|_reg_3);
   assign  _net_1856 = (in_do|_reg_3);
   assign  _net_1857 = (in_do|_reg_3);
   assign  _net_1858 = (in_do|_reg_3);
   assign  _net_1859 = (in_do|_reg_3);
   assign  _net_1860 = (in_do|_reg_3);
   assign  _net_1861 = (in_do|_reg_3);
   assign  _net_1862 = (in_do|_reg_3);
   assign  _net_1863 = (in_do|_reg_3);
   assign  _net_1864 = (in_do|_reg_3);
   assign  _net_1865 = (in_do|_reg_3);
   assign  _net_1866 = (in_do|_reg_3);
   assign  _net_1867 = (in_do|_reg_3);
   assign  _net_1868 = (in_do|_reg_3);
   assign  _net_1869 = (in_do|_reg_3);
   assign  _net_1870 = (in_do|_reg_3);
   assign  _net_1871 = (in_do|_reg_3);
   assign  _net_1872 = (in_do|_reg_3);
   assign  _net_1873 = (in_do|_reg_3);
   assign  _net_1874 = (in_do|_reg_3);
   assign  _net_1875 = (in_do|_reg_3);
   assign  _net_1876 = (in_do|_reg_3);
   assign  _net_1877 = (in_do|_reg_3);
   assign  _net_1878 = (in_do|_reg_3);
   assign  _net_1879 = (in_do|_reg_3);
   assign  _net_1880 = (in_do|_reg_3);
   assign  _net_1881 = (in_do|_reg_3);
   assign  _net_1882 = (in_do|_reg_3);
   assign  _net_1883 = (in_do|_reg_3);
   assign  _net_1884 = (in_do|_reg_3);
   assign  _net_1885 = (in_do|_reg_3);
   assign  _net_1886 = (in_do|_reg_3);
   assign  _net_1887 = (in_do|_reg_3);
   assign  _net_1888 = (in_do|_reg_3);
   assign  _net_1889 = (in_do|_reg_3);
   assign  _net_1890 = (in_do|_reg_3);
   assign  _net_1891 = (in_do|_reg_3);
   assign  _net_1892 = (in_do|_reg_3);
   assign  _net_1893 = (in_do|_reg_3);
   assign  _net_1894 = (in_do|_reg_3);
   assign  _net_1895 = (in_do|_reg_3);
   assign  _net_1896 = (in_do|_reg_3);
   assign  _net_1897 = (in_do|_reg_3);
   assign  _net_1898 = (in_do|_reg_3);
   assign  _net_1899 = (in_do|_reg_3);
   assign  _net_1900 = (in_do|_reg_3);
   assign  _net_1901 = (in_do|_reg_3);
   assign  _net_1902 = (in_do|_reg_3);
   assign  _net_1903 = (in_do|_reg_3);
   assign  _net_1904 = (in_do|_reg_3);
   assign  _net_1905 = (in_do|_reg_3);
   assign  _net_1906 = (in_do|_reg_3);
   assign  _net_1907 = (in_do|_reg_3);
   assign  _net_1908 = (in_do|_reg_3);
   assign  _net_1909 = (in_do|_reg_3);
   assign  _net_1910 = (in_do|_reg_3);
   assign  _net_1911 = (in_do|_reg_3);
   assign  _net_1912 = (in_do|_reg_3);
   assign  _net_1913 = (in_do|_reg_3);
   assign  _net_1914 = (in_do|_reg_3);
   assign  _net_1915 = (in_do|_reg_3);
   assign  _net_1916 = (in_do|_reg_3);
   assign  _net_1917 = (in_do|_reg_3);
   assign  _net_1918 = (in_do|_reg_3);
   assign  _net_1919 = (in_do|_reg_3);
   assign  _net_1920 = (in_do|_reg_3);
   assign  _net_1921 = (in_do|_reg_3);
   assign  _net_1922 = (in_do|_reg_3);
   assign  _net_1923 = (in_do|_reg_3);
   assign  _net_1924 = (in_do|_reg_3);
   assign  _net_1925 = (in_do|_reg_3);
   assign  _net_1926 = (in_do|_reg_3);
   assign  _net_1927 = (in_do|_reg_3);
   assign  _net_1928 = (in_do|_reg_3);
   assign  _net_1929 = (in_do|_reg_3);
   assign  _net_1930 = (in_do|_reg_3);
   assign  _net_1931 = (in_do|_reg_3);
   assign  _net_1932 = (in_do|_reg_3);
   assign  _net_1933 = (in_do|_reg_3);
   assign  _net_1934 = (in_do|_reg_3);
   assign  _net_1935 = (in_do|_reg_3);
   assign  _net_1936 = (in_do|_reg_3);
   assign  _net_1937 = (in_do|_reg_3);
   assign  _net_1938 = (in_do|_reg_3);
   assign  _net_1939 = (in_do|_reg_3);
   assign  _net_1940 = (in_do|_reg_3);
   assign  _net_1941 = (in_do|_reg_3);
   assign  _net_1942 = (in_do|_reg_3);
   assign  _net_1943 = (in_do|_reg_3);
   assign  _net_1944 = (in_do|_reg_3);
   assign  _net_1945 = (in_do|_reg_3);
   assign  _net_1946 = (in_do|_reg_3);
   assign  _net_1947 = (in_do|_reg_3);
   assign  _net_1948 = (in_do|_reg_3);
   assign  _net_1949 = (in_do|_reg_3);
   assign  _net_1950 = (in_do|_reg_3);
   assign  _net_1951 = (in_do|_reg_3);
   assign  _net_1952 = (in_do|_reg_3);
   assign  _net_1953 = (in_do|_reg_3);
   assign  _net_1954 = (in_do|_reg_3);
   assign  _net_1955 = (in_do|_reg_3);
   assign  _net_1956 = (in_do|_reg_3);
   assign  _net_1957 = (in_do|_reg_3);
   assign  _net_1958 = (in_do|_reg_3);
   assign  _net_1959 = (in_do|_reg_3);
   assign  _net_1960 = (in_do|_reg_3);
   assign  _net_1961 = (in_do|_reg_3);
   assign  _net_1962 = (in_do|_reg_3);
   assign  _net_1963 = (in_do|_reg_3);
   assign  _net_1964 = (in_do|_reg_3);
   assign  _net_1965 = (in_do|_reg_3);
   assign  _net_1966 = (in_do|_reg_3);
   assign  _net_1967 = (in_do|_reg_3);
   assign  _net_1968 = (in_do|_reg_3);
   assign  _net_1969 = (in_do|_reg_3);
   assign  _net_1970 = (in_do|_reg_3);
   assign  _net_1971 = (in_do|_reg_3);
   assign  _net_1972 = (in_do|_reg_3);
   assign  _net_1973 = (in_do|_reg_3);
   assign  _net_1974 = (in_do|_reg_3);
   assign  _net_1975 = (in_do|_reg_3);
   assign  _net_1976 = (in_do|_reg_3);
   assign  _net_1977 = (in_do|_reg_3);
   assign  _net_1978 = (in_do|_reg_3);
   assign  _net_1979 = (in_do|_reg_3);
   assign  _net_1980 = (in_do|_reg_3);
   assign  _net_1981 = (in_do|_reg_3);
   assign  _net_1982 = (in_do|_reg_3);
   assign  _net_1983 = (in_do|_reg_3);
   assign  _net_1984 = (in_do|_reg_3);
   assign  _net_1985 = (in_do|_reg_3);
   assign  _net_1986 = (in_do|_reg_3);
   assign  _net_1987 = (in_do|_reg_3);
   assign  _net_1988 = (in_do|_reg_3);
   assign  _net_1989 = (in_do|_reg_3);
   assign  _net_1990 = (in_do|_reg_3);
   assign  _net_1991 = (in_do|_reg_3);
   assign  _net_1992 = (in_do|_reg_3);
   assign  _net_1993 = (in_do|_reg_3);
   assign  _net_1994 = (in_do|_reg_3);
   assign  _net_1995 = (in_do|_reg_3);
   assign  _net_1996 = (in_do|_reg_3);
   assign  _net_1997 = (in_do|_reg_3);
   assign  _net_1998 = (in_do|_reg_3);
   assign  _net_1999 = (in_do|_reg_3);
   assign  _net_2000 = (in_do|_reg_3);
   assign  _net_2001 = (in_do|_reg_3);
   assign  _net_2002 = (in_do|_reg_3);
   assign  _net_2003 = (in_do|_reg_3);
   assign  _net_2004 = (in_do|_reg_3);
   assign  _net_2005 = (in_do|_reg_3);
   assign  _net_2006 = (in_do|_reg_3);
   assign  _net_2007 = (in_do|_reg_3);
   assign  _net_2008 = (in_do|_reg_3);
   assign  _net_2009 = (in_do|_reg_3);
   assign  _net_2010 = (in_do|_reg_3);
   assign  _net_2011 = (in_do|_reg_3);
   assign  _net_2012 = (in_do|_reg_3);
   assign  _net_2013 = (in_do|_reg_3);
   assign  _net_2014 = (in_do|_reg_3);
   assign  _net_2015 = (in_do|_reg_3);
   assign  _net_2016 = (in_do|_reg_3);
   assign  _net_2017 = (in_do|_reg_3);
   assign  _net_2018 = (in_do|_reg_3);
   assign  _net_2019 = (in_do|_reg_3);
   assign  _net_2020 = (in_do|_reg_3);
   assign  _net_2021 = (in_do|_reg_3);
   assign  _net_2022 = (in_do|_reg_3);
   assign  _net_2023 = (in_do|_reg_3);
   assign  _net_2024 = (in_do|_reg_3);
   assign  _net_2025 = (in_do|_reg_3);
   assign  _net_2026 = (in_do|_reg_3);
   assign  _net_2027 = (in_do|_reg_3);
   assign  _net_2028 = (in_do|_reg_3);
   assign  _net_2029 = (in_do|_reg_3);
   assign  _net_2030 = (in_do|_reg_3);
   assign  _net_2031 = (in_do|_reg_3);
   assign  _net_2032 = (in_do|_reg_3);
   assign  _net_2033 = (in_do|_reg_3);
   assign  _net_2034 = (in_do|_reg_3);
   assign  _net_2035 = (in_do|_reg_3);
   assign  _net_2036 = (in_do|_reg_3);
   assign  _net_2037 = (in_do|_reg_3);
   assign  _net_2038 = (in_do|_reg_3);
   assign  _net_2039 = (in_do|_reg_3);
   assign  _net_2040 = (in_do|_reg_3);
   assign  _net_2041 = (in_do|_reg_3);
   assign  _net_2042 = (in_do|_reg_3);
   assign  _net_2043 = (in_do|_reg_3);
   assign  _net_2044 = (in_do|_reg_3);
   assign  _net_2045 = (in_do|_reg_3);
   assign  _net_2046 = (in_do|_reg_3);
   assign  _net_2047 = (in_do|_reg_3);
   assign  _net_2048 = (in_do|_reg_3);
   assign  _net_2049 = (in_do|_reg_3);
   assign  _net_2050 = (in_do|_reg_3);
   assign  _net_2051 = (in_do|_reg_3);
   assign  _net_2052 = (in_do|_reg_3);
   assign  _net_2053 = (in_do|_reg_3);
   assign  _net_2054 = (in_do|_reg_3);
   assign  _net_2055 = (in_do|_reg_3);
   assign  _net_2056 = (in_do|_reg_3);
   assign  _net_2057 = (in_do|_reg_3);
   assign  _net_2058 = (in_do|_reg_3);
   assign  _net_2059 = (in_do|_reg_3);
   assign  _net_2060 = (in_do|_reg_3);
   assign  _net_2061 = (in_do|_reg_3);
   assign  _net_2062 = (in_do|_reg_3);
   assign  _net_2063 = (in_do|_reg_3);
   assign  _net_2064 = (in_do|_reg_3);
   assign  _net_2065 = (in_do|_reg_3);
   assign  _net_2066 = (in_do|_reg_3);
   assign  _net_2067 = (in_do|_reg_3);
   assign  _net_2068 = (in_do|_reg_3);
   assign  _net_2069 = (in_do|_reg_3);
   assign  _net_2070 = (in_do|_reg_3);
   assign  _net_2071 = (in_do|_reg_3);
   assign  _net_2072 = (in_do|_reg_3);
   assign  _net_2073 = (in_do|_reg_3);
   assign  _net_2074 = (in_do|_reg_3);
   assign  _net_2075 = (in_do|_reg_3);
   assign  _net_2076 = (in_do|_reg_3);
   assign  _net_2077 = (in_do|_reg_3);
   assign  _net_2078 = (in_do|_reg_3);
   assign  _net_2079 = (in_do|_reg_3);
   assign  _net_2080 = (in_do|_reg_3);
   assign  _net_2081 = (in_do|_reg_3);
   assign  _net_2082 = (in_do|_reg_3);
   assign  _net_2083 = (in_do|_reg_3);
   assign  _net_2084 = (in_do|_reg_3);
   assign  _net_2085 = (in_do|_reg_3);
   assign  _net_2086 = (in_do|_reg_3);
   assign  _net_2087 = (in_do|_reg_3);
   assign  _net_2088 = (in_do|_reg_3);
   assign  _net_2089 = (in_do|_reg_3);
   assign  _net_2090 = (in_do|_reg_3);
   assign  _net_2091 = (in_do|_reg_3);
   assign  _net_2092 = (in_do|_reg_3);
   assign  _net_2093 = (in_do|_reg_3);
   assign  _net_2094 = (in_do|_reg_3);
   assign  _net_2095 = (in_do|_reg_3);
   assign  _net_2096 = (in_do|_reg_3);
   assign  _net_2097 = (in_do|_reg_3);
   assign  _net_2098 = (in_do|_reg_3);
   assign  _net_2099 = (in_do|_reg_3);
   assign  _net_2100 = (in_do|_reg_3);
   assign  _net_2101 = (in_do|_reg_3);
   assign  _net_2102 = (in_do|_reg_3);
   assign  _net_2103 = (in_do|_reg_3);
   assign  _net_2104 = (in_do|_reg_3);
   assign  _net_2105 = (in_do|_reg_3);
   assign  _net_2106 = (in_do|_reg_3);
   assign  _net_2107 = (in_do|_reg_3);
   assign  _net_2108 = (in_do|_reg_3);
   assign  _net_2109 = (in_do|_reg_3);
   assign  _net_2110 = (in_do|_reg_3);
   assign  _net_2111 = (in_do|_reg_3);
   assign  _net_2112 = (in_do|_reg_3);
   assign  _net_2113 = (in_do|_reg_3);
   assign  _net_2114 = (in_do|_reg_3);
   assign  _net_2115 = (in_do|_reg_3);
   assign  _net_2116 = (in_do|_reg_3);
   assign  _net_2117 = (in_do|_reg_3);
   assign  _net_2118 = (in_do|_reg_3);
   assign  _net_2119 = (in_do|_reg_3);
   assign  _net_2120 = (in_do|_reg_3);
   assign  _net_2121 = (in_do|_reg_3);
   assign  _net_2122 = (in_do|_reg_3);
   assign  _net_2123 = (in_do|_reg_3);
   assign  _net_2124 = (in_do|_reg_3);
   assign  _net_2125 = (in_do|_reg_3);
   assign  _net_2126 = (in_do|_reg_3);
   assign  _net_2127 = (in_do|_reg_3);
   assign  _net_2128 = (in_do|_reg_3);
   assign  _net_2129 = (in_do|_reg_3);
   assign  _net_2130 = (in_do|_reg_3);
   assign  _net_2131 = (in_do|_reg_3);
   assign  _net_2132 = (in_do|_reg_3);
   assign  _net_2133 = (in_do|_reg_3);
   assign  _net_2134 = (in_do|_reg_3);
   assign  _net_2135 = (in_do|_reg_3);
   assign  _net_2136 = (in_do|_reg_3);
   assign  _net_2137 = (in_do|_reg_3);
   assign  _net_2138 = (in_do|_reg_3);
   assign  _net_2139 = (in_do|_reg_3);
   assign  _net_2140 = (in_do|_reg_3);
   assign  _net_2141 = (in_do|_reg_3);
   assign  _net_2142 = (in_do|_reg_3);
   assign  _net_2143 = (in_do|_reg_3);
   assign  _net_2144 = (in_do|_reg_3);
   assign  _net_2145 = (in_do|_reg_3);
   assign  _net_2146 = (in_do|_reg_3);
   assign  _net_2147 = (in_do|_reg_3);
   assign  _net_2148 = (in_do|_reg_3);
   assign  _net_2149 = (in_do|_reg_3);
   assign  _net_2150 = (in_do|_reg_3);
   assign  _net_2151 = (in_do|_reg_3);
   assign  _net_2152 = (in_do|_reg_3);
   assign  _net_2153 = (in_do|_reg_3);
   assign  _net_2154 = (in_do|_reg_3);
   assign  _net_2155 = (in_do|_reg_3);
   assign  _net_2156 = (in_do|_reg_3);
   assign  _net_2157 = (in_do|_reg_3);
   assign  _net_2158 = (in_do|_reg_3);
   assign  _net_2159 = (in_do|_reg_3);
   assign  _net_2160 = (in_do|_reg_3);
   assign  _net_2161 = (in_do|_reg_3);
   assign  _net_2162 = (in_do|_reg_3);
   assign  _net_2163 = (in_do|_reg_3);
   assign  _net_2164 = (in_do|_reg_3);
   assign  _net_2165 = (in_do|_reg_3);
   assign  _net_2166 = (in_do|_reg_3);
   assign  _net_2167 = (in_do|_reg_3);
   assign  _net_2168 = (in_do|_reg_3);
   assign  _net_2169 = (in_do|_reg_3);
   assign  _net_2170 = (in_do|_reg_3);
   assign  _net_2171 = (in_do|_reg_3);
   assign  _net_2172 = (in_do|_reg_3);
   assign  _net_2173 = (in_do|_reg_3);
   assign  _net_2174 = (in_do|_reg_3);
   assign  _net_2175 = (in_do|_reg_3);
   assign  _net_2176 = (in_do|_reg_3);
   assign  _net_2177 = (in_do|_reg_3);
   assign  _net_2178 = (in_do|_reg_3);
   assign  _net_2179 = (in_do|_reg_3);
   assign  _net_2180 = (in_do|_reg_3);
   assign  _net_2181 = (in_do|_reg_3);
   assign  _net_2182 = (in_do|_reg_3);
   assign  _net_2183 = (in_do|_reg_3);
   assign  _net_2184 = (in_do|_reg_3);
   assign  _net_2185 = (in_do|_reg_3);
   assign  _net_2186 = (in_do|_reg_3);
   assign  _net_2187 = (in_do|_reg_3);
   assign  _net_2188 = (in_do|_reg_3);
   assign  _net_2189 = (in_do|_reg_3);
   assign  _net_2190 = (in_do|_reg_3);
   assign  _net_2191 = (in_do|_reg_3);
   assign  _net_2192 = (in_do|_reg_3);
   assign  _net_2193 = (in_do|_reg_3);
   assign  _net_2194 = (in_do|_reg_3);
   assign  _net_2195 = (in_do|_reg_3);
   assign  _net_2196 = (in_do|_reg_3);
   assign  _net_2197 = (in_do|_reg_3);
   assign  _net_2198 = (in_do|_reg_3);
   assign  _net_2199 = (in_do|_reg_3);
   assign  _net_2200 = (in_do|_reg_3);
   assign  _net_2201 = (in_do|_reg_3);
   assign  _net_2202 = (in_do|_reg_3);
   assign  _net_2203 = (in_do|_reg_3);
   assign  _net_2204 = (in_do|_reg_3);
   assign  _net_2205 = (in_do|_reg_3);
   assign  _net_2206 = (in_do|_reg_3);
   assign  _net_2207 = (in_do|_reg_3);
   assign  _net_2208 = (in_do|_reg_3);
   assign  _net_2209 = (in_do|_reg_3);
   assign  _net_2210 = (in_do|_reg_3);
   assign  _net_2211 = (in_do|_reg_3);
   assign  _net_2212 = (in_do|_reg_3);
   assign  _net_2213 = (in_do|_reg_3);
   assign  _net_2214 = (in_do|_reg_3);
   assign  _net_2215 = (in_do|_reg_3);
   assign  _net_2216 = (in_do|_reg_3);
   assign  _net_2217 = (in_do|_reg_3);
   assign  _net_2218 = (in_do|_reg_3);
   assign  _net_2219 = (in_do|_reg_3);
   assign  _net_2220 = (in_do|_reg_3);
   assign  _net_2221 = (in_do|_reg_3);
   assign  _net_2222 = (in_do|_reg_3);
   assign  _net_2223 = (in_do|_reg_3);
   assign  _net_2224 = (in_do|_reg_3);
   assign  _net_2225 = (in_do|_reg_3);
   assign  _net_2226 = (in_do|_reg_3);
   assign  _net_2227 = (in_do|_reg_3);
   assign  _net_2228 = (in_do|_reg_3);
   assign  _net_2229 = (in_do|_reg_3);
   assign  _net_2230 = (in_do|_reg_3);
   assign  _net_2231 = (in_do|_reg_3);
   assign  _net_2232 = (in_do|_reg_3);
   assign  _net_2233 = (in_do|_reg_3);
   assign  _net_2234 = (in_do|_reg_3);
   assign  _net_2235 = (in_do|_reg_3);
   assign  _net_2236 = (in_do|_reg_3);
   assign  _net_2237 = (in_do|_reg_3);
   assign  _net_2238 = (in_do|_reg_3);
   assign  _net_2239 = (in_do|_reg_3);
   assign  _net_2240 = (in_do|_reg_3);
   assign  _net_2241 = (in_do|_reg_3);
   assign  _net_2242 = (in_do|_reg_3);
   assign  _net_2243 = (in_do|_reg_3);
   assign  _net_2244 = (in_do|_reg_3);
   assign  _net_2245 = (in_do|_reg_3);
   assign  _net_2246 = (in_do|_reg_3);
   assign  _net_2247 = (in_do|_reg_3);
   assign  _net_2248 = (in_do|_reg_3);
   assign  _net_2249 = (in_do|_reg_3);
   assign  _net_2250 = (in_do|_reg_3);
   assign  _net_2251 = (in_do|_reg_3);
   assign  _net_2252 = (in_do|_reg_3);
   assign  _net_2253 = (in_do|_reg_3);
   assign  _net_2254 = (in_do|_reg_3);
   assign  _net_2255 = (in_do|_reg_3);
   assign  _net_2256 = (in_do|_reg_3);
   assign  _net_2257 = (in_do|_reg_3);
   assign  _net_2258 = (in_do|_reg_3);
   assign  _net_2259 = (in_do|_reg_3);
   assign  _net_2260 = (in_do|_reg_3);
   assign  _net_2261 = (in_do|_reg_3);
   assign  _net_2262 = (in_do|_reg_3);
   assign  _net_2263 = (in_do|_reg_3);
   assign  _net_2264 = (in_do|_reg_3);
   assign  _net_2265 = (in_do|_reg_3);
   assign  _net_2266 = (in_do|_reg_3);
   assign  _net_2267 = (in_do|_reg_3);
   assign  _net_2268 = (in_do|_reg_3);
   assign  _net_2269 = (in_do|_reg_3);
   assign  _net_2270 = (in_do|_reg_3);
   assign  _net_2271 = (in_do|_reg_3);
   assign  _net_2272 = (in_do|_reg_3);
   assign  _net_2273 = (in_do|_reg_3);
   assign  _net_2274 = (in_do|_reg_3);
   assign  _net_2275 = (in_do|_reg_3);
   assign  _net_2276 = (in_do|_reg_3);
   assign  _net_2277 = (in_do|_reg_3);
   assign  _net_2278 = (in_do|_reg_3);
   assign  _net_2279 = (in_do|_reg_3);
   assign  _net_2280 = (in_do|_reg_3);
   assign  _net_2281 = (in_do|_reg_3);
   assign  _net_2282 = (in_do|_reg_3);
   assign  _net_2283 = (in_do|_reg_3);
   assign  _net_2284 = (in_do|_reg_3);
   assign  _net_2285 = (in_do|_reg_3);
   assign  _net_2286 = (in_do|_reg_3);
   assign  _net_2287 = (in_do|_reg_3);
   assign  _net_2288 = (in_do|_reg_3);
   assign  _net_2289 = (in_do|_reg_3);
   assign  _net_2290 = (in_do|_reg_3);
   assign  _net_2291 = (in_do|_reg_3);
   assign  _net_2292 = (in_do|_reg_3);
   assign  _net_2293 = (in_do|_reg_3);
   assign  _net_2294 = (in_do|_reg_3);
   assign  _net_2295 = (in_do|_reg_3);
   assign  _net_2296 = (in_do|_reg_3);
   assign  _net_2297 = (in_do|_reg_3);
   assign  _net_2298 = (in_do|_reg_3);
   assign  _net_2299 = (in_do|_reg_3);
   assign  _net_2300 = (in_do|_reg_3);
   assign  _net_2301 = (in_do|_reg_3);
   assign  _net_2302 = (in_do|_reg_3);
   assign  _net_2303 = (in_do|_reg_3);
   assign  _net_2304 = (in_do|_reg_3);
   assign  _net_2305 = (in_do|_reg_3);
   assign  _net_2306 = (in_do|_reg_3);
   assign  _net_2307 = (in_do|_reg_3);
   assign  _net_2308 = (in_do|_reg_3);
   assign  _net_2309 = (in_do|_reg_3);
   assign  _net_2310 = (in_do|_reg_3);
   assign  _net_2311 = (in_do|_reg_3);
   assign  _net_2312 = (in_do|_reg_3);
   assign  _net_2313 = (in_do|_reg_3);
   assign  _net_2314 = (in_do|_reg_3);
   assign  _net_2315 = (in_do|_reg_3);
   assign  _net_2316 = (in_do|_reg_3);
   assign  _net_2317 = (in_do|_reg_3);
   assign  _net_2318 = (in_do|_reg_3);
   assign  _net_2319 = (in_do|_reg_3);
   assign  _net_2320 = (in_do|_reg_3);
   assign  _net_2321 = (in_do|_reg_3);
   assign  _net_2322 = (in_do|_reg_3);
   assign  _net_2323 = (in_do|_reg_3);
   assign  _net_2324 = (in_do|_reg_3);
   assign  _net_2325 = (in_do|_reg_3);
   assign  _net_2326 = (in_do|_reg_3);
   assign  _net_2327 = (in_do|_reg_3);
   assign  _net_2328 = (in_do|_reg_3);
   assign  _net_2329 = (in_do|_reg_3);
   assign  _net_2330 = (in_do|_reg_3);
   assign  _net_2331 = (in_do|_reg_3);
   assign  _net_2332 = (in_do|_reg_3);
   assign  _net_2333 = (in_do|_reg_3);
   assign  _net_2334 = (in_do|_reg_3);
   assign  _net_2335 = (in_do|_reg_3);
   assign  _net_2336 = (in_do|_reg_3);
   assign  _net_2337 = (in_do|_reg_3);
   assign  _net_2338 = (in_do|_reg_3);
   assign  _net_2339 = (in_do|_reg_3);
   assign  _net_2340 = (in_do|_reg_3);
   assign  _net_2341 = (in_do|_reg_3);
   assign  _net_2342 = (in_do|_reg_3);
   assign  _net_2343 = (in_do|_reg_3);
   assign  _net_2344 = (in_do|_reg_3);
   assign  _net_2345 = (in_do|_reg_3);
   assign  _net_2346 = (in_do|_reg_3);
   assign  _net_2347 = (in_do|_reg_3);
   assign  _net_2348 = (in_do|_reg_3);
   assign  _net_2349 = (in_do|_reg_3);
   assign  _net_2350 = (in_do|_reg_3);
   assign  _net_2351 = (in_do|_reg_3);
   assign  _net_2352 = (in_do|_reg_3);
   assign  _net_2353 = (in_do|_reg_3);
   assign  _net_2354 = (in_do|_reg_3);
   assign  _net_2355 = (in_do|_reg_3);
   assign  _net_2356 = (in_do|_reg_3);
   assign  _net_2357 = (in_do|_reg_3);
   assign  _net_2358 = (in_do|_reg_3);
   assign  _net_2359 = (in_do|_reg_3);
   assign  _net_2360 = (in_do|_reg_3);
   assign  _net_2361 = (in_do|_reg_3);
   assign  _net_2362 = (in_do|_reg_3);
   assign  _net_2363 = (in_do|_reg_3);
   assign  _net_2364 = (in_do|_reg_3);
   assign  _net_2365 = (in_do|_reg_3);
   assign  _net_2366 = (in_do|_reg_3);
   assign  _net_2367 = (in_do|_reg_3);
   assign  _net_2368 = (in_do|_reg_3);
   assign  _net_2369 = (in_do|_reg_3);
   assign  _net_2370 = (in_do|_reg_3);
   assign  _net_2371 = (in_do|_reg_3);
   assign  _net_2372 = (in_do|_reg_3);
   assign  _net_2373 = (in_do|_reg_3);
   assign  _net_2374 = (in_do|_reg_3);
   assign  _net_2375 = (in_do|_reg_3);
   assign  _net_2376 = (in_do|_reg_3);
   assign  _net_2377 = (in_do|_reg_3);
   assign  _net_2378 = (in_do|_reg_3);
   assign  _net_2379 = (in_do|_reg_3);
   assign  _net_2380 = (in_do|_reg_3);
   assign  _net_2381 = (in_do|_reg_3);
   assign  _net_2382 = (in_do|_reg_3);
   assign  _net_2383 = (in_do|_reg_3);
   assign  _net_2384 = (in_do|_reg_3);
   assign  _net_2385 = (in_do|_reg_3);
   assign  _net_2386 = (in_do|_reg_3);
   assign  _net_2387 = (in_do|_reg_3);
   assign  _net_2388 = (in_do|_reg_3);
   assign  _net_2389 = (in_do|_reg_3);
   assign  _net_2390 = (in_do|_reg_3);
   assign  _net_2391 = (in_do|_reg_3);
   assign  _net_2392 = (in_do|_reg_3);
   assign  _net_2393 = (in_do|_reg_3);
   assign  _net_2394 = (in_do|_reg_3);
   assign  _net_2395 = (in_do|_reg_3);
   assign  _net_2396 = (in_do|_reg_3);
   assign  _net_2397 = (in_do|_reg_3);
   assign  _net_2398 = (in_do|_reg_3);
   assign  _net_2399 = (in_do|_reg_3);
   assign  _net_2400 = (in_do|_reg_3);
   assign  _net_2401 = (in_do|_reg_3);
   assign  _net_2402 = (in_do|_reg_3);
   assign  _net_2403 = (in_do|_reg_3);
   assign  _net_2404 = (in_do|_reg_3);
   assign  _net_2405 = (in_do|_reg_3);
   assign  _net_2406 = (in_do|_reg_3);
   assign  _net_2407 = (in_do|_reg_3);
   assign  _net_2408 = (in_do|_reg_3);
   assign  _net_2409 = (in_do|_reg_3);
   assign  _net_2410 = (in_do|_reg_3);
   assign  _net_2411 = (in_do|_reg_3);
   assign  _net_2412 = (in_do|_reg_3);
   assign  _net_2413 = (in_do|_reg_3);
   assign  _net_2414 = (in_do|_reg_3);
   assign  _net_2415 = (in_do|_reg_3);
   assign  _net_2416 = (in_do|_reg_3);
   assign  _net_2417 = (in_do|_reg_3);
   assign  _net_2418 = (in_do|_reg_3);
   assign  _net_2419 = (in_do|_reg_3);
   assign  _net_2420 = (in_do|_reg_3);
   assign  _net_2421 = (in_do|_reg_3);
   assign  _net_2422 = (in_do|_reg_3);
   assign  _net_2423 = (in_do|_reg_3);
   assign  _net_2424 = (in_do|_reg_3);
   assign  _net_2425 = (in_do|_reg_3);
   assign  _net_2426 = (in_do|_reg_3);
   assign  _net_2427 = (in_do|_reg_3);
   assign  _net_2428 = (in_do|_reg_3);
   assign  _net_2429 = (in_do|_reg_3);
   assign  _net_2430 = (in_do|_reg_3);
   assign  _net_2431 = (in_do|_reg_3);
   assign  _net_2432 = (in_do|_reg_3);
   assign  _net_2433 = (in_do|_reg_3);
   assign  _net_2434 = (in_do|_reg_3);
   assign  _net_2435 = (in_do|_reg_3);
   assign  _net_2436 = (in_do|_reg_3);
   assign  _net_2437 = (in_do|_reg_3);
   assign  _net_2438 = (in_do|_reg_3);
   assign  _net_2439 = (in_do|_reg_3);
   assign  _net_2440 = (in_do|_reg_3);
   assign  _net_2441 = (in_do|_reg_3);
   assign  _net_2442 = (in_do|_reg_3);
   assign  _net_2443 = (in_do|_reg_3);
   assign  _net_2444 = (in_do|_reg_3);
   assign  _net_2445 = (in_do|_reg_3);
   assign  _net_2446 = (in_do|_reg_3);
   assign  _net_2447 = (in_do|_reg_3);
   assign  _net_2448 = (in_do|_reg_3);
   assign  _net_2449 = (in_do|_reg_3);
   assign  _net_2450 = (in_do|_reg_3);
   assign  _net_2451 = (in_do|_reg_3);
   assign  _net_2452 = (in_do|_reg_3);
   assign  _net_2453 = (in_do|_reg_3);
   assign  _net_2454 = (in_do|_reg_3);
   assign  _net_2455 = (in_do|_reg_3);
   assign  _net_2456 = (in_do|_reg_3);
   assign  _net_2457 = (in_do|_reg_3);
   assign  _net_2458 = (in_do|_reg_3);
   assign  _net_2459 = (in_do|_reg_3);
   assign  _net_2460 = (in_do|_reg_3);
   assign  _net_2461 = (in_do|_reg_3);
   assign  _net_2462 = (in_do|_reg_3);
   assign  _net_2463 = (in_do|_reg_3);
   assign  _net_2464 = (in_do|_reg_3);
   assign  _net_2465 = (in_do|_reg_3);
   assign  _net_2466 = (in_do|_reg_3);
   assign  _net_2467 = (in_do|_reg_3);
   assign  _net_2468 = (in_do|_reg_3);
   assign  _net_2469 = (in_do|_reg_3);
   assign  _net_2470 = (in_do|_reg_3);
   assign  _net_2471 = (in_do|_reg_3);
   assign  _net_2472 = (in_do|_reg_3);
   assign  _net_2473 = (in_do|_reg_3);
   assign  _net_2474 = (in_do|_reg_3);
   assign  _net_2475 = (in_do|_reg_3);
   assign  _net_2476 = (in_do|_reg_3);
   assign  _net_2477 = (in_do|_reg_3);
   assign  _net_2478 = (in_do|_reg_3);
   assign  _net_2479 = (in_do|_reg_3);
   assign  _net_2480 = (in_do|_reg_3);
   assign  _net_2481 = (in_do|_reg_3);
   assign  _net_2482 = (in_do|_reg_3);
   assign  _net_2483 = (in_do|_reg_3);
   assign  _net_2484 = (in_do|_reg_3);
   assign  _net_2485 = (in_do|_reg_3);
   assign  _net_2486 = (in_do|_reg_3);
   assign  _net_2487 = (in_do|_reg_3);
   assign  _net_2488 = (in_do|_reg_3);
   assign  _net_2489 = (in_do|_reg_3);
   assign  _net_2490 = (in_do|_reg_3);
   assign  _net_2491 = (in_do|_reg_3);
   assign  _net_2492 = (in_do|_reg_3);
   assign  _net_2493 = (in_do|_reg_3);
   assign  _net_2494 = (in_do|_reg_3);
   assign  _net_2495 = (in_do|_reg_3);
   assign  _net_2496 = (in_do|_reg_3);
   assign  _net_2497 = (in_do|_reg_3);
   assign  _net_2498 = (in_do|_reg_3);
   assign  _net_2499 = (in_do|_reg_3);
   assign  _net_2500 = (in_do|_reg_3);
   assign  _net_2501 = (in_do|_reg_3);
   assign  _net_2502 = (in_do|_reg_3);
   assign  _net_2503 = (in_do|_reg_3);
   assign  _net_2504 = (in_do|_reg_3);
   assign  _net_2505 = (in_do|_reg_3);
   assign  _net_2506 = (in_do|_reg_3);
   assign  _net_2507 = (in_do|_reg_3);
   assign  _net_2508 = (in_do|_reg_3);
   assign  _net_2509 = (in_do|_reg_3);
   assign  _net_2510 = (in_do|_reg_3);
   assign  _net_2511 = (in_do|_reg_3);
   assign  _net_2512 = (in_do|_reg_3);
   assign  _net_2513 = (in_do|_reg_3);
   assign  _net_2514 = (in_do|_reg_3);
   assign  _net_2515 = (in_do|_reg_3);
   assign  _net_2516 = (in_do|_reg_3);
   assign  _net_2517 = (in_do|_reg_3);
   assign  _net_2518 = (in_do|_reg_3);
   assign  _net_2519 = (in_do|_reg_3);
   assign  _net_2520 = (in_do|_reg_3);
   assign  _net_2521 = (in_do|_reg_3);
   assign  _net_2522 = (in_do|_reg_3);
   assign  _net_2523 = (in_do|_reg_3);
   assign  _net_2524 = (in_do|_reg_3);
   assign  _net_2525 = (in_do|_reg_3);
   assign  _net_2526 = (in_do|_reg_3);
   assign  _net_2527 = (in_do|_reg_3);
   assign  _net_2528 = (in_do|_reg_3);
   assign  _net_2529 = (in_do|_reg_3);
   assign  _net_2530 = (in_do|_reg_3);
   assign  _net_2531 = (in_do|_reg_3);
   assign  _net_2532 = (in_do|_reg_3);
   assign  _net_2533 = (in_do|_reg_3);
   assign  _net_2534 = (in_do|_reg_3);
   assign  _net_2535 = (in_do|_reg_3);
   assign  _net_2536 = (in_do|_reg_3);
   assign  _net_2537 = (in_do|_reg_3);
   assign  _net_2538 = (in_do|_reg_3);
   assign  _net_2539 = (in_do|_reg_3);
   assign  _net_2540 = (in_do|_reg_3);
   assign  _net_2541 = (in_do|_reg_3);
   assign  _net_2542 = (((_reg_1&_net_4)|in_do)|(_reg_2|_reg_3));
   assign  _net_2543 = (_reg_1|_reg_2);
   assign  _net_2544 = (_reg_0|_reg_1);

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_reg_2545)
    begin
    $display("h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\n",_add_all_x_sg_out33,_add_all_x_sg_out34,_add_all_x_sg_out35,_add_all_x_sg_out36,_add_all_x_sg_out37,_add_all_x_sg_out38,_add_all_x_sg_out39,_add_all_x_sg_out40,_add_all_x_sg_out41,_add_all_x_sg_out42,_add_all_x_sg_out43,_add_all_x_sg_out44,_add_all_x_sg_out45,_add_all_x_sg_out46,_add_all_x_sg_out47,_add_all_x_sg_out48,_add_all_x_sg_out49,_add_all_x_sg_out50,_add_all_x_sg_out51,_add_all_x_sg_out52,_add_all_x_sg_out53,_add_all_x_sg_out54,_add_all_x_sg_out55,_add_all_x_sg_out56,_add_all_x_sg_out57,_add_all_x_sg_out58,_add_all_x_sg_out59,_add_all_x_sg_out60,_add_all_x_sg_out61,_add_all_x_sg_out62,_add_all_x_sg_out65,_add_all_x_sg_out66,_add_all_x_sg_out67,_add_all_x_sg_out68,_add_all_x_sg_out69,_add_all_x_sg_out70,_add_all_x_sg_out71,_add_all_x_sg_out72,_add_all_x_sg_out73,_add_all_x_sg_out74,_add_all_x_sg_out75,_add_all_x_sg_out76,_add_all_x_sg_out77,_add_all_x_sg_out78,_add_all_x_sg_out79,_add_all_x_sg_out80,_add_all_x_sg_out81,_add_all_x_sg_out82,_add_all_x_sg_out83,_add_all_x_sg_out84,_add_all_x_sg_out85,_add_all_x_sg_out86,_add_all_x_sg_out87,_add_all_x_sg_out88,_add_all_x_sg_out89,_add_all_x_sg_out90,_add_all_x_sg_out91,_add_all_x_sg_out92,_add_all_x_sg_out93,_add_all_x_sg_out94,_add_all_x_sg_out97,_add_all_x_sg_out98,_add_all_x_sg_out99,_add_all_x_sg_out100,_add_all_x_sg_out101,_add_all_x_sg_out102,_add_all_x_sg_out103,_add_all_x_sg_out104,_add_all_x_sg_out105,_add_all_x_sg_out106,_add_all_x_sg_out107,_add_all_x_sg_out108,_add_all_x_sg_out109,_add_all_x_sg_out110,_add_all_x_sg_out111,_add_all_x_sg_out112,_add_all_x_sg_out113,_add_all_x_sg_out114,_add_all_x_sg_out115,_add_all_x_sg_out116,_add_all_x_sg_out117,_add_all_x_sg_out118,_add_all_x_sg_out119,_add_all_x_sg_out120,_add_all_x_sg_out121,_add_all_x_sg_out122,_add_all_x_sg_out123,_add_all_x_sg_out124,_add_all_x_sg_out125,_add_all_x_sg_out126,_add_all_x_sg_out129,_add_all_x_sg_out130,_add_all_x_sg_out131,_add_all_x_sg_out132,_add_all_x_sg_out133,_add_all_x_sg_out134,_add_all_x_sg_out135,_add_all_x_sg_out136,_add_all_x_sg_out137,_add_all_x_sg_out138,_add_all_x_sg_out139,_add_all_x_sg_out140,_add_all_x_sg_out141,_add_all_x_sg_out142,_add_all_x_sg_out143,_add_all_x_sg_out144,_add_all_x_sg_out145,_add_all_x_sg_out146,_add_all_x_sg_out147,_add_all_x_sg_out148,_add_all_x_sg_out149,_add_all_x_sg_out150,_add_all_x_sg_out151,_add_all_x_sg_out152,_add_all_x_sg_out153,_add_all_x_sg_out154,_add_all_x_sg_out155,_add_all_x_sg_out156,_add_all_x_sg_out157,_add_all_x_sg_out158,_add_all_x_sg_out161,_add_all_x_sg_out162,_add_all_x_sg_out163,_add_all_x_sg_out164,_add_all_x_sg_out165,_add_all_x_sg_out166,_add_all_x_sg_out167,_add_all_x_sg_out168,_add_all_x_sg_out169,_add_all_x_sg_out170,_add_all_x_sg_out171,_add_all_x_sg_out172,_add_all_x_sg_out173,_add_all_x_sg_out174,_add_all_x_sg_out175,_add_all_x_sg_out176,_add_all_x_sg_out177,_add_all_x_sg_out178,_add_all_x_sg_out179,_add_all_x_sg_out180,_add_all_x_sg_out181,_add_all_x_sg_out182,_add_all_x_sg_out183,_add_all_x_sg_out184,_add_all_x_sg_out185,_add_all_x_sg_out186,_add_all_x_sg_out187,_add_all_x_sg_out188,_add_all_x_sg_out189,_add_all_x_sg_out190,_add_all_x_sg_out193,_add_all_x_sg_out194,_add_all_x_sg_out195,_add_all_x_sg_out196,_add_all_x_sg_out197,_add_all_x_sg_out198,_add_all_x_sg_out199,_add_all_x_sg_out200,_add_all_x_sg_out201,_add_all_x_sg_out202,_add_all_x_sg_out203,_add_all_x_sg_out204,_add_all_x_sg_out205,_add_all_x_sg_out206,_add_all_x_sg_out207,_add_all_x_sg_out208,_add_all_x_sg_out209,_add_all_x_sg_out210,_add_all_x_sg_out211,_add_all_x_sg_out212,_add_all_x_sg_out213,_add_all_x_sg_out214,_add_all_x_sg_out215,_add_all_x_sg_out216,_add_all_x_sg_out217,_add_all_x_sg_out218,_add_all_x_sg_out219,_add_all_x_sg_out220,_add_all_x_sg_out221,_add_all_x_sg_out222,_add_all_x_sg_out225,_add_all_x_sg_out226,_add_all_x_sg_out227,_add_all_x_sg_out228,_add_all_x_sg_out229,_add_all_x_sg_out230,_add_all_x_sg_out231,_add_all_x_sg_out232,_add_all_x_sg_out233,_add_all_x_sg_out234,_add_all_x_sg_out235,_add_all_x_sg_out236,_add_all_x_sg_out237,_add_all_x_sg_out238,_add_all_x_sg_out239,_add_all_x_sg_out240,_add_all_x_sg_out241,_add_all_x_sg_out242,_add_all_x_sg_out243,_add_all_x_sg_out244,_add_all_x_sg_out245,_add_all_x_sg_out246,_add_all_x_sg_out247,_add_all_x_sg_out248,_add_all_x_sg_out249,_add_all_x_sg_out250,_add_all_x_sg_out251,_add_all_x_sg_out252,_add_all_x_sg_out253,_add_all_x_sg_out254,_add_all_x_sg_out257,_add_all_x_sg_out258,_add_all_x_sg_out259,_add_all_x_sg_out260,_add_all_x_sg_out261,_add_all_x_sg_out262,_add_all_x_sg_out263,_add_all_x_sg_out264,_add_all_x_sg_out265,_add_all_x_sg_out266,_add_all_x_sg_out267,_add_all_x_sg_out268,_add_all_x_sg_out269,_add_all_x_sg_out270,_add_all_x_sg_out271,_add_all_x_sg_out272,_add_all_x_sg_out273,_add_all_x_sg_out274,_add_all_x_sg_out275,_add_all_x_sg_out276,_add_all_x_sg_out277,_add_all_x_sg_out278,_add_all_x_sg_out279,_add_all_x_sg_out280,_add_all_x_sg_out281,_add_all_x_sg_out282,_add_all_x_sg_out283,_add_all_x_sg_out284,_add_all_x_sg_out285,_add_all_x_sg_out286,_add_all_x_sg_out289,_add_all_x_sg_out290,_add_all_x_sg_out291,_add_all_x_sg_out292,_add_all_x_sg_out293,_add_all_x_sg_out294,_add_all_x_sg_out295,_add_all_x_sg_out296,_add_all_x_sg_out297,_add_all_x_sg_out298,_add_all_x_sg_out299,_add_all_x_sg_out300,_add_all_x_sg_out301,_add_all_x_sg_out302,_add_all_x_sg_out303,_add_all_x_sg_out304,_add_all_x_sg_out305,_add_all_x_sg_out306,_add_all_x_sg_out307,_add_all_x_sg_out308,_add_all_x_sg_out309,_add_all_x_sg_out310,_add_all_x_sg_out311,_add_all_x_sg_out312,_add_all_x_sg_out313,_add_all_x_sg_out314,_add_all_x_sg_out315,_add_all_x_sg_out316,_add_all_x_sg_out317,_add_all_x_sg_out318,_add_all_x_sg_out321,_add_all_x_sg_out322,_add_all_x_sg_out323,_add_all_x_sg_out324,_add_all_x_sg_out325,_add_all_x_sg_out326,_add_all_x_sg_out327,_add_all_x_sg_out328,_add_all_x_sg_out329,_add_all_x_sg_out330,_add_all_x_sg_out331,_add_all_x_sg_out332,_add_all_x_sg_out333,_add_all_x_sg_out334,_add_all_x_sg_out335,_add_all_x_sg_out336,_add_all_x_sg_out337,_add_all_x_sg_out338,_add_all_x_sg_out339,_add_all_x_sg_out340,_add_all_x_sg_out341,_add_all_x_sg_out342,_add_all_x_sg_out343,_add_all_x_sg_out344,_add_all_x_sg_out345,_add_all_x_sg_out346,_add_all_x_sg_out347,_add_all_x_sg_out348,_add_all_x_sg_out349,_add_all_x_sg_out350,_add_all_x_sg_out353,_add_all_x_sg_out354,_add_all_x_sg_out355,_add_all_x_sg_out356,_add_all_x_sg_out357,_add_all_x_sg_out358,_add_all_x_sg_out359,_add_all_x_sg_out360,_add_all_x_sg_out361,_add_all_x_sg_out362,_add_all_x_sg_out363,_add_all_x_sg_out364,_add_all_x_sg_out365,_add_all_x_sg_out366,_add_all_x_sg_out367,_add_all_x_sg_out368,_add_all_x_sg_out369,_add_all_x_sg_out370,_add_all_x_sg_out371,_add_all_x_sg_out372,_add_all_x_sg_out373,_add_all_x_sg_out374,_add_all_x_sg_out375,_add_all_x_sg_out376,_add_all_x_sg_out377,_add_all_x_sg_out378,_add_all_x_sg_out379,_add_all_x_sg_out380,_add_all_x_sg_out381,_add_all_x_sg_out382,_add_all_x_sg_out385,_add_all_x_sg_out386,_add_all_x_sg_out387,_add_all_x_sg_out388,_add_all_x_sg_out389,_add_all_x_sg_out390,_add_all_x_sg_out391,_add_all_x_sg_out392,_add_all_x_sg_out393,_add_all_x_sg_out394,_add_all_x_sg_out395,_add_all_x_sg_out396,_add_all_x_sg_out397,_add_all_x_sg_out398,_add_all_x_sg_out399,_add_all_x_sg_out400,_add_all_x_sg_out401,_add_all_x_sg_out402,_add_all_x_sg_out403,_add_all_x_sg_out404,_add_all_x_sg_out405,_add_all_x_sg_out406,_add_all_x_sg_out407,_add_all_x_sg_out408,_add_all_x_sg_out409,_add_all_x_sg_out410,_add_all_x_sg_out411,_add_all_x_sg_out412,_add_all_x_sg_out413,_add_all_x_sg_out414,_add_all_x_sg_out417,_add_all_x_sg_out418,_add_all_x_sg_out419,_add_all_x_sg_out420,_add_all_x_sg_out421,_add_all_x_sg_out422,_add_all_x_sg_out423,_add_all_x_sg_out424,_add_all_x_sg_out425,_add_all_x_sg_out426,_add_all_x_sg_out427,_add_all_x_sg_out428,_add_all_x_sg_out429,_add_all_x_sg_out430,_add_all_x_sg_out431,_add_all_x_sg_out432,_add_all_x_sg_out433,_add_all_x_sg_out434,_add_all_x_sg_out435,_add_all_x_sg_out436,_add_all_x_sg_out437,_add_all_x_sg_out438,_add_all_x_sg_out439,_add_all_x_sg_out440,_add_all_x_sg_out441,_add_all_x_sg_out442,_add_all_x_sg_out443,_add_all_x_sg_out444,_add_all_x_sg_out445,_add_all_x_sg_out446,_add_all_x_sg_out449,_add_all_x_sg_out450,_add_all_x_sg_out451,_add_all_x_sg_out452,_add_all_x_sg_out453,_add_all_x_sg_out454,_add_all_x_sg_out455,_add_all_x_sg_out456,_add_all_x_sg_out457,_add_all_x_sg_out458,_add_all_x_sg_out459,_add_all_x_sg_out460,_add_all_x_sg_out461,_add_all_x_sg_out462,_add_all_x_sg_out463,_add_all_x_sg_out464,_add_all_x_sg_out465,_add_all_x_sg_out466,_add_all_x_sg_out467,_add_all_x_sg_out468,_add_all_x_sg_out469,_add_all_x_sg_out470,_add_all_x_sg_out471,_add_all_x_sg_out472,_add_all_x_sg_out473,_add_all_x_sg_out474,_add_all_x_sg_out475,_add_all_x_sg_out476,_add_all_x_sg_out477,_add_all_x_sg_out478);
    end
  end

// synthesis translate_on
// synopsys translate_on

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_reg_2545)
    begin
    $display("h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\nh,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,h,\n",_add_all_x_data_out_index33,_add_all_x_data_out_index34,_add_all_x_data_out_index35,_add_all_x_data_out_index36,_add_all_x_data_out_index37,_add_all_x_data_out_index38,_add_all_x_data_out_index39,_add_all_x_data_out_index40,_add_all_x_data_out_index41,_add_all_x_data_out_index42,_add_all_x_data_out_index43,_add_all_x_data_out_index44,_add_all_x_data_out_index45,_add_all_x_data_out_index46,_add_all_x_data_out_index47,_add_all_x_data_out_index48,_add_all_x_data_out_index49,_add_all_x_data_out_index50,_add_all_x_data_out_index51,_add_all_x_data_out_index52,_add_all_x_data_out_index53,_add_all_x_data_out_index54,_add_all_x_data_out_index55,_add_all_x_data_out_index56,_add_all_x_data_out_index57,_add_all_x_data_out_index58,_add_all_x_data_out_index59,_add_all_x_data_out_index60,_add_all_x_data_out_index61,_add_all_x_data_out_index62,_add_all_x_data_out_index65,_add_all_x_data_out_index66,_add_all_x_data_out_index67,_add_all_x_data_out_index68,_add_all_x_data_out_index69,_add_all_x_data_out_index70,_add_all_x_data_out_index71,_add_all_x_data_out_index72,_add_all_x_data_out_index73,_add_all_x_data_out_index74,_add_all_x_data_out_index75,_add_all_x_data_out_index76,_add_all_x_data_out_index77,_add_all_x_data_out_index78,_add_all_x_data_out_index79,_add_all_x_data_out_index80,_add_all_x_data_out_index81,_add_all_x_data_out_index82,_add_all_x_data_out_index83,_add_all_x_data_out_index84,_add_all_x_data_out_index85,_add_all_x_data_out_index86,_add_all_x_data_out_index87,_add_all_x_data_out_index88,_add_all_x_data_out_index89,_add_all_x_data_out_index90,_add_all_x_data_out_index91,_add_all_x_data_out_index92,_add_all_x_data_out_index93,_add_all_x_data_out_index94,_add_all_x_data_out_index97,_add_all_x_data_out_index98,_add_all_x_data_out_index99,_add_all_x_data_out_index100,_add_all_x_data_out_index101,_add_all_x_data_out_index102,_add_all_x_data_out_index103,_add_all_x_data_out_index104,_add_all_x_data_out_index105,_add_all_x_data_out_index106,_add_all_x_data_out_index107,_add_all_x_data_out_index108,_add_all_x_data_out_index109,_add_all_x_data_out_index110,_add_all_x_data_out_index111,_add_all_x_data_out_index112,_add_all_x_data_out_index113,_add_all_x_data_out_index114,_add_all_x_data_out_index115,_add_all_x_data_out_index116,_add_all_x_data_out_index117,_add_all_x_data_out_index118,_add_all_x_data_out_index119,_add_all_x_data_out_index120,_add_all_x_data_out_index121,_add_all_x_data_out_index122,_add_all_x_data_out_index123,_add_all_x_data_out_index124,_add_all_x_data_out_index125,_add_all_x_data_out_index126,_add_all_x_data_out_index129,_add_all_x_data_out_index130,_add_all_x_data_out_index131,_add_all_x_data_out_index132,_add_all_x_data_out_index133,_add_all_x_data_out_index134,_add_all_x_data_out_index135,_add_all_x_data_out_index136,_add_all_x_data_out_index137,_add_all_x_data_out_index138,_add_all_x_data_out_index139,_add_all_x_data_out_index140,_add_all_x_data_out_index141,_add_all_x_data_out_index142,_add_all_x_data_out_index143,_add_all_x_data_out_index144,_add_all_x_data_out_index145,_add_all_x_data_out_index146,_add_all_x_data_out_index147,_add_all_x_data_out_index148,_add_all_x_data_out_index149,_add_all_x_data_out_index150,_add_all_x_data_out_index151,_add_all_x_data_out_index152,_add_all_x_data_out_index153,_add_all_x_data_out_index154,_add_all_x_data_out_index155,_add_all_x_data_out_index156,_add_all_x_data_out_index157,_add_all_x_data_out_index158,_add_all_x_data_out_index161,_add_all_x_data_out_index162,_add_all_x_data_out_index163,_add_all_x_data_out_index164,_add_all_x_data_out_index165,_add_all_x_data_out_index166,_add_all_x_data_out_index167,_add_all_x_data_out_index168,_add_all_x_data_out_index169,_add_all_x_data_out_index170,_add_all_x_data_out_index171,_add_all_x_data_out_index172,_add_all_x_data_out_index173,_add_all_x_data_out_index174,_add_all_x_data_out_index175,_add_all_x_data_out_index176,_add_all_x_data_out_index177,_add_all_x_data_out_index178,_add_all_x_data_out_index179,_add_all_x_data_out_index180,_add_all_x_data_out_index181,_add_all_x_data_out_index182,_add_all_x_data_out_index183,_add_all_x_data_out_index184,_add_all_x_data_out_index185,_add_all_x_data_out_index186,_add_all_x_data_out_index187,_add_all_x_data_out_index188,_add_all_x_data_out_index189,_add_all_x_data_out_index190,_add_all_x_data_out_index193,_add_all_x_data_out_index194,_add_all_x_data_out_index195,_add_all_x_data_out_index196,_add_all_x_data_out_index197,_add_all_x_data_out_index198,_add_all_x_data_out_index199,_add_all_x_data_out_index200,_add_all_x_data_out_index201,_add_all_x_data_out_index202,_add_all_x_data_out_index203,_add_all_x_data_out_index204,_add_all_x_data_out_index205,_add_all_x_data_out_index206,_add_all_x_data_out_index207,_add_all_x_data_out_index208,_add_all_x_data_out_index209,_add_all_x_data_out_index210,_add_all_x_data_out_index211,_add_all_x_data_out_index212,_add_all_x_data_out_index213,_add_all_x_data_out_index214,_add_all_x_data_out_index215,_add_all_x_data_out_index216,_add_all_x_data_out_index217,_add_all_x_data_out_index218,_add_all_x_data_out_index219,_add_all_x_data_out_index220,_add_all_x_data_out_index221,_add_all_x_data_out_index222,_add_all_x_data_out_index225,_add_all_x_data_out_index226,_add_all_x_data_out_index227,_add_all_x_data_out_index228,_add_all_x_data_out_index229,_add_all_x_data_out_index230,_add_all_x_data_out_index231,_add_all_x_data_out_index232,_add_all_x_data_out_index233,_add_all_x_data_out_index234,_add_all_x_data_out_index235,_add_all_x_data_out_index236,_add_all_x_data_out_index237,_add_all_x_data_out_index238,_add_all_x_data_out_index239,_add_all_x_data_out_index240,_add_all_x_data_out_index241,_add_all_x_data_out_index242,_add_all_x_data_out_index243,_add_all_x_data_out_index244,_add_all_x_data_out_index245,_add_all_x_data_out_index246,_add_all_x_data_out_index247,_add_all_x_data_out_index248,_add_all_x_data_out_index249,_add_all_x_data_out_index250,_add_all_x_data_out_index251,_add_all_x_data_out_index252,_add_all_x_data_out_index253,_add_all_x_data_out_index254,_add_all_x_data_out_index257,_add_all_x_data_out_index258,_add_all_x_data_out_index259,_add_all_x_data_out_index260,_add_all_x_data_out_index261,_add_all_x_data_out_index262,_add_all_x_data_out_index263,_add_all_x_data_out_index264,_add_all_x_data_out_index265,_add_all_x_data_out_index266,_add_all_x_data_out_index267,_add_all_x_data_out_index268,_add_all_x_data_out_index269,_add_all_x_data_out_index270,_add_all_x_data_out_index271,_add_all_x_data_out_index272,_add_all_x_data_out_index273,_add_all_x_data_out_index274,_add_all_x_data_out_index275,_add_all_x_data_out_index276,_add_all_x_data_out_index277,_add_all_x_data_out_index278,_add_all_x_data_out_index279,_add_all_x_data_out_index280,_add_all_x_data_out_index281,_add_all_x_data_out_index282,_add_all_x_data_out_index283,_add_all_x_data_out_index284,_add_all_x_data_out_index285,_add_all_x_data_out_index286,_add_all_x_data_out_index289,_add_all_x_data_out_index290,_add_all_x_data_out_index291,_add_all_x_data_out_index292,_add_all_x_data_out_index293,_add_all_x_data_out_index294,_add_all_x_data_out_index295,_add_all_x_data_out_index296,_add_all_x_data_out_index297,_add_all_x_data_out_index298,_add_all_x_data_out_index299,_add_all_x_data_out_index300,_add_all_x_data_out_index301,_add_all_x_data_out_index302,_add_all_x_data_out_index303,_add_all_x_data_out_index304,_add_all_x_data_out_index305,_add_all_x_data_out_index306,_add_all_x_data_out_index307,_add_all_x_data_out_index308,_add_all_x_data_out_index309,_add_all_x_data_out_index310,_add_all_x_data_out_index311,_add_all_x_data_out_index312,_add_all_x_data_out_index313,_add_all_x_data_out_index314,_add_all_x_data_out_index315,_add_all_x_data_out_index316,_add_all_x_data_out_index317,_add_all_x_data_out_index318,_add_all_x_data_out_index321,_add_all_x_data_out_index322,_add_all_x_data_out_index323,_add_all_x_data_out_index324,_add_all_x_data_out_index325,_add_all_x_data_out_index326,_add_all_x_data_out_index327,_add_all_x_data_out_index328,_add_all_x_data_out_index329,_add_all_x_data_out_index330,_add_all_x_data_out_index331,_add_all_x_data_out_index332,_add_all_x_data_out_index333,_add_all_x_data_out_index334,_add_all_x_data_out_index335,_add_all_x_data_out_index336,_add_all_x_data_out_index337,_add_all_x_data_out_index338,_add_all_x_data_out_index339,_add_all_x_data_out_index340,_add_all_x_data_out_index341,_add_all_x_data_out_index342,_add_all_x_data_out_index343,_add_all_x_data_out_index344,_add_all_x_data_out_index345,_add_all_x_data_out_index346,_add_all_x_data_out_index347,_add_all_x_data_out_index348,_add_all_x_data_out_index349,_add_all_x_data_out_index350,_add_all_x_data_out_index353,_add_all_x_data_out_index354,_add_all_x_data_out_index355,_add_all_x_data_out_index356,_add_all_x_data_out_index357,_add_all_x_data_out_index358,_add_all_x_data_out_index359,_add_all_x_data_out_index360,_add_all_x_data_out_index361,_add_all_x_data_out_index362,_add_all_x_data_out_index363,_add_all_x_data_out_index364,_add_all_x_data_out_index365,_add_all_x_data_out_index366,_add_all_x_data_out_index367,_add_all_x_data_out_index368,_add_all_x_data_out_index369,_add_all_x_data_out_index370,_add_all_x_data_out_index371,_add_all_x_data_out_index372,_add_all_x_data_out_index373,_add_all_x_data_out_index374,_add_all_x_data_out_index375,_add_all_x_data_out_index376,_add_all_x_data_out_index377,_add_all_x_data_out_index378,_add_all_x_data_out_index379,_add_all_x_data_out_index380,_add_all_x_data_out_index381,_add_all_x_data_out_index382,_add_all_x_data_out_index385,_add_all_x_data_out_index386,_add_all_x_data_out_index387,_add_all_x_data_out_index388,_add_all_x_data_out_index389,_add_all_x_data_out_index390,_add_all_x_data_out_index391,_add_all_x_data_out_index392,_add_all_x_data_out_index393,_add_all_x_data_out_index394,_add_all_x_data_out_index395,_add_all_x_data_out_index396,_add_all_x_data_out_index397,_add_all_x_data_out_index398,_add_all_x_data_out_index399,_add_all_x_data_out_index400,_add_all_x_data_out_index401,_add_all_x_data_out_index402,_add_all_x_data_out_index403,_add_all_x_data_out_index404,_add_all_x_data_out_index405,_add_all_x_data_out_index406,_add_all_x_data_out_index407,_add_all_x_data_out_index408,_add_all_x_data_out_index409,_add_all_x_data_out_index410,_add_all_x_data_out_index411,_add_all_x_data_out_index412,_add_all_x_data_out_index413,_add_all_x_data_out_index414,_add_all_x_data_out_index417,_add_all_x_data_out_index418,_add_all_x_data_out_index419,_add_all_x_data_out_index420,_add_all_x_data_out_index421,_add_all_x_data_out_index422,_add_all_x_data_out_index423,_add_all_x_data_out_index424,_add_all_x_data_out_index425,_add_all_x_data_out_index426,_add_all_x_data_out_index427,_add_all_x_data_out_index428,_add_all_x_data_out_index429,_add_all_x_data_out_index430,_add_all_x_data_out_index431,_add_all_x_data_out_index432,_add_all_x_data_out_index433,_add_all_x_data_out_index434,_add_all_x_data_out_index435,_add_all_x_data_out_index436,_add_all_x_data_out_index437,_add_all_x_data_out_index438,_add_all_x_data_out_index439,_add_all_x_data_out_index440,_add_all_x_data_out_index441,_add_all_x_data_out_index442,_add_all_x_data_out_index443,_add_all_x_data_out_index444,_add_all_x_data_out_index445,_add_all_x_data_out_index446,_add_all_x_data_out_index449,_add_all_x_data_out_index450,_add_all_x_data_out_index451,_add_all_x_data_out_index452,_add_all_x_data_out_index453,_add_all_x_data_out_index454,_add_all_x_data_out_index455,_add_all_x_data_out_index456,_add_all_x_data_out_index457,_add_all_x_data_out_index458,_add_all_x_data_out_index459,_add_all_x_data_out_index460,_add_all_x_data_out_index461,_add_all_x_data_out_index462,_add_all_x_data_out_index463,_add_all_x_data_out_index464,_add_all_x_data_out_index465,_add_all_x_data_out_index466,_add_all_x_data_out_index467,_add_all_x_data_out_index468,_add_all_x_data_out_index469,_add_all_x_data_out_index470,_add_all_x_data_out_index471,_add_all_x_data_out_index472,_add_all_x_data_out_index473,_add_all_x_data_out_index474,_add_all_x_data_out_index475,_add_all_x_data_out_index476,_add_all_x_data_out_index477,_add_all_x_data_out_index478);
    end
  end

// synthesis translate_on
// synopsys translate_on
   assign  _net_2549 = (~even);
   assign  _net_2550 = (_reg_2545&_net_2549);
   assign  _net_2551 = (_reg_2545&_net_2549);
   assign  _net_2552 = (_reg_2545&_net_2549);
   assign  _net_2553 = (_reg_2545&_net_2549);
   assign  _net_2554 = (_reg_2545&_net_2549);
   assign  _net_2555 = (_reg_2545&_net_2549);
   assign  _net_2556 = (_reg_2545&_net_2549);
   assign  _net_2557 = (_reg_2545&_net_2549);
   assign  _net_2558 = (_reg_2545&_net_2549);
   assign  _net_2559 = (_reg_2545&_net_2549);
   assign  _net_2560 = (_reg_2545&_net_2549);
   assign  _net_2561 = (_reg_2545&_net_2549);
   assign  _net_2562 = (_reg_2545&_net_2549);
   assign  _net_2563 = (_reg_2545&_net_2549);
   assign  _net_2564 = (_reg_2545&_net_2549);
   assign  _net_2565 = (_reg_2545&_net_2549);
   assign  _net_2566 = (_reg_2545&_net_2549);
   assign  _net_2567 = (_reg_2545&_net_2549);
   assign  _net_2568 = (_reg_2545&_net_2549);
   assign  _net_2569 = (_reg_2545&_net_2549);
   assign  _net_2570 = (_reg_2545&_net_2549);
   assign  _net_2571 = (_reg_2545&_net_2549);
   assign  _net_2572 = (_reg_2545&_net_2549);
   assign  _net_2573 = (_reg_2545&_net_2549);
   assign  _net_2574 = (_reg_2545&_net_2549);
   assign  _net_2575 = (_reg_2545&_net_2549);
   assign  _net_2576 = (_reg_2545&_net_2549);
   assign  _net_2577 = (_reg_2545&_net_2549);
   assign  _net_2578 = (_reg_2545&_net_2549);
   assign  _net_2579 = (_reg_2545&_net_2549);
   assign  _net_2580 = (_reg_2545&_net_2549);
   assign  _net_2581 = (_reg_2545&_net_2549);
   assign  _net_2582 = (_reg_2545&_net_2549);
   assign  _net_2583 = (_reg_2545&_net_2549);
   assign  _net_2584 = (_reg_2545&_net_2549);
   assign  _net_2585 = (_reg_2545&_net_2549);
   assign  _net_2586 = (_reg_2545&_net_2549);
   assign  _net_2587 = (_reg_2545&_net_2549);
   assign  _net_2588 = (_reg_2545&_net_2549);
   assign  _net_2589 = (_reg_2545&_net_2549);
   assign  _net_2590 = (_reg_2545&_net_2549);
   assign  _net_2591 = (_reg_2545&_net_2549);
   assign  _net_2592 = (_reg_2545&_net_2549);
   assign  _net_2593 = (_reg_2545&_net_2549);
   assign  _net_2594 = (_reg_2545&_net_2549);
   assign  _net_2595 = (_reg_2545&_net_2549);
   assign  _net_2596 = (_reg_2545&_net_2549);
   assign  _net_2597 = (_reg_2545&_net_2549);
   assign  _net_2598 = (_reg_2545&_net_2549);
   assign  _net_2599 = (_reg_2545&_net_2549);
   assign  _net_2600 = (_reg_2545&_net_2549);
   assign  _net_2601 = (_reg_2545&_net_2549);
   assign  _net_2602 = (_reg_2545&_net_2549);
   assign  _net_2603 = (_reg_2545&_net_2549);
   assign  _net_2604 = (_reg_2545&_net_2549);
   assign  _net_2605 = (_reg_2545&_net_2549);
   assign  _net_2606 = (_reg_2545&_net_2549);
   assign  _net_2607 = (_reg_2545&_net_2549);
   assign  _net_2608 = (_reg_2545&_net_2549);
   assign  _net_2609 = (_reg_2545&_net_2549);
   assign  _net_2610 = (_reg_2545&_net_2549);
   assign  _net_2611 = (_reg_2545&_net_2549);
   assign  _net_2612 = (_reg_2545&_net_2549);
   assign  _net_2613 = (_reg_2545&_net_2549);
   assign  _net_2614 = (_reg_2545&_net_2549);
   assign  _net_2615 = (_reg_2545&_net_2549);
   assign  _net_2616 = (_reg_2545&_net_2549);
   assign  _net_2617 = (_reg_2545&_net_2549);
   assign  _net_2618 = (_reg_2545&_net_2549);
   assign  _net_2619 = (_reg_2545&_net_2549);
   assign  _net_2620 = (_reg_2545&_net_2549);
   assign  _net_2621 = (_reg_2545&_net_2549);
   assign  _net_2622 = (_reg_2545&_net_2549);
   assign  _net_2623 = (_reg_2545&_net_2549);
   assign  _net_2624 = (_reg_2545&_net_2549);
   assign  _net_2625 = (_reg_2545&_net_2549);
   assign  _net_2626 = (_reg_2545&_net_2549);
   assign  _net_2627 = (_reg_2545&_net_2549);
   assign  _net_2628 = (_reg_2545&_net_2549);
   assign  _net_2629 = (_reg_2545&_net_2549);
   assign  _net_2630 = (_reg_2545&_net_2549);
   assign  _net_2631 = (_reg_2545&_net_2549);
   assign  _net_2632 = (_reg_2545&_net_2549);
   assign  _net_2633 = (_reg_2545&_net_2549);
   assign  _net_2634 = (_reg_2545&_net_2549);
   assign  _net_2635 = (_reg_2545&_net_2549);
   assign  _net_2636 = (_reg_2545&_net_2549);
   assign  _net_2637 = (_reg_2545&_net_2549);
   assign  _net_2638 = (_reg_2545&_net_2549);
   assign  _net_2639 = (_reg_2545&_net_2549);
   assign  _net_2640 = (_reg_2545&_net_2549);
   assign  _net_2641 = (_reg_2545&_net_2549);
   assign  _net_2642 = (_reg_2545&_net_2549);
   assign  _net_2643 = (_reg_2545&_net_2549);
   assign  _net_2644 = (_reg_2545&_net_2549);
   assign  _net_2645 = (_reg_2545&_net_2549);
   assign  _net_2646 = (_reg_2545&_net_2549);
   assign  _net_2647 = (_reg_2545&_net_2549);
   assign  _net_2648 = (_reg_2545&_net_2549);
   assign  _net_2649 = (_reg_2545&_net_2549);
   assign  _net_2650 = (_reg_2545&_net_2549);
   assign  _net_2651 = (_reg_2545&_net_2549);
   assign  _net_2652 = (_reg_2545&_net_2549);
   assign  _net_2653 = (_reg_2545&_net_2549);
   assign  _net_2654 = (_reg_2545&_net_2549);
   assign  _net_2655 = (_reg_2545&_net_2549);
   assign  _net_2656 = (_reg_2545&_net_2549);
   assign  _net_2657 = (_reg_2545&_net_2549);
   assign  _net_2658 = (_reg_2545&_net_2549);
   assign  _net_2659 = (_reg_2545&_net_2549);
   assign  _net_2660 = (_reg_2545&_net_2549);
   assign  _net_2661 = (_reg_2545&_net_2549);
   assign  _net_2662 = (_reg_2545&_net_2549);
   assign  _net_2663 = (_reg_2545&_net_2549);
   assign  _net_2664 = (_reg_2545&_net_2549);
   assign  _net_2665 = (_reg_2545&_net_2549);
   assign  _net_2666 = (_reg_2545&_net_2549);
   assign  _net_2667 = (_reg_2545&_net_2549);
   assign  _net_2668 = (_reg_2545&_net_2549);
   assign  _net_2669 = (_reg_2545&_net_2549);
   assign  _net_2670 = (_reg_2545&_net_2549);
   assign  _net_2671 = (_reg_2545&_net_2549);
   assign  _net_2672 = (_reg_2545&_net_2549);
   assign  _net_2673 = (_reg_2545&_net_2549);
   assign  _net_2674 = (_reg_2545&_net_2549);
   assign  _net_2675 = (_reg_2545&_net_2549);
   assign  _net_2676 = (_reg_2545&_net_2549);
   assign  _net_2677 = (_reg_2545&_net_2549);
   assign  _net_2678 = (_reg_2545&_net_2549);
   assign  _net_2679 = (_reg_2545&_net_2549);
   assign  _net_2680 = (_reg_2545&_net_2549);
   assign  _net_2681 = (_reg_2545&_net_2549);
   assign  _net_2682 = (_reg_2545&_net_2549);
   assign  _net_2683 = (_reg_2545&_net_2549);
   assign  _net_2684 = (_reg_2545&_net_2549);
   assign  _net_2685 = (_reg_2545&_net_2549);
   assign  _net_2686 = (_reg_2545&_net_2549);
   assign  _net_2687 = (_reg_2545&_net_2549);
   assign  _net_2688 = (_reg_2545&_net_2549);
   assign  _net_2689 = (_reg_2545&_net_2549);
   assign  _net_2690 = (_reg_2545&_net_2549);
   assign  _net_2691 = (_reg_2545&_net_2549);
   assign  _net_2692 = (_reg_2545&_net_2549);
   assign  _net_2693 = (_reg_2545&_net_2549);
   assign  _net_2694 = (_reg_2545&_net_2549);
   assign  _net_2695 = (_reg_2545&_net_2549);
   assign  _net_2696 = (_reg_2545&_net_2549);
   assign  _net_2697 = (_reg_2545&_net_2549);
   assign  _net_2698 = (_reg_2545&_net_2549);
   assign  _net_2699 = (_reg_2545&_net_2549);
   assign  _net_2700 = (_reg_2545&_net_2549);
   assign  _net_2701 = (_reg_2545&_net_2549);
   assign  _net_2702 = (_reg_2545&_net_2549);
   assign  _net_2703 = (_reg_2545&_net_2549);
   assign  _net_2704 = (_reg_2545&_net_2549);
   assign  _net_2705 = (_reg_2545&_net_2549);
   assign  _net_2706 = (_reg_2545&_net_2549);
   assign  _net_2707 = (_reg_2545&_net_2549);
   assign  _net_2708 = (_reg_2545&_net_2549);
   assign  _net_2709 = (_reg_2545&_net_2549);
   assign  _net_2710 = (_reg_2545&_net_2549);
   assign  _net_2711 = (_reg_2545&_net_2549);
   assign  _net_2712 = (_reg_2545&_net_2549);
   assign  _net_2713 = (_reg_2545&_net_2549);
   assign  _net_2714 = (_reg_2545&_net_2549);
   assign  _net_2715 = (_reg_2545&_net_2549);
   assign  _net_2716 = (_reg_2545&_net_2549);
   assign  _net_2717 = (_reg_2545&_net_2549);
   assign  _net_2718 = (_reg_2545&_net_2549);
   assign  _net_2719 = (_reg_2545&_net_2549);
   assign  _net_2720 = (_reg_2545&_net_2549);
   assign  _net_2721 = (_reg_2545&_net_2549);
   assign  _net_2722 = (_reg_2545&_net_2549);
   assign  _net_2723 = (_reg_2545&_net_2549);
   assign  _net_2724 = (_reg_2545&_net_2549);
   assign  _net_2725 = (_reg_2545&_net_2549);
   assign  _net_2726 = (_reg_2545&_net_2549);
   assign  _net_2727 = (_reg_2545&_net_2549);
   assign  _net_2728 = (_reg_2545&_net_2549);
   assign  _net_2729 = (_reg_2545&_net_2549);
   assign  _net_2730 = (_reg_2545&_net_2549);
   assign  _net_2731 = (_reg_2545&_net_2549);
   assign  _net_2732 = (_reg_2545&_net_2549);
   assign  _net_2733 = (_reg_2545&_net_2549);
   assign  _net_2734 = (_reg_2545&_net_2549);
   assign  _net_2735 = (_reg_2545&_net_2549);
   assign  _net_2736 = (_reg_2545&_net_2549);
   assign  _net_2737 = (_reg_2545&_net_2549);
   assign  _net_2738 = (_reg_2545&_net_2549);
   assign  _net_2739 = (_reg_2545&_net_2549);
   assign  _net_2740 = (_reg_2545&_net_2549);
   assign  _net_2741 = (_reg_2545&_net_2549);
   assign  _net_2742 = (_reg_2545&_net_2549);
   assign  _net_2743 = (_reg_2545&_net_2549);
   assign  _net_2744 = (_reg_2545&_net_2549);
   assign  _net_2745 = (_reg_2545&_net_2549);
   assign  _net_2746 = (_reg_2545&_net_2549);
   assign  _net_2747 = (_reg_2545&_net_2549);
   assign  _net_2748 = (_reg_2545&_net_2549);
   assign  _net_2749 = (_reg_2545&_net_2549);
   assign  _net_2750 = (_reg_2545&_net_2549);
   assign  _net_2751 = (_reg_2545&_net_2549);
   assign  _net_2752 = (_reg_2545&_net_2549);
   assign  _net_2753 = (_reg_2545&_net_2549);
   assign  _net_2754 = (_reg_2545&_net_2549);
   assign  _net_2755 = (_reg_2545&_net_2549);
   assign  _net_2756 = (_reg_2545&_net_2549);
   assign  _net_2757 = (_reg_2545&_net_2549);
   assign  _net_2758 = (_reg_2545&_net_2549);
   assign  _net_2759 = (_reg_2545&_net_2549);
   assign  _net_2760 = (_reg_2545&_net_2549);
   assign  _net_2761 = (_reg_2545&_net_2549);
   assign  _net_2762 = (_reg_2545&_net_2549);
   assign  _net_2763 = (_reg_2545&_net_2549);
   assign  _net_2764 = (_reg_2545&_net_2549);
   assign  _net_2765 = (_reg_2545&_net_2549);
   assign  _net_2766 = (_reg_2545&_net_2549);
   assign  _net_2767 = (_reg_2545&_net_2549);
   assign  _net_2768 = (_reg_2545&_net_2549);
   assign  _net_2769 = (_reg_2545&_net_2549);
   assign  _net_2770 = (_reg_2545&_net_2549);
   assign  _net_2771 = (_reg_2545&_net_2549);
   assign  _net_2772 = (_reg_2545&_net_2549);
   assign  _net_2773 = (_reg_2545&_net_2549);
   assign  _net_2774 = (_reg_2545&_net_2549);
   assign  _net_2775 = (_reg_2545&_net_2549);
   assign  _net_2776 = (_reg_2545&_net_2549);
   assign  _net_2777 = (_reg_2545&_net_2549);
   assign  _net_2778 = (_reg_2545&_net_2549);
   assign  _net_2779 = (_reg_2545&_net_2549);
   assign  _net_2780 = (_reg_2545&_net_2549);
   assign  _net_2781 = (_reg_2545&_net_2549);
   assign  _net_2782 = (_reg_2545&_net_2549);
   assign  _net_2783 = (_reg_2545&_net_2549);
   assign  _net_2784 = (_reg_2545&_net_2549);
   assign  _net_2785 = (_reg_2545&_net_2549);
   assign  _net_2786 = (_reg_2545&_net_2549);
   assign  _net_2787 = (_reg_2545&_net_2549);
   assign  _net_2788 = (_reg_2545&_net_2549);
   assign  _net_2789 = (_reg_2545&_net_2549);
   assign  _net_2790 = (_reg_2545&_net_2549);
   assign  _net_2791 = (_reg_2545&_net_2549);
   assign  _net_2792 = (_reg_2545&_net_2549);
   assign  _net_2793 = (_reg_2545&_net_2549);
   assign  _net_2794 = (_reg_2545&_net_2549);
   assign  _net_2795 = (_reg_2545&_net_2549);
   assign  _net_2796 = (_reg_2545&_net_2549);
   assign  _net_2797 = (_reg_2545&_net_2549);
   assign  _net_2798 = (_reg_2545&_net_2549);
   assign  _net_2799 = (_reg_2545&_net_2549);
   assign  _net_2800 = (_reg_2545&_net_2549);
   assign  _net_2801 = (_reg_2545&_net_2549);
   assign  _net_2802 = (_reg_2545&_net_2549);
   assign  _net_2803 = (_reg_2545&_net_2549);
   assign  _net_2804 = (_reg_2545&_net_2549);
   assign  _net_2805 = (_reg_2545&_net_2549);
   assign  _net_2806 = (_reg_2545&_net_2549);
   assign  _net_2807 = (_reg_2545&_net_2549);
   assign  _net_2808 = (_reg_2545&_net_2549);
   assign  _net_2809 = (_reg_2545&_net_2549);
   assign  _net_2810 = (_reg_2545&_net_2549);
   assign  _net_2811 = (_reg_2545&_net_2549);
   assign  _net_2812 = (_reg_2545&_net_2549);
   assign  _net_2813 = (_reg_2545&_net_2549);
   assign  _net_2814 = (_reg_2545&_net_2549);
   assign  _net_2815 = (_reg_2545&_net_2549);
   assign  _net_2816 = (_reg_2545&_net_2549);
   assign  _net_2817 = (_reg_2545&_net_2549);
   assign  _net_2818 = (_reg_2545&_net_2549);
   assign  _net_2819 = (_reg_2545&_net_2549);
   assign  _net_2820 = (_reg_2545&_net_2549);
   assign  _net_2821 = (_reg_2545&_net_2549);
   assign  _net_2822 = (_reg_2545&_net_2549);
   assign  _net_2823 = (_reg_2545&_net_2549);
   assign  _net_2824 = (_reg_2545&_net_2549);
   assign  _net_2825 = (_reg_2545&_net_2549);
   assign  _net_2826 = (_reg_2545&_net_2549);
   assign  _net_2827 = (_reg_2545&_net_2549);
   assign  _net_2828 = (_reg_2545&_net_2549);
   assign  _net_2829 = (_reg_2545&_net_2549);
   assign  _net_2830 = (_reg_2545&_net_2549);
   assign  _net_2831 = (_reg_2545&_net_2549);
   assign  _net_2832 = (_reg_2545&_net_2549);
   assign  _net_2833 = (_reg_2545&_net_2549);
   assign  _net_2834 = (_reg_2545&_net_2549);
   assign  _net_2835 = (_reg_2545&_net_2549);
   assign  _net_2836 = (_reg_2545&_net_2549);
   assign  _net_2837 = (_reg_2545&_net_2549);
   assign  _net_2838 = (_reg_2545&_net_2549);
   assign  _net_2839 = (_reg_2545&_net_2549);
   assign  _net_2840 = (_reg_2545&_net_2549);
   assign  _net_2841 = (_reg_2545&_net_2549);
   assign  _net_2842 = (_reg_2545&_net_2549);
   assign  _net_2843 = (_reg_2545&_net_2549);
   assign  _net_2844 = (_reg_2545&_net_2549);
   assign  _net_2845 = (_reg_2545&_net_2549);
   assign  _net_2846 = (_reg_2545&_net_2549);
   assign  _net_2847 = (_reg_2545&_net_2549);
   assign  _net_2848 = (_reg_2545&_net_2549);
   assign  _net_2849 = (_reg_2545&_net_2549);
   assign  _net_2850 = (_reg_2545&_net_2549);
   assign  _net_2851 = (_reg_2545&_net_2549);
   assign  _net_2852 = (_reg_2545&_net_2549);
   assign  _net_2853 = (_reg_2545&_net_2549);
   assign  _net_2854 = (_reg_2545&_net_2549);
   assign  _net_2855 = (_reg_2545&_net_2549);
   assign  _net_2856 = (_reg_2545&_net_2549);
   assign  _net_2857 = (_reg_2545&_net_2549);
   assign  _net_2858 = (_reg_2545&_net_2549);
   assign  _net_2859 = (_reg_2545&_net_2549);
   assign  _net_2860 = (_reg_2545&_net_2549);
   assign  _net_2861 = (_reg_2545&_net_2549);
   assign  _net_2862 = (_reg_2545&_net_2549);
   assign  _net_2863 = (_reg_2545&_net_2549);
   assign  _net_2864 = (_reg_2545&_net_2549);
   assign  _net_2865 = (_reg_2545&_net_2549);
   assign  _net_2866 = (_reg_2545&_net_2549);
   assign  _net_2867 = (_reg_2545&_net_2549);
   assign  _net_2868 = (_reg_2545&_net_2549);
   assign  _net_2869 = (_reg_2545&_net_2549);
   assign  _net_2870 = (_reg_2545&_net_2549);
   assign  _net_2871 = (_reg_2545&_net_2549);
   assign  _net_2872 = (_reg_2545&_net_2549);
   assign  _net_2873 = (_reg_2545&_net_2549);
   assign  _net_2874 = (_reg_2545&_net_2549);
   assign  _net_2875 = (_reg_2545&_net_2549);
   assign  _net_2876 = (_reg_2545&_net_2549);
   assign  _net_2877 = (_reg_2545&_net_2549);
   assign  _net_2878 = (_reg_2545&_net_2549);
   assign  _net_2879 = (_reg_2545&_net_2549);
   assign  _net_2880 = (_reg_2545&_net_2549);
   assign  _net_2881 = (_reg_2545&_net_2549);
   assign  _net_2882 = (_reg_2545&_net_2549);
   assign  _net_2883 = (_reg_2545&_net_2549);
   assign  _net_2884 = (_reg_2545&_net_2549);
   assign  _net_2885 = (_reg_2545&_net_2549);
   assign  _net_2886 = (_reg_2545&_net_2549);
   assign  _net_2887 = (_reg_2545&_net_2549);
   assign  _net_2888 = (_reg_2545&_net_2549);
   assign  _net_2889 = (_reg_2545&_net_2549);
   assign  _net_2890 = (_reg_2545&_net_2549);
   assign  _net_2891 = (_reg_2545&_net_2549);
   assign  _net_2892 = (_reg_2545&_net_2549);
   assign  _net_2893 = (_reg_2545&_net_2549);
   assign  _net_2894 = (_reg_2545&_net_2549);
   assign  _net_2895 = (_reg_2545&_net_2549);
   assign  _net_2896 = (_reg_2545&_net_2549);
   assign  _net_2897 = (_reg_2545&_net_2549);
   assign  _net_2898 = (_reg_2545&_net_2549);
   assign  _net_2899 = (_reg_2545&_net_2549);
   assign  _net_2900 = (_reg_2545&_net_2549);
   assign  _net_2901 = (_reg_2545&_net_2549);
   assign  _net_2902 = (_reg_2545&_net_2549);
   assign  _net_2903 = (_reg_2545&_net_2549);
   assign  _net_2904 = (_reg_2545&_net_2549);
   assign  _net_2905 = (_reg_2545&_net_2549);
   assign  _net_2906 = (_reg_2545&_net_2549);
   assign  _net_2907 = (_reg_2545&_net_2549);
   assign  _net_2908 = (_reg_2545&_net_2549);
   assign  _net_2909 = (_reg_2545&_net_2549);
   assign  _net_2910 = (_reg_2545&_net_2549);
   assign  _net_2911 = (_reg_2545&_net_2549);
   assign  _net_2912 = (_reg_2545&_net_2549);
   assign  _net_2913 = (_reg_2545&_net_2549);
   assign  _net_2914 = (_reg_2545&_net_2549);
   assign  _net_2915 = (_reg_2545&_net_2549);
   assign  _net_2916 = (_reg_2545&_net_2549);
   assign  _net_2917 = (_reg_2545&_net_2549);
   assign  _net_2918 = (_reg_2545&_net_2549);
   assign  _net_2919 = (_reg_2545&_net_2549);
   assign  _net_2920 = (_reg_2545&_net_2549);
   assign  _net_2921 = (_reg_2545&_net_2549);
   assign  _net_2922 = (_reg_2545&_net_2549);
   assign  _net_2923 = (_reg_2545&_net_2549);
   assign  _net_2924 = (_reg_2545&_net_2549);
   assign  _net_2925 = (_reg_2545&_net_2549);
   assign  _net_2926 = (_reg_2545&_net_2549);
   assign  _net_2927 = (_reg_2545&_net_2549);
   assign  _net_2928 = (_reg_2545&_net_2549);
   assign  _net_2929 = (_reg_2545&_net_2549);
   assign  _net_2930 = (_reg_2545&_net_2549);
   assign  _net_2931 = (_reg_2545&_net_2549);
   assign  _net_2932 = (_reg_2545&_net_2549);
   assign  _net_2933 = (_reg_2545&_net_2549);
   assign  _net_2934 = (_reg_2545&_net_2549);
   assign  _net_2935 = (_reg_2545&_net_2549);
   assign  _net_2936 = (_reg_2545&_net_2549);
   assign  _net_2937 = (_reg_2545&_net_2549);
   assign  _net_2938 = (_reg_2545&_net_2549);
   assign  _net_2939 = (_reg_2545&_net_2549);
   assign  _net_2940 = (_reg_2545&_net_2549);
   assign  _net_2941 = (_reg_2545&_net_2549);
   assign  _net_2942 = (_reg_2545&_net_2549);
   assign  _net_2943 = (_reg_2545&_net_2549);
   assign  _net_2944 = (_reg_2545&_net_2549);
   assign  _net_2945 = (_reg_2545&_net_2549);
   assign  _net_2946 = (_reg_2545&_net_2549);
   assign  _net_2947 = (_reg_2545&_net_2549);
   assign  _net_2948 = (_reg_2545&_net_2549);
   assign  _net_2949 = (_reg_2545&_net_2549);
   assign  _net_2950 = (_reg_2545&_net_2549);
   assign  _net_2951 = (_reg_2545&_net_2549);
   assign  _net_2952 = (_reg_2545&_net_2549);
   assign  _net_2953 = (_reg_2545&_net_2549);
   assign  _net_2954 = (_reg_2545&_net_2549);
   assign  _net_2955 = (_reg_2545&_net_2549);
   assign  _net_2956 = (_reg_2545&_net_2549);
   assign  _net_2957 = (_reg_2545&_net_2549);
   assign  _net_2958 = (_reg_2545&_net_2549);
   assign  _net_2959 = (_reg_2545&_net_2549);
   assign  _net_2960 = (_reg_2545&_net_2549);
   assign  _net_2961 = (_reg_2545&_net_2549);
   assign  _net_2962 = (_reg_2545&_net_2549);
   assign  _net_2963 = (_reg_2545&_net_2549);
   assign  _net_2964 = (_reg_2545&_net_2549);
   assign  _net_2965 = (_reg_2545&_net_2549);
   assign  _net_2966 = (_reg_2545&_net_2549);
   assign  _net_2967 = (_reg_2545&_net_2549);
   assign  _net_2968 = (_reg_2545&_net_2549);
   assign  _net_2969 = (_reg_2545&_net_2549);
   assign  _net_2970 = (_reg_2545&_net_2549);
   assign  _net_2971 = (_reg_2545&(~_net_2549));
   assign  _net_2972 = (_reg_2545&(~_net_2549));
   assign  _net_2973 = (_reg_2545&(~_net_2549));
   assign  _net_2974 = (_reg_2545&(~_net_2549));
   assign  _net_2975 = (_reg_2545&(~_net_2549));
   assign  _net_2976 = (_reg_2545&(~_net_2549));
   assign  _net_2977 = (_reg_2545&(~_net_2549));
   assign  _net_2978 = (_reg_2545&(~_net_2549));
   assign  _net_2979 = (_reg_2545&(~_net_2549));
   assign  _net_2980 = (_reg_2545&(~_net_2549));
   assign  _net_2981 = (_reg_2545&(~_net_2549));
   assign  _net_2982 = (_reg_2545&(~_net_2549));
   assign  _net_2983 = (_reg_2545&(~_net_2549));
   assign  _net_2984 = (_reg_2545&(~_net_2549));
   assign  _net_2985 = (_reg_2545&(~_net_2549));
   assign  _net_2986 = (_reg_2545&(~_net_2549));
   assign  _net_2987 = (_reg_2545&(~_net_2549));
   assign  _net_2988 = (_reg_2545&(~_net_2549));
   assign  _net_2989 = (_reg_2545&(~_net_2549));
   assign  _net_2990 = (_reg_2545&(~_net_2549));
   assign  _net_2991 = (_reg_2545&(~_net_2549));
   assign  _net_2992 = (_reg_2545&(~_net_2549));
   assign  _net_2993 = (_reg_2545&(~_net_2549));
   assign  _net_2994 = (_reg_2545&(~_net_2549));
   assign  _net_2995 = (_reg_2545&(~_net_2549));
   assign  _net_2996 = (_reg_2545&(~_net_2549));
   assign  _net_2997 = (_reg_2545&(~_net_2549));
   assign  _net_2998 = (_reg_2545&(~_net_2549));
   assign  _net_2999 = (_reg_2545&(~_net_2549));
   assign  _net_3000 = (_reg_2545&(~_net_2549));
   assign  _net_3001 = (_reg_2545&(~_net_2549));
   assign  _net_3002 = (_reg_2545&(~_net_2549));
   assign  _net_3003 = (_reg_2545&(~_net_2549));
   assign  _net_3004 = (_reg_2545&(~_net_2549));
   assign  _net_3005 = (_reg_2545&(~_net_2549));
   assign  _net_3006 = (_reg_2545&(~_net_2549));
   assign  _net_3007 = (_reg_2545&(~_net_2549));
   assign  _net_3008 = (_reg_2545&(~_net_2549));
   assign  _net_3009 = (_reg_2545&(~_net_2549));
   assign  _net_3010 = (_reg_2545&(~_net_2549));
   assign  _net_3011 = (_reg_2545&(~_net_2549));
   assign  _net_3012 = (_reg_2545&(~_net_2549));
   assign  _net_3013 = (_reg_2545&(~_net_2549));
   assign  _net_3014 = (_reg_2545&(~_net_2549));
   assign  _net_3015 = (_reg_2545&(~_net_2549));
   assign  _net_3016 = (_reg_2545&(~_net_2549));
   assign  _net_3017 = (_reg_2545&(~_net_2549));
   assign  _net_3018 = (_reg_2545&(~_net_2549));
   assign  _net_3019 = (_reg_2545&(~_net_2549));
   assign  _net_3020 = (_reg_2545&(~_net_2549));
   assign  _net_3021 = (_reg_2545&(~_net_2549));
   assign  _net_3022 = (_reg_2545&(~_net_2549));
   assign  _net_3023 = (_reg_2545&(~_net_2549));
   assign  _net_3024 = (_reg_2545&(~_net_2549));
   assign  _net_3025 = (_reg_2545&(~_net_2549));
   assign  _net_3026 = (_reg_2545&(~_net_2549));
   assign  _net_3027 = (_reg_2545&(~_net_2549));
   assign  _net_3028 = (_reg_2545&(~_net_2549));
   assign  _net_3029 = (_reg_2545&(~_net_2549));
   assign  _net_3030 = (_reg_2545&(~_net_2549));
   assign  _net_3031 = (_reg_2545&(~_net_2549));
   assign  _net_3032 = (_reg_2545&(~_net_2549));
   assign  _net_3033 = (_reg_2545&(~_net_2549));
   assign  _net_3034 = (_reg_2545&(~_net_2549));
   assign  _net_3035 = (_reg_2545&(~_net_2549));
   assign  _net_3036 = (_reg_2545&(~_net_2549));
   assign  _net_3037 = (_reg_2545&(~_net_2549));
   assign  _net_3038 = (_reg_2545&(~_net_2549));
   assign  _net_3039 = (_reg_2545&(~_net_2549));
   assign  _net_3040 = (_reg_2545&(~_net_2549));
   assign  _net_3041 = (_reg_2545&(~_net_2549));
   assign  _net_3042 = (_reg_2545&(~_net_2549));
   assign  _net_3043 = (_reg_2545&(~_net_2549));
   assign  _net_3044 = (_reg_2545&(~_net_2549));
   assign  _net_3045 = (_reg_2545&(~_net_2549));
   assign  _net_3046 = (_reg_2545&(~_net_2549));
   assign  _net_3047 = (_reg_2545&(~_net_2549));
   assign  _net_3048 = (_reg_2545&(~_net_2549));
   assign  _net_3049 = (_reg_2545&(~_net_2549));
   assign  _net_3050 = (_reg_2545&(~_net_2549));
   assign  _net_3051 = (_reg_2545&(~_net_2549));
   assign  _net_3052 = (_reg_2545&(~_net_2549));
   assign  _net_3053 = (_reg_2545&(~_net_2549));
   assign  _net_3054 = (_reg_2545&(~_net_2549));
   assign  _net_3055 = (_reg_2545&(~_net_2549));
   assign  _net_3056 = (_reg_2545&(~_net_2549));
   assign  _net_3057 = (_reg_2545&(~_net_2549));
   assign  _net_3058 = (_reg_2545&(~_net_2549));
   assign  _net_3059 = (_reg_2545&(~_net_2549));
   assign  _net_3060 = (_reg_2545&(~_net_2549));
   assign  _net_3061 = (_reg_2545&(~_net_2549));
   assign  _net_3062 = (_reg_2545&(~_net_2549));
   assign  _net_3063 = (_reg_2545&(~_net_2549));
   assign  _net_3064 = (_reg_2545&(~_net_2549));
   assign  _net_3065 = (_reg_2545&(~_net_2549));
   assign  _net_3066 = (_reg_2545&(~_net_2549));
   assign  _net_3067 = (_reg_2545&(~_net_2549));
   assign  _net_3068 = (_reg_2545&(~_net_2549));
   assign  _net_3069 = (_reg_2545&(~_net_2549));
   assign  _net_3070 = (_reg_2545&(~_net_2549));
   assign  _net_3071 = (_reg_2545&(~_net_2549));
   assign  _net_3072 = (_reg_2545&(~_net_2549));
   assign  _net_3073 = (_reg_2545&(~_net_2549));
   assign  _net_3074 = (_reg_2545&(~_net_2549));
   assign  _net_3075 = (_reg_2545&(~_net_2549));
   assign  _net_3076 = (_reg_2545&(~_net_2549));
   assign  _net_3077 = (_reg_2545&(~_net_2549));
   assign  _net_3078 = (_reg_2545&(~_net_2549));
   assign  _net_3079 = (_reg_2545&(~_net_2549));
   assign  _net_3080 = (_reg_2545&(~_net_2549));
   assign  _net_3081 = (_reg_2545&(~_net_2549));
   assign  _net_3082 = (_reg_2545&(~_net_2549));
   assign  _net_3083 = (_reg_2545&(~_net_2549));
   assign  _net_3084 = (_reg_2545&(~_net_2549));
   assign  _net_3085 = (_reg_2545&(~_net_2549));
   assign  _net_3086 = (_reg_2545&(~_net_2549));
   assign  _net_3087 = (_reg_2545&(~_net_2549));
   assign  _net_3088 = (_reg_2545&(~_net_2549));
   assign  _net_3089 = (_reg_2545&(~_net_2549));
   assign  _net_3090 = (_reg_2545&(~_net_2549));
   assign  _net_3091 = (_reg_2545&(~_net_2549));
   assign  _net_3092 = (_reg_2545&(~_net_2549));
   assign  _net_3093 = (_reg_2545&(~_net_2549));
   assign  _net_3094 = (_reg_2545&(~_net_2549));
   assign  _net_3095 = (_reg_2545&(~_net_2549));
   assign  _net_3096 = (_reg_2545&(~_net_2549));
   assign  _net_3097 = (_reg_2545&(~_net_2549));
   assign  _net_3098 = (_reg_2545&(~_net_2549));
   assign  _net_3099 = (_reg_2545&(~_net_2549));
   assign  _net_3100 = (_reg_2545&(~_net_2549));
   assign  _net_3101 = (_reg_2545&(~_net_2549));
   assign  _net_3102 = (_reg_2545&(~_net_2549));
   assign  _net_3103 = (_reg_2545&(~_net_2549));
   assign  _net_3104 = (_reg_2545&(~_net_2549));
   assign  _net_3105 = (_reg_2545&(~_net_2549));
   assign  _net_3106 = (_reg_2545&(~_net_2549));
   assign  _net_3107 = (_reg_2545&(~_net_2549));
   assign  _net_3108 = (_reg_2545&(~_net_2549));
   assign  _net_3109 = (_reg_2545&(~_net_2549));
   assign  _net_3110 = (_reg_2545&(~_net_2549));
   assign  _net_3111 = (_reg_2545&(~_net_2549));
   assign  _net_3112 = (_reg_2545&(~_net_2549));
   assign  _net_3113 = (_reg_2545&(~_net_2549));
   assign  _net_3114 = (_reg_2545&(~_net_2549));
   assign  _net_3115 = (_reg_2545&(~_net_2549));
   assign  _net_3116 = (_reg_2545&(~_net_2549));
   assign  _net_3117 = (_reg_2545&(~_net_2549));
   assign  _net_3118 = (_reg_2545&(~_net_2549));
   assign  _net_3119 = (_reg_2545&(~_net_2549));
   assign  _net_3120 = (_reg_2545&(~_net_2549));
   assign  _net_3121 = (_reg_2545&(~_net_2549));
   assign  _net_3122 = (_reg_2545&(~_net_2549));
   assign  _net_3123 = (_reg_2545&(~_net_2549));
   assign  _net_3124 = (_reg_2545&(~_net_2549));
   assign  _net_3125 = (_reg_2545&(~_net_2549));
   assign  _net_3126 = (_reg_2545&(~_net_2549));
   assign  _net_3127 = (_reg_2545&(~_net_2549));
   assign  _net_3128 = (_reg_2545&(~_net_2549));
   assign  _net_3129 = (_reg_2545&(~_net_2549));
   assign  _net_3130 = (_reg_2545&(~_net_2549));
   assign  _net_3131 = (_reg_2545&(~_net_2549));
   assign  _net_3132 = (_reg_2545&(~_net_2549));
   assign  _net_3133 = (_reg_2545&(~_net_2549));
   assign  _net_3134 = (_reg_2545&(~_net_2549));
   assign  _net_3135 = (_reg_2545&(~_net_2549));
   assign  _net_3136 = (_reg_2545&(~_net_2549));
   assign  _net_3137 = (_reg_2545&(~_net_2549));
   assign  _net_3138 = (_reg_2545&(~_net_2549));
   assign  _net_3139 = (_reg_2545&(~_net_2549));
   assign  _net_3140 = (_reg_2545&(~_net_2549));
   assign  _net_3141 = (_reg_2545&(~_net_2549));
   assign  _net_3142 = (_reg_2545&(~_net_2549));
   assign  _net_3143 = (_reg_2545&(~_net_2549));
   assign  _net_3144 = (_reg_2545&(~_net_2549));
   assign  _net_3145 = (_reg_2545&(~_net_2549));
   assign  _net_3146 = (_reg_2545&(~_net_2549));
   assign  _net_3147 = (_reg_2545&(~_net_2549));
   assign  _net_3148 = (_reg_2545&(~_net_2549));
   assign  _net_3149 = (_reg_2545&(~_net_2549));
   assign  _net_3150 = (_reg_2545&(~_net_2549));
   assign  _net_3151 = (_reg_2545&(~_net_2549));
   assign  _net_3152 = (_reg_2545&(~_net_2549));
   assign  _net_3153 = (_reg_2545&(~_net_2549));
   assign  _net_3154 = (_reg_2545&(~_net_2549));
   assign  _net_3155 = (_reg_2545&(~_net_2549));
   assign  _net_3156 = (_reg_2545&(~_net_2549));
   assign  _net_3157 = (_reg_2545&(~_net_2549));
   assign  _net_3158 = (_reg_2545&(~_net_2549));
   assign  _net_3159 = (_reg_2545&(~_net_2549));
   assign  _net_3160 = (_reg_2545&(~_net_2549));
   assign  _net_3161 = (_reg_2545&(~_net_2549));
   assign  _net_3162 = (_reg_2545&(~_net_2549));
   assign  _net_3163 = (_reg_2545&(~_net_2549));
   assign  _net_3164 = (_reg_2545&(~_net_2549));
   assign  _net_3165 = (_reg_2545&(~_net_2549));
   assign  _net_3166 = (_reg_2545&(~_net_2549));
   assign  _net_3167 = (_reg_2545&(~_net_2549));
   assign  _net_3168 = (_reg_2545&(~_net_2549));
   assign  _net_3169 = (_reg_2545&(~_net_2549));
   assign  _net_3170 = (_reg_2545&(~_net_2549));
   assign  _net_3171 = (_reg_2545&(~_net_2549));
   assign  _net_3172 = (_reg_2545&(~_net_2549));
   assign  _net_3173 = (_reg_2545&(~_net_2549));
   assign  _net_3174 = (_reg_2545&(~_net_2549));
   assign  _net_3175 = (_reg_2545&(~_net_2549));
   assign  _net_3176 = (_reg_2545&(~_net_2549));
   assign  _net_3177 = (_reg_2545&(~_net_2549));
   assign  _net_3178 = (_reg_2545&(~_net_2549));
   assign  _net_3179 = (_reg_2545&(~_net_2549));
   assign  _net_3180 = (_reg_2545&(~_net_2549));
   assign  _net_3181 = (_reg_2545&(~_net_2549));
   assign  _net_3182 = (_reg_2545&(~_net_2549));
   assign  _net_3183 = (_reg_2545&(~_net_2549));
   assign  _net_3184 = (_reg_2545&(~_net_2549));
   assign  _net_3185 = (_reg_2545&(~_net_2549));
   assign  _net_3186 = (_reg_2545&(~_net_2549));
   assign  _net_3187 = (_reg_2545&(~_net_2549));
   assign  _net_3188 = (_reg_2545&(~_net_2549));
   assign  _net_3189 = (_reg_2545&(~_net_2549));
   assign  _net_3190 = (_reg_2545&(~_net_2549));
   assign  _net_3191 = (_reg_2545&(~_net_2549));
   assign  _net_3192 = (_reg_2545&(~_net_2549));
   assign  _net_3193 = (_reg_2545&(~_net_2549));
   assign  _net_3194 = (_reg_2545&(~_net_2549));
   assign  _net_3195 = (_reg_2545&(~_net_2549));
   assign  _net_3196 = (_reg_2545&(~_net_2549));
   assign  _net_3197 = (_reg_2545&(~_net_2549));
   assign  _net_3198 = (_reg_2545&(~_net_2549));
   assign  _net_3199 = (_reg_2545&(~_net_2549));
   assign  _net_3200 = (_reg_2545&(~_net_2549));
   assign  _net_3201 = (_reg_2545&(~_net_2549));
   assign  _net_3202 = (_reg_2545&(~_net_2549));
   assign  _net_3203 = (_reg_2545&(~_net_2549));
   assign  _net_3204 = (_reg_2545&(~_net_2549));
   assign  _net_3205 = (_reg_2545&(~_net_2549));
   assign  _net_3206 = (_reg_2545&(~_net_2549));
   assign  _net_3207 = (_reg_2545&(~_net_2549));
   assign  _net_3208 = (_reg_2545&(~_net_2549));
   assign  _net_3209 = (_reg_2545&(~_net_2549));
   assign  _net_3210 = (_reg_2545&(~_net_2549));
   assign  _net_3211 = (_reg_2545&(~_net_2549));
   assign  _net_3212 = (_reg_2545&(~_net_2549));
   assign  _net_3213 = (_reg_2545&(~_net_2549));
   assign  _net_3214 = (_reg_2545&(~_net_2549));
   assign  _net_3215 = (_reg_2545&(~_net_2549));
   assign  _net_3216 = (_reg_2545&(~_net_2549));
   assign  _net_3217 = (_reg_2545&(~_net_2549));
   assign  _net_3218 = (_reg_2545&(~_net_2549));
   assign  _net_3219 = (_reg_2545&(~_net_2549));
   assign  _net_3220 = (_reg_2545&(~_net_2549));
   assign  _net_3221 = (_reg_2545&(~_net_2549));
   assign  _net_3222 = (_reg_2545&(~_net_2549));
   assign  _net_3223 = (_reg_2545&(~_net_2549));
   assign  _net_3224 = (_reg_2545&(~_net_2549));
   assign  _net_3225 = (_reg_2545&(~_net_2549));
   assign  _net_3226 = (_reg_2545&(~_net_2549));
   assign  _net_3227 = (_reg_2545&(~_net_2549));
   assign  _net_3228 = (_reg_2545&(~_net_2549));
   assign  _net_3229 = (_reg_2545&(~_net_2549));
   assign  _net_3230 = (_reg_2545&(~_net_2549));
   assign  _net_3231 = (_reg_2545&(~_net_2549));
   assign  _net_3232 = (_reg_2545&(~_net_2549));
   assign  _net_3233 = (_reg_2545&(~_net_2549));
   assign  _net_3234 = (_reg_2545&(~_net_2549));
   assign  _net_3235 = (_reg_2545&(~_net_2549));
   assign  _net_3236 = (_reg_2545&(~_net_2549));
   assign  _net_3237 = (_reg_2545&(~_net_2549));
   assign  _net_3238 = (_reg_2545&(~_net_2549));
   assign  _net_3239 = (_reg_2545&(~_net_2549));
   assign  _net_3240 = (_reg_2545&(~_net_2549));
   assign  _net_3241 = (_reg_2545&(~_net_2549));
   assign  _net_3242 = (_reg_2545&(~_net_2549));
   assign  _net_3243 = (_reg_2545&(~_net_2549));
   assign  _net_3244 = (_reg_2545&(~_net_2549));
   assign  _net_3245 = (_reg_2545&(~_net_2549));
   assign  _net_3246 = (_reg_2545&(~_net_2549));
   assign  _net_3247 = (_reg_2545&(~_net_2549));
   assign  _net_3248 = (_reg_2545&(~_net_2549));
   assign  _net_3249 = (_reg_2545&(~_net_2549));
   assign  _net_3250 = (_reg_2545&(~_net_2549));
   assign  _net_3251 = (_reg_2545&(~_net_2549));
   assign  _net_3252 = (_reg_2545&(~_net_2549));
   assign  _net_3253 = (_reg_2545&(~_net_2549));
   assign  _net_3254 = (_reg_2545&(~_net_2549));
   assign  _net_3255 = (_reg_2545&(~_net_2549));
   assign  _net_3256 = (_reg_2545&(~_net_2549));
   assign  _net_3257 = (_reg_2545&(~_net_2549));
   assign  _net_3258 = (_reg_2545&(~_net_2549));
   assign  _net_3259 = (_reg_2545&(~_net_2549));
   assign  _net_3260 = (_reg_2545&(~_net_2549));
   assign  _net_3261 = (_reg_2545&(~_net_2549));
   assign  _net_3262 = (_reg_2545&(~_net_2549));
   assign  _net_3263 = (_reg_2545&(~_net_2549));
   assign  _net_3264 = (_reg_2545&(~_net_2549));
   assign  _net_3265 = (_reg_2545&(~_net_2549));
   assign  _net_3266 = (_reg_2545&(~_net_2549));
   assign  _net_3267 = (_reg_2545&(~_net_2549));
   assign  _net_3268 = (_reg_2545&(~_net_2549));
   assign  _net_3269 = (_reg_2545&(~_net_2549));
   assign  _net_3270 = (_reg_2545&(~_net_2549));
   assign  _net_3271 = (_reg_2545&(~_net_2549));
   assign  _net_3272 = (_reg_2545&(~_net_2549));
   assign  _net_3273 = (_reg_2545&(~_net_2549));
   assign  _net_3274 = (_reg_2545&(~_net_2549));
   assign  _net_3275 = (_reg_2545&(~_net_2549));
   assign  _net_3276 = (_reg_2545&(~_net_2549));
   assign  _net_3277 = (_reg_2545&(~_net_2549));
   assign  _net_3278 = (_reg_2545&(~_net_2549));
   assign  _net_3279 = (_reg_2545&(~_net_2549));
   assign  _net_3280 = (_reg_2545&(~_net_2549));
   assign  _net_3281 = (_reg_2545&(~_net_2549));
   assign  _net_3282 = (_reg_2545&(~_net_2549));
   assign  _net_3283 = (_reg_2545&(~_net_2549));
   assign  _net_3284 = (_reg_2545&(~_net_2549));
   assign  _net_3285 = (_reg_2545&(~_net_2549));
   assign  _net_3286 = (_reg_2545&(~_net_2549));
   assign  _net_3287 = (_reg_2545&(~_net_2549));
   assign  _net_3288 = (_reg_2545&(~_net_2549));
   assign  _net_3289 = (_reg_2545&(~_net_2549));
   assign  _net_3290 = (_reg_2545&(~_net_2549));
   assign  _net_3291 = (_reg_2545&(~_net_2549));
   assign  _net_3292 = (_reg_2545&(~_net_2549));
   assign  _net_3293 = (_reg_2545&(~_net_2549));
   assign  _net_3294 = (_reg_2545&(~_net_2549));
   assign  _net_3295 = (_reg_2545&(~_net_2549));
   assign  _net_3296 = (_reg_2545&(~_net_2549));
   assign  _net_3297 = (_reg_2545&(~_net_2549));
   assign  _net_3298 = (_reg_2545&(~_net_2549));
   assign  _net_3299 = (_reg_2545&(~_net_2549));
   assign  _net_3300 = (_reg_2545&(~_net_2549));
   assign  _net_3301 = (_reg_2545&(~_net_2549));
   assign  _net_3302 = (_reg_2545&(~_net_2549));
   assign  _net_3303 = (_reg_2545&(~_net_2549));
   assign  _net_3304 = (_reg_2545&(~_net_2549));
   assign  _net_3305 = (_reg_2545&(~_net_2549));
   assign  _net_3306 = (_reg_2545&(~_net_2549));
   assign  _net_3307 = (_reg_2545&(~_net_2549));
   assign  _net_3308 = (_reg_2545&(~_net_2549));
   assign  _net_3309 = (_reg_2545&(~_net_2549));
   assign  _net_3310 = (_reg_2545&(~_net_2549));
   assign  _net_3311 = (_reg_2545&(~_net_2549));
   assign  _net_3312 = (_reg_2545&(~_net_2549));
   assign  _net_3313 = (_reg_2545&(~_net_2549));
   assign  _net_3314 = (_reg_2545&(~_net_2549));
   assign  _net_3315 = (_reg_2545&(~_net_2549));
   assign  _net_3316 = (_reg_2545&(~_net_2549));
   assign  _net_3317 = (_reg_2545&(~_net_2549));
   assign  _net_3318 = (_reg_2545&(~_net_2549));
   assign  _net_3319 = (_reg_2545&(~_net_2549));
   assign  _net_3320 = (_reg_2545&(~_net_2549));
   assign  _net_3321 = (_reg_2545&(~_net_2549));
   assign  _net_3322 = (_reg_2545&(~_net_2549));
   assign  _net_3323 = (_reg_2545&(~_net_2549));
   assign  _net_3324 = (_reg_2545&(~_net_2549));
   assign  _net_3325 = (_reg_2545&(~_net_2549));
   assign  _net_3326 = (_reg_2545&(~_net_2549));
   assign  _net_3327 = (_reg_2545&(~_net_2549));
   assign  _net_3328 = (_reg_2545&(~_net_2549));
   assign  _net_3329 = (_reg_2545&(~_net_2549));
   assign  _net_3330 = (_reg_2545&(~_net_2549));
   assign  _net_3331 = (_reg_2545&(~_net_2549));
   assign  _net_3332 = (_reg_2545&(~_net_2549));
   assign  _net_3333 = (_reg_2545&(~_net_2549));
   assign  _net_3334 = (_reg_2545&(~_net_2549));
   assign  _net_3335 = (_reg_2545&(~_net_2549));
   assign  _net_3336 = (_reg_2545&(~_net_2549));
   assign  _net_3337 = (_reg_2545&(~_net_2549));
   assign  _net_3338 = (_reg_2545&(~_net_2549));
   assign  _net_3339 = (_reg_2545&(~_net_2549));
   assign  _net_3340 = (_reg_2545&(~_net_2549));
   assign  _net_3341 = (_reg_2545&(~_net_2549));
   assign  _net_3342 = (_reg_2545&(~_net_2549));
   assign  _net_3343 = (_reg_2545&(~_net_2549));
   assign  _net_3344 = (_reg_2545&(~_net_2549));
   assign  _net_3345 = (_reg_2545&(~_net_2549));
   assign  _net_3346 = (_reg_2545&(~_net_2549));
   assign  _net_3347 = (_reg_2545&(~_net_2549));
   assign  _net_3348 = (_reg_2545&(~_net_2549));
   assign  _net_3349 = (_reg_2545&(~_net_2549));
   assign  _net_3350 = (_reg_2545&(~_net_2549));
   assign  _net_3351 = (_reg_2545&(~_net_2549));
   assign  _net_3352 = (_reg_2545&(~_net_2549));
   assign  _net_3353 = (_reg_2545&(~_net_2549));
   assign  _net_3354 = (_reg_2545&(~_net_2549));
   assign  _net_3355 = (_reg_2545&(~_net_2549));
   assign  _net_3356 = (_reg_2545&(~_net_2549));
   assign  _net_3357 = (_reg_2545&(~_net_2549));
   assign  _net_3358 = (_reg_2545&(~_net_2549));
   assign  _net_3359 = (_reg_2545&(~_net_2549));
   assign  _net_3360 = (_reg_2545&(~_net_2549));
   assign  _net_3361 = (_reg_2545&(~_net_2549));
   assign  _net_3362 = (_reg_2545&(~_net_2549));
   assign  _net_3363 = (_reg_2545&(~_net_2549));
   assign  _net_3364 = (_reg_2545&(~_net_2549));
   assign  _net_3365 = (_reg_2545&(~_net_2549));
   assign  _net_3366 = (_reg_2545&(~_net_2549));
   assign  _net_3367 = (_reg_2545&(~_net_2549));
   assign  _net_3368 = (_reg_2545&(~_net_2549));
   assign  _net_3369 = (_reg_2545&(~_net_2549));
   assign  _net_3370 = (_reg_2545&(~_net_2549));
   assign  _net_3371 = (_reg_2545&(~_net_2549));
   assign  _net_3372 = (_reg_2545&(~_net_2549));
   assign  _net_3373 = (_reg_2545&(~_net_2549));
   assign  _net_3374 = (_reg_2545&(~_net_2549));
   assign  _net_3375 = (_reg_2545&(~_net_2549));
   assign  _net_3376 = (_reg_2545&(~_net_2549));
   assign  _net_3377 = (_reg_2545&(~_net_2549));
   assign  _net_3378 = (_reg_2545&(~_net_2549));
   assign  _net_3379 = (_reg_2545&(~_net_2549));
   assign  _net_3380 = (_reg_2545&(~_net_2549));
   assign  _net_3381 = (_reg_2545&(~_net_2549));
   assign  _net_3382 = (_reg_2545&(~_net_2549));
   assign  _net_3383 = (_reg_2545&(~_net_2549));
   assign  _net_3384 = (_reg_2545&(~_net_2549));
   assign  _net_3385 = (_reg_2545&(~_net_2549));
   assign  _net_3386 = (_reg_2545&(~_net_2549));
   assign  _net_3387 = (_reg_2545&(~_net_2549));
   assign  _net_3388 = (_reg_2545&(~_net_2549));
   assign  _net_3389 = (_reg_2545&(~_net_2549));
   assign  _net_3390 = (_reg_2545&(~_net_2549));
   assign  _net_3391 = (_reg_2545&(~_net_2549));
   assign  _net_3392 = (dig_exit==1'b0);
   assign  _net_3393 = (_reg_2545&_net_3392);
   assign  _net_3394 = (_sub_x_sub_array_out < 10'b0000000001);
   assign  _net_3395 = (_reg_2545&(~_net_3392));
   assign  _net_3396 = ((_reg_2545&(~_net_3392))&_net_3394);

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_reg_2545)
    begin
    $display("sub %d",_sub_x_sub_array_out);
    end
  end

// synthesis translate_on
// synopsys translate_on
   assign  _net_3398 = (_add_all_x_out_do|(_reg_2545|_reg_2546));
   assign  data_out33 = _add_all_x_data_out_index33;
   assign  data_out34 = _add_all_x_data_out_index34;
   assign  data_out35 = _add_all_x_data_out_index35;
   assign  data_out36 = _add_all_x_data_out_index36;
   assign  data_out37 = _add_all_x_data_out_index37;
   assign  data_out38 = _add_all_x_data_out_index38;
   assign  data_out39 = _add_all_x_data_out_index39;
   assign  data_out40 = _add_all_x_data_out_index40;
   assign  data_out41 = _add_all_x_data_out_index41;
   assign  data_out42 = _add_all_x_data_out_index42;
   assign  data_out43 = _add_all_x_data_out_index43;
   assign  data_out44 = _add_all_x_data_out_index44;
   assign  data_out45 = _add_all_x_data_out_index45;
   assign  data_out46 = _add_all_x_data_out_index46;
   assign  data_out47 = _add_all_x_data_out_index47;
   assign  data_out48 = _add_all_x_data_out_index48;
   assign  data_out49 = _add_all_x_data_out_index49;
   assign  data_out50 = _add_all_x_data_out_index50;
   assign  data_out51 = _add_all_x_data_out_index51;
   assign  data_out52 = _add_all_x_data_out_index52;
   assign  data_out53 = _add_all_x_data_out_index53;
   assign  data_out54 = _add_all_x_data_out_index54;
   assign  data_out55 = _add_all_x_data_out_index55;
   assign  data_out56 = _add_all_x_data_out_index56;
   assign  data_out57 = _add_all_x_data_out_index57;
   assign  data_out58 = _add_all_x_data_out_index58;
   assign  data_out59 = _add_all_x_data_out_index59;
   assign  data_out60 = _add_all_x_data_out_index60;
   assign  data_out61 = _add_all_x_data_out_index61;
   assign  data_out62 = _add_all_x_data_out_index62;
   assign  data_out65 = _add_all_x_data_out_index65;
   assign  data_out66 = _add_all_x_data_out_index66;
   assign  data_out67 = _add_all_x_data_out_index67;
   assign  data_out68 = _add_all_x_data_out_index68;
   assign  data_out69 = _add_all_x_data_out_index69;
   assign  data_out70 = _add_all_x_data_out_index70;
   assign  data_out71 = _add_all_x_data_out_index71;
   assign  data_out72 = _add_all_x_data_out_index72;
   assign  data_out73 = _add_all_x_data_out_index73;
   assign  data_out74 = _add_all_x_data_out_index74;
   assign  data_out75 = _add_all_x_data_out_index75;
   assign  data_out76 = _add_all_x_data_out_index76;
   assign  data_out77 = _add_all_x_data_out_index77;
   assign  data_out78 = _add_all_x_data_out_index78;
   assign  data_out79 = _add_all_x_data_out_index79;
   assign  data_out80 = _add_all_x_data_out_index80;
   assign  data_out81 = _add_all_x_data_out_index81;
   assign  data_out82 = _add_all_x_data_out_index82;
   assign  data_out83 = _add_all_x_data_out_index83;
   assign  data_out84 = _add_all_x_data_out_index84;
   assign  data_out85 = _add_all_x_data_out_index85;
   assign  data_out86 = _add_all_x_data_out_index86;
   assign  data_out87 = _add_all_x_data_out_index87;
   assign  data_out88 = _add_all_x_data_out_index88;
   assign  data_out89 = _add_all_x_data_out_index89;
   assign  data_out90 = _add_all_x_data_out_index90;
   assign  data_out91 = _add_all_x_data_out_index91;
   assign  data_out92 = _add_all_x_data_out_index92;
   assign  data_out93 = _add_all_x_data_out_index93;
   assign  data_out94 = _add_all_x_data_out_index94;
   assign  data_out97 = _add_all_x_data_out_index97;
   assign  data_out98 = _add_all_x_data_out_index98;
   assign  data_out99 = _add_all_x_data_out_index99;
   assign  data_out100 = _add_all_x_data_out_index100;
   assign  data_out101 = _add_all_x_data_out_index101;
   assign  data_out102 = _add_all_x_data_out_index102;
   assign  data_out103 = _add_all_x_data_out_index103;
   assign  data_out104 = _add_all_x_data_out_index104;
   assign  data_out105 = _add_all_x_data_out_index105;
   assign  data_out106 = _add_all_x_data_out_index106;
   assign  data_out107 = _add_all_x_data_out_index107;
   assign  data_out108 = _add_all_x_data_out_index108;
   assign  data_out109 = _add_all_x_data_out_index109;
   assign  data_out110 = _add_all_x_data_out_index110;
   assign  data_out111 = _add_all_x_data_out_index111;
   assign  data_out112 = _add_all_x_data_out_index112;
   assign  data_out113 = _add_all_x_data_out_index113;
   assign  data_out114 = _add_all_x_data_out_index114;
   assign  data_out115 = _add_all_x_data_out_index115;
   assign  data_out116 = _add_all_x_data_out_index116;
   assign  data_out117 = _add_all_x_data_out_index117;
   assign  data_out118 = _add_all_x_data_out_index118;
   assign  data_out119 = _add_all_x_data_out_index119;
   assign  data_out120 = _add_all_x_data_out_index120;
   assign  data_out121 = _add_all_x_data_out_index121;
   assign  data_out122 = _add_all_x_data_out_index122;
   assign  data_out123 = _add_all_x_data_out_index123;
   assign  data_out124 = _add_all_x_data_out_index124;
   assign  data_out125 = _add_all_x_data_out_index125;
   assign  data_out126 = _add_all_x_data_out_index126;
   assign  data_out129 = _add_all_x_data_out_index129;
   assign  data_out130 = _add_all_x_data_out_index130;
   assign  data_out131 = _add_all_x_data_out_index131;
   assign  data_out132 = _add_all_x_data_out_index132;
   assign  data_out133 = _add_all_x_data_out_index133;
   assign  data_out134 = _add_all_x_data_out_index134;
   assign  data_out135 = _add_all_x_data_out_index135;
   assign  data_out136 = _add_all_x_data_out_index136;
   assign  data_out137 = _add_all_x_data_out_index137;
   assign  data_out138 = _add_all_x_data_out_index138;
   assign  data_out139 = _add_all_x_data_out_index139;
   assign  data_out140 = _add_all_x_data_out_index140;
   assign  data_out141 = _add_all_x_data_out_index141;
   assign  data_out142 = _add_all_x_data_out_index142;
   assign  data_out143 = _add_all_x_data_out_index143;
   assign  data_out144 = _add_all_x_data_out_index144;
   assign  data_out145 = _add_all_x_data_out_index145;
   assign  data_out146 = _add_all_x_data_out_index146;
   assign  data_out147 = _add_all_x_data_out_index147;
   assign  data_out148 = _add_all_x_data_out_index148;
   assign  data_out149 = _add_all_x_data_out_index149;
   assign  data_out150 = _add_all_x_data_out_index150;
   assign  data_out151 = _add_all_x_data_out_index151;
   assign  data_out152 = _add_all_x_data_out_index152;
   assign  data_out153 = _add_all_x_data_out_index153;
   assign  data_out154 = _add_all_x_data_out_index154;
   assign  data_out155 = _add_all_x_data_out_index155;
   assign  data_out156 = _add_all_x_data_out_index156;
   assign  data_out157 = _add_all_x_data_out_index157;
   assign  data_out158 = _add_all_x_data_out_index158;
   assign  data_out161 = _add_all_x_data_out_index161;
   assign  data_out162 = _add_all_x_data_out_index162;
   assign  data_out163 = _add_all_x_data_out_index163;
   assign  data_out164 = _add_all_x_data_out_index164;
   assign  data_out165 = _add_all_x_data_out_index165;
   assign  data_out166 = _add_all_x_data_out_index166;
   assign  data_out167 = _add_all_x_data_out_index167;
   assign  data_out168 = _add_all_x_data_out_index168;
   assign  data_out169 = _add_all_x_data_out_index169;
   assign  data_out170 = _add_all_x_data_out_index170;
   assign  data_out171 = _add_all_x_data_out_index171;
   assign  data_out172 = _add_all_x_data_out_index172;
   assign  data_out173 = _add_all_x_data_out_index173;
   assign  data_out174 = _add_all_x_data_out_index174;
   assign  data_out175 = _add_all_x_data_out_index175;
   assign  data_out176 = _add_all_x_data_out_index176;
   assign  data_out177 = _add_all_x_data_out_index177;
   assign  data_out178 = _add_all_x_data_out_index178;
   assign  data_out179 = _add_all_x_data_out_index179;
   assign  data_out180 = _add_all_x_data_out_index180;
   assign  data_out181 = _add_all_x_data_out_index181;
   assign  data_out182 = _add_all_x_data_out_index182;
   assign  data_out183 = _add_all_x_data_out_index183;
   assign  data_out184 = _add_all_x_data_out_index184;
   assign  data_out185 = _add_all_x_data_out_index185;
   assign  data_out186 = _add_all_x_data_out_index186;
   assign  data_out187 = _add_all_x_data_out_index187;
   assign  data_out188 = _add_all_x_data_out_index188;
   assign  data_out189 = _add_all_x_data_out_index189;
   assign  data_out190 = _add_all_x_data_out_index190;
   assign  data_out193 = _add_all_x_data_out_index193;
   assign  data_out194 = _add_all_x_data_out_index194;
   assign  data_out195 = _add_all_x_data_out_index195;
   assign  data_out196 = _add_all_x_data_out_index196;
   assign  data_out197 = _add_all_x_data_out_index197;
   assign  data_out198 = _add_all_x_data_out_index198;
   assign  data_out199 = _add_all_x_data_out_index199;
   assign  data_out200 = _add_all_x_data_out_index200;
   assign  data_out201 = _add_all_x_data_out_index201;
   assign  data_out202 = _add_all_x_data_out_index202;
   assign  data_out203 = _add_all_x_data_out_index203;
   assign  data_out204 = _add_all_x_data_out_index204;
   assign  data_out205 = _add_all_x_data_out_index205;
   assign  data_out206 = _add_all_x_data_out_index206;
   assign  data_out207 = _add_all_x_data_out_index207;
   assign  data_out208 = _add_all_x_data_out_index208;
   assign  data_out209 = _add_all_x_data_out_index209;
   assign  data_out210 = _add_all_x_data_out_index210;
   assign  data_out211 = _add_all_x_data_out_index211;
   assign  data_out212 = _add_all_x_data_out_index212;
   assign  data_out213 = _add_all_x_data_out_index213;
   assign  data_out214 = _add_all_x_data_out_index214;
   assign  data_out215 = _add_all_x_data_out_index215;
   assign  data_out216 = _add_all_x_data_out_index216;
   assign  data_out217 = _add_all_x_data_out_index217;
   assign  data_out218 = _add_all_x_data_out_index218;
   assign  data_out219 = _add_all_x_data_out_index219;
   assign  data_out220 = _add_all_x_data_out_index220;
   assign  data_out221 = _add_all_x_data_out_index221;
   assign  data_out222 = _add_all_x_data_out_index222;
   assign  data_out225 = _add_all_x_data_out_index225;
   assign  data_out226 = _add_all_x_data_out_index226;
   assign  data_out227 = _add_all_x_data_out_index227;
   assign  data_out228 = _add_all_x_data_out_index228;
   assign  data_out229 = _add_all_x_data_out_index229;
   assign  data_out230 = _add_all_x_data_out_index230;
   assign  data_out231 = _add_all_x_data_out_index231;
   assign  data_out232 = _add_all_x_data_out_index232;
   assign  data_out233 = _add_all_x_data_out_index233;
   assign  data_out234 = _add_all_x_data_out_index234;
   assign  data_out235 = _add_all_x_data_out_index235;
   assign  data_out236 = _add_all_x_data_out_index236;
   assign  data_out237 = _add_all_x_data_out_index237;
   assign  data_out238 = _add_all_x_data_out_index238;
   assign  data_out239 = _add_all_x_data_out_index239;
   assign  data_out240 = _add_all_x_data_out_index240;
   assign  data_out241 = _add_all_x_data_out_index241;
   assign  data_out242 = _add_all_x_data_out_index242;
   assign  data_out243 = _add_all_x_data_out_index243;
   assign  data_out244 = _add_all_x_data_out_index244;
   assign  data_out245 = _add_all_x_data_out_index245;
   assign  data_out246 = _add_all_x_data_out_index246;
   assign  data_out247 = _add_all_x_data_out_index247;
   assign  data_out248 = _add_all_x_data_out_index248;
   assign  data_out249 = _add_all_x_data_out_index249;
   assign  data_out250 = _add_all_x_data_out_index250;
   assign  data_out251 = _add_all_x_data_out_index251;
   assign  data_out252 = _add_all_x_data_out_index252;
   assign  data_out253 = _add_all_x_data_out_index253;
   assign  data_out254 = _add_all_x_data_out_index254;
   assign  data_out257 = _add_all_x_data_out_index257;
   assign  data_out258 = _add_all_x_data_out_index258;
   assign  data_out259 = _add_all_x_data_out_index259;
   assign  data_out260 = _add_all_x_data_out_index260;
   assign  data_out261 = _add_all_x_data_out_index261;
   assign  data_out262 = _add_all_x_data_out_index262;
   assign  data_out263 = _add_all_x_data_out_index263;
   assign  data_out264 = _add_all_x_data_out_index264;
   assign  data_out265 = _add_all_x_data_out_index265;
   assign  data_out266 = _add_all_x_data_out_index266;
   assign  data_out267 = _add_all_x_data_out_index267;
   assign  data_out268 = _add_all_x_data_out_index268;
   assign  data_out269 = _add_all_x_data_out_index269;
   assign  data_out270 = _add_all_x_data_out_index270;
   assign  data_out271 = _add_all_x_data_out_index271;
   assign  data_out272 = _add_all_x_data_out_index272;
   assign  data_out273 = _add_all_x_data_out_index273;
   assign  data_out274 = _add_all_x_data_out_index274;
   assign  data_out275 = _add_all_x_data_out_index275;
   assign  data_out276 = _add_all_x_data_out_index276;
   assign  data_out277 = _add_all_x_data_out_index277;
   assign  data_out278 = _add_all_x_data_out_index278;
   assign  data_out279 = _add_all_x_data_out_index279;
   assign  data_out280 = _add_all_x_data_out_index280;
   assign  data_out281 = _add_all_x_data_out_index281;
   assign  data_out282 = _add_all_x_data_out_index282;
   assign  data_out283 = _add_all_x_data_out_index283;
   assign  data_out284 = _add_all_x_data_out_index284;
   assign  data_out285 = _add_all_x_data_out_index285;
   assign  data_out286 = _add_all_x_data_out_index286;
   assign  data_out289 = _add_all_x_data_out_index289;
   assign  data_out290 = _add_all_x_data_out_index290;
   assign  data_out291 = _add_all_x_data_out_index291;
   assign  data_out292 = _add_all_x_data_out_index292;
   assign  data_out293 = _add_all_x_data_out_index293;
   assign  data_out294 = _add_all_x_data_out_index294;
   assign  data_out295 = _add_all_x_data_out_index295;
   assign  data_out296 = _add_all_x_data_out_index296;
   assign  data_out297 = _add_all_x_data_out_index297;
   assign  data_out298 = _add_all_x_data_out_index298;
   assign  data_out299 = _add_all_x_data_out_index299;
   assign  data_out300 = _add_all_x_data_out_index300;
   assign  data_out301 = _add_all_x_data_out_index301;
   assign  data_out302 = _add_all_x_data_out_index302;
   assign  data_out303 = _add_all_x_data_out_index303;
   assign  data_out304 = _add_all_x_data_out_index304;
   assign  data_out305 = _add_all_x_data_out_index305;
   assign  data_out306 = _add_all_x_data_out_index306;
   assign  data_out307 = _add_all_x_data_out_index307;
   assign  data_out308 = _add_all_x_data_out_index308;
   assign  data_out309 = _add_all_x_data_out_index309;
   assign  data_out310 = _add_all_x_data_out_index310;
   assign  data_out311 = _add_all_x_data_out_index311;
   assign  data_out312 = _add_all_x_data_out_index312;
   assign  data_out313 = _add_all_x_data_out_index313;
   assign  data_out314 = _add_all_x_data_out_index314;
   assign  data_out315 = _add_all_x_data_out_index315;
   assign  data_out316 = _add_all_x_data_out_index316;
   assign  data_out317 = _add_all_x_data_out_index317;
   assign  data_out318 = _add_all_x_data_out_index318;
   assign  data_out321 = _add_all_x_data_out_index321;
   assign  data_out322 = _add_all_x_data_out_index322;
   assign  data_out323 = _add_all_x_data_out_index323;
   assign  data_out324 = _add_all_x_data_out_index324;
   assign  data_out325 = _add_all_x_data_out_index325;
   assign  data_out326 = _add_all_x_data_out_index326;
   assign  data_out327 = _add_all_x_data_out_index327;
   assign  data_out328 = _add_all_x_data_out_index328;
   assign  data_out329 = _add_all_x_data_out_index329;
   assign  data_out330 = _add_all_x_data_out_index330;
   assign  data_out331 = _add_all_x_data_out_index331;
   assign  data_out332 = _add_all_x_data_out_index332;
   assign  data_out333 = _add_all_x_data_out_index333;
   assign  data_out334 = _add_all_x_data_out_index334;
   assign  data_out335 = _add_all_x_data_out_index335;
   assign  data_out336 = _add_all_x_data_out_index336;
   assign  data_out337 = _add_all_x_data_out_index337;
   assign  data_out338 = _add_all_x_data_out_index338;
   assign  data_out339 = _add_all_x_data_out_index339;
   assign  data_out340 = _add_all_x_data_out_index340;
   assign  data_out341 = _add_all_x_data_out_index341;
   assign  data_out342 = _add_all_x_data_out_index342;
   assign  data_out343 = _add_all_x_data_out_index343;
   assign  data_out344 = _add_all_x_data_out_index344;
   assign  data_out345 = _add_all_x_data_out_index345;
   assign  data_out346 = _add_all_x_data_out_index346;
   assign  data_out347 = _add_all_x_data_out_index347;
   assign  data_out348 = _add_all_x_data_out_index348;
   assign  data_out349 = _add_all_x_data_out_index349;
   assign  data_out350 = _add_all_x_data_out_index350;
   assign  data_out353 = _add_all_x_data_out_index353;
   assign  data_out354 = _add_all_x_data_out_index354;
   assign  data_out355 = _add_all_x_data_out_index355;
   assign  data_out356 = _add_all_x_data_out_index356;
   assign  data_out357 = _add_all_x_data_out_index357;
   assign  data_out358 = _add_all_x_data_out_index358;
   assign  data_out359 = _add_all_x_data_out_index359;
   assign  data_out360 = _add_all_x_data_out_index360;
   assign  data_out361 = _add_all_x_data_out_index361;
   assign  data_out362 = _add_all_x_data_out_index362;
   assign  data_out363 = _add_all_x_data_out_index363;
   assign  data_out364 = _add_all_x_data_out_index364;
   assign  data_out365 = _add_all_x_data_out_index365;
   assign  data_out366 = _add_all_x_data_out_index366;
   assign  data_out367 = _add_all_x_data_out_index367;
   assign  data_out368 = _add_all_x_data_out_index368;
   assign  data_out369 = _add_all_x_data_out_index369;
   assign  data_out370 = _add_all_x_data_out_index370;
   assign  data_out371 = _add_all_x_data_out_index371;
   assign  data_out372 = _add_all_x_data_out_index372;
   assign  data_out373 = _add_all_x_data_out_index373;
   assign  data_out374 = _add_all_x_data_out_index374;
   assign  data_out375 = _add_all_x_data_out_index375;
   assign  data_out376 = _add_all_x_data_out_index376;
   assign  data_out377 = _add_all_x_data_out_index377;
   assign  data_out378 = _add_all_x_data_out_index378;
   assign  data_out379 = _add_all_x_data_out_index379;
   assign  data_out380 = _add_all_x_data_out_index380;
   assign  data_out381 = _add_all_x_data_out_index381;
   assign  data_out382 = _add_all_x_data_out_index382;
   assign  data_out385 = _add_all_x_data_out_index385;
   assign  data_out386 = _add_all_x_data_out_index386;
   assign  data_out387 = _add_all_x_data_out_index387;
   assign  data_out388 = _add_all_x_data_out_index388;
   assign  data_out389 = _add_all_x_data_out_index389;
   assign  data_out390 = _add_all_x_data_out_index390;
   assign  data_out391 = _add_all_x_data_out_index391;
   assign  data_out392 = _add_all_x_data_out_index392;
   assign  data_out393 = _add_all_x_data_out_index393;
   assign  data_out394 = _add_all_x_data_out_index394;
   assign  data_out395 = _add_all_x_data_out_index395;
   assign  data_out396 = _add_all_x_data_out_index396;
   assign  data_out397 = _add_all_x_data_out_index397;
   assign  data_out398 = _add_all_x_data_out_index398;
   assign  data_out399 = _add_all_x_data_out_index399;
   assign  data_out400 = _add_all_x_data_out_index400;
   assign  data_out401 = _add_all_x_data_out_index401;
   assign  data_out402 = _add_all_x_data_out_index402;
   assign  data_out403 = _add_all_x_data_out_index403;
   assign  data_out404 = _add_all_x_data_out_index404;
   assign  data_out405 = _add_all_x_data_out_index405;
   assign  data_out406 = _add_all_x_data_out_index406;
   assign  data_out407 = _add_all_x_data_out_index407;
   assign  data_out408 = _add_all_x_data_out_index408;
   assign  data_out409 = _add_all_x_data_out_index409;
   assign  data_out410 = _add_all_x_data_out_index410;
   assign  data_out411 = _add_all_x_data_out_index411;
   assign  data_out412 = _add_all_x_data_out_index412;
   assign  data_out413 = _add_all_x_data_out_index413;
   assign  data_out414 = _add_all_x_data_out_index414;
   assign  data_out417 = _add_all_x_data_out_index417;
   assign  data_out418 = _add_all_x_data_out_index418;
   assign  data_out419 = _add_all_x_data_out_index419;
   assign  data_out420 = _add_all_x_data_out_index420;
   assign  data_out421 = _add_all_x_data_out_index421;
   assign  data_out422 = _add_all_x_data_out_index422;
   assign  data_out423 = _add_all_x_data_out_index423;
   assign  data_out424 = _add_all_x_data_out_index424;
   assign  data_out425 = _add_all_x_data_out_index425;
   assign  data_out426 = _add_all_x_data_out_index426;
   assign  data_out427 = _add_all_x_data_out_index427;
   assign  data_out428 = _add_all_x_data_out_index428;
   assign  data_out429 = _add_all_x_data_out_index429;
   assign  data_out430 = _add_all_x_data_out_index430;
   assign  data_out431 = _add_all_x_data_out_index431;
   assign  data_out432 = _add_all_x_data_out_index432;
   assign  data_out433 = _add_all_x_data_out_index433;
   assign  data_out434 = _add_all_x_data_out_index434;
   assign  data_out435 = _add_all_x_data_out_index435;
   assign  data_out436 = _add_all_x_data_out_index436;
   assign  data_out437 = _add_all_x_data_out_index437;
   assign  data_out438 = _add_all_x_data_out_index438;
   assign  data_out439 = _add_all_x_data_out_index439;
   assign  data_out440 = _add_all_x_data_out_index440;
   assign  data_out441 = _add_all_x_data_out_index441;
   assign  data_out442 = _add_all_x_data_out_index442;
   assign  data_out443 = _add_all_x_data_out_index443;
   assign  data_out444 = _add_all_x_data_out_index444;
   assign  data_out445 = _add_all_x_data_out_index445;
   assign  data_out446 = _add_all_x_data_out_index446;
   assign  data_out449 = _add_all_x_data_out_index449;
   assign  data_out450 = _add_all_x_data_out_index450;
   assign  data_out451 = _add_all_x_data_out_index451;
   assign  data_out452 = _add_all_x_data_out_index452;
   assign  data_out453 = _add_all_x_data_out_index453;
   assign  data_out454 = _add_all_x_data_out_index454;
   assign  data_out455 = _add_all_x_data_out_index455;
   assign  data_out456 = _add_all_x_data_out_index456;
   assign  data_out457 = _add_all_x_data_out_index457;
   assign  data_out458 = _add_all_x_data_out_index458;
   assign  data_out459 = _add_all_x_data_out_index459;
   assign  data_out460 = _add_all_x_data_out_index460;
   assign  data_out461 = _add_all_x_data_out_index461;
   assign  data_out462 = _add_all_x_data_out_index462;
   assign  data_out463 = _add_all_x_data_out_index463;
   assign  data_out464 = _add_all_x_data_out_index464;
   assign  data_out465 = _add_all_x_data_out_index465;
   assign  data_out466 = _add_all_x_data_out_index466;
   assign  data_out467 = _add_all_x_data_out_index467;
   assign  data_out468 = _add_all_x_data_out_index468;
   assign  data_out469 = _add_all_x_data_out_index469;
   assign  data_out470 = _add_all_x_data_out_index470;
   assign  data_out471 = _add_all_x_data_out_index471;
   assign  data_out472 = _add_all_x_data_out_index472;
   assign  data_out473 = _add_all_x_data_out_index473;
   assign  data_out474 = _add_all_x_data_out_index474;
   assign  data_out475 = _add_all_x_data_out_index475;
   assign  data_out476 = _add_all_x_data_out_index476;
   assign  data_out477 = _add_all_x_data_out_index477;
   assign  data_out478 = _add_all_x_data_out_index478;
   assign  out_do = _reg_0;
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     kanwa_exit <= 2'b00;
else if ((_net_3396)|(_net_3393)) 
      kanwa_exit <= ((_net_3396) ?(kanwa_exit+2'b01):2'b0)|
    ((_net_3393) ?2'b00:2'b0);

end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     start_reg <= 10'b0000000000;
else if ((_net_2540)) 
      start_reg <= start;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     goal_reg <= 10'b0000000000;
else if ((_net_2541)) 
      goal_reg <= goal;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     even <= 1'b0;
else if ((kanwa_s)) 
      even <= even_w1;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_0 <= 1'b0;
else if ((_net_2544)) 
      _reg_0 <= (_reg_1&(~_reg_1_goto));
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_1 <= 1'b0;
else if ((_net_2543)) 
      _reg_1 <= _reg_2;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_2 <= 1'b0;
else if ((_net_2542)) 
      _reg_2 <= (((_reg_1&_net_4)|_reg_3)|in_do);
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_3 <= 1'b0;
else if ((_reg_3)) 
      _reg_3 <= 1'b0;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_2545 <= 1'b0;
else if ((_net_3398)) 
      _reg_2545 <= (_reg_2546|_add_all_x_out_do);
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_2546 <= 1'b0;
else if ((_reg_2546)) 
      _reg_2546 <= 1'b0;
end
endmodule

/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 19:04:52 2023
 Licensed to :EVALUATION USER*/
