
/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 19:04:52 2023
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module test ( p_reset , m_clock , HEX0 );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  output HEX0;
  wire HEX0;
  reg [9:0] map_test [0:511];
  wire fpga_512_start;
  reg out_put_flag;
  reg [3:0] first;
  reg [3:0] second;
  reg [3:0] third;
  reg [31:0] count;
  reg [7:0] encode [0:15];
  wire out_put;
  reg [1:0] end_reg;
  wire [21:0] _mul_bit_x_mul_bit1;
  wire [21:0] _mul_bit_x_mul_bit2;
  wire [24:0] _mul_bit_x_mul_bit_result;
  wire _mul_bit_x_mul_bit_exe;
  wire _mul_bit_x_p_reset;
  wire _mul_bit_x_m_clock;
  wire [21:0] _mul_bit_x_1_mul_bit1;
  wire [21:0] _mul_bit_x_1_mul_bit2;
  wire [24:0] _mul_bit_x_1_mul_bit_result;
  wire _mul_bit_x_1_mul_bit_exe;
  wire _mul_bit_x_1_p_reset;
  wire _mul_bit_x_1_m_clock;
  wire [9:0] _meirotest_map_value_arg0;
  wire [9:0] _meirotest_map_value_arg1;
  wire [9:0] _meirotest_map_value_arg2;
  wire [9:0] _meirotest_map_value_arg3;
  wire [9:0] _meirotest_map_value_arg4;
  wire [9:0] _meirotest_map_value_arg5;
  wire [9:0] _meirotest_map_value_arg6;
  wire [9:0] _meirotest_map_value_arg7;
  wire [9:0] _meirotest_map_value_arg8;
  wire [9:0] _meirotest_map_value_arg9;
  wire [9:0] _meirotest_map_value_arg10;
  wire [9:0] _meirotest_map_value_arg11;
  wire [9:0] _meirotest_map_value_arg12;
  wire [9:0] _meirotest_map_value_arg13;
  wire [9:0] _meirotest_map_value_arg14;
  wire [9:0] _meirotest_map_value_arg15;
  wire [9:0] _meirotest_map_value_arg16;
  wire [9:0] _meirotest_map_value_arg17;
  wire [9:0] _meirotest_map_value_arg18;
  wire [9:0] _meirotest_map_value_arg19;
  wire [9:0] _meirotest_map_value_arg20;
  wire [9:0] _meirotest_map_value_arg21;
  wire [9:0] _meirotest_map_value_arg22;
  wire [9:0] _meirotest_map_value_arg23;
  wire [9:0] _meirotest_map_value_arg24;
  wire [9:0] _meirotest_map_value_arg25;
  wire [9:0] _meirotest_map_value_arg26;
  wire [9:0] _meirotest_map_value_arg27;
  wire [9:0] _meirotest_map_value_arg28;
  wire [9:0] _meirotest_map_value_arg29;
  wire [9:0] _meirotest_map_value_arg30;
  wire [9:0] _meirotest_map_value_arg31;
  wire [9:0] _meirotest_map_value_arg32;
  wire [9:0] _meirotest_map_value_arg33;
  wire [9:0] _meirotest_map_value_arg34;
  wire [9:0] _meirotest_map_value_arg35;
  wire [9:0] _meirotest_map_value_arg36;
  wire [9:0] _meirotest_map_value_arg37;
  wire [9:0] _meirotest_map_value_arg38;
  wire [9:0] _meirotest_map_value_arg39;
  wire [9:0] _meirotest_map_value_arg40;
  wire [9:0] _meirotest_map_value_arg41;
  wire [9:0] _meirotest_map_value_arg42;
  wire [9:0] _meirotest_map_value_arg43;
  wire [9:0] _meirotest_map_value_arg44;
  wire [9:0] _meirotest_map_value_arg45;
  wire [9:0] _meirotest_map_value_arg46;
  wire [9:0] _meirotest_map_value_arg47;
  wire [9:0] _meirotest_map_value_arg48;
  wire [9:0] _meirotest_map_value_arg49;
  wire [9:0] _meirotest_map_value_arg50;
  wire [9:0] _meirotest_map_value_arg51;
  wire [9:0] _meirotest_map_value_arg52;
  wire [9:0] _meirotest_map_value_arg53;
  wire [9:0] _meirotest_map_value_arg54;
  wire [9:0] _meirotest_map_value_arg55;
  wire [9:0] _meirotest_map_value_arg56;
  wire [9:0] _meirotest_map_value_arg57;
  wire [9:0] _meirotest_map_value_arg58;
  wire [9:0] _meirotest_map_value_arg59;
  wire [9:0] _meirotest_map_value_arg60;
  wire [9:0] _meirotest_map_value_arg61;
  wire [9:0] _meirotest_map_value_arg62;
  wire [9:0] _meirotest_map_value_arg63;
  wire [9:0] _meirotest_map_value_arg64;
  wire [9:0] _meirotest_map_value_arg65;
  wire [9:0] _meirotest_map_value_arg66;
  wire [9:0] _meirotest_map_value_arg67;
  wire [9:0] _meirotest_map_value_arg68;
  wire [9:0] _meirotest_map_value_arg69;
  wire [9:0] _meirotest_map_value_arg70;
  wire [9:0] _meirotest_map_value_arg71;
  wire [9:0] _meirotest_map_value_arg72;
  wire [9:0] _meirotest_map_value_arg73;
  wire [9:0] _meirotest_map_value_arg74;
  wire [9:0] _meirotest_map_value_arg75;
  wire [9:0] _meirotest_map_value_arg76;
  wire [9:0] _meirotest_map_value_arg77;
  wire [9:0] _meirotest_map_value_arg78;
  wire [9:0] _meirotest_map_value_arg79;
  wire [9:0] _meirotest_map_value_arg80;
  wire [9:0] _meirotest_map_value_arg81;
  wire [9:0] _meirotest_map_value_arg82;
  wire [9:0] _meirotest_map_value_arg83;
  wire [9:0] _meirotest_map_value_arg84;
  wire [9:0] _meirotest_map_value_arg85;
  wire [9:0] _meirotest_map_value_arg86;
  wire [9:0] _meirotest_map_value_arg87;
  wire [9:0] _meirotest_map_value_arg88;
  wire [9:0] _meirotest_map_value_arg89;
  wire [9:0] _meirotest_map_value_arg90;
  wire [9:0] _meirotest_map_value_arg91;
  wire [9:0] _meirotest_map_value_arg92;
  wire [9:0] _meirotest_map_value_arg93;
  wire [9:0] _meirotest_map_value_arg94;
  wire [9:0] _meirotest_map_value_arg95;
  wire [9:0] _meirotest_map_value_arg96;
  wire [9:0] _meirotest_map_value_arg97;
  wire [9:0] _meirotest_map_value_arg98;
  wire [9:0] _meirotest_map_value_arg99;
  wire [9:0] _meirotest_map_value_arg100;
  wire [9:0] _meirotest_map_value_arg101;
  wire [9:0] _meirotest_map_value_arg102;
  wire [9:0] _meirotest_map_value_arg103;
  wire [9:0] _meirotest_map_value_arg104;
  wire [9:0] _meirotest_map_value_arg105;
  wire [9:0] _meirotest_map_value_arg106;
  wire [9:0] _meirotest_map_value_arg107;
  wire [9:0] _meirotest_map_value_arg108;
  wire [9:0] _meirotest_map_value_arg109;
  wire [9:0] _meirotest_map_value_arg110;
  wire [9:0] _meirotest_map_value_arg111;
  wire [9:0] _meirotest_map_value_arg112;
  wire [9:0] _meirotest_map_value_arg113;
  wire [9:0] _meirotest_map_value_arg114;
  wire [9:0] _meirotest_map_value_arg115;
  wire [9:0] _meirotest_map_value_arg116;
  wire [9:0] _meirotest_map_value_arg117;
  wire [9:0] _meirotest_map_value_arg118;
  wire [9:0] _meirotest_map_value_arg119;
  wire [9:0] _meirotest_map_value_arg120;
  wire [9:0] _meirotest_map_value_arg121;
  wire [9:0] _meirotest_map_value_arg122;
  wire [9:0] _meirotest_map_value_arg123;
  wire [9:0] _meirotest_map_value_arg124;
  wire [9:0] _meirotest_map_value_arg125;
  wire [9:0] _meirotest_map_value_arg126;
  wire [9:0] _meirotest_map_value_arg127;
  wire [9:0] _meirotest_map_value_arg128;
  wire [9:0] _meirotest_map_value_arg129;
  wire [9:0] _meirotest_map_value_arg130;
  wire [9:0] _meirotest_map_value_arg131;
  wire [9:0] _meirotest_map_value_arg132;
  wire [9:0] _meirotest_map_value_arg133;
  wire [9:0] _meirotest_map_value_arg134;
  wire [9:0] _meirotest_map_value_arg135;
  wire [9:0] _meirotest_map_value_arg136;
  wire [9:0] _meirotest_map_value_arg137;
  wire [9:0] _meirotest_map_value_arg138;
  wire [9:0] _meirotest_map_value_arg139;
  wire [9:0] _meirotest_map_value_arg140;
  wire [9:0] _meirotest_map_value_arg141;
  wire [9:0] _meirotest_map_value_arg142;
  wire [9:0] _meirotest_map_value_arg143;
  wire [9:0] _meirotest_map_value_arg144;
  wire [9:0] _meirotest_map_value_arg145;
  wire [9:0] _meirotest_map_value_arg146;
  wire [9:0] _meirotest_map_value_arg147;
  wire [9:0] _meirotest_map_value_arg148;
  wire [9:0] _meirotest_map_value_arg149;
  wire [9:0] _meirotest_map_value_arg150;
  wire [9:0] _meirotest_map_value_arg151;
  wire [9:0] _meirotest_map_value_arg152;
  wire [9:0] _meirotest_map_value_arg153;
  wire [9:0] _meirotest_map_value_arg154;
  wire [9:0] _meirotest_map_value_arg155;
  wire [9:0] _meirotest_map_value_arg156;
  wire [9:0] _meirotest_map_value_arg157;
  wire [9:0] _meirotest_map_value_arg158;
  wire [9:0] _meirotest_map_value_arg159;
  wire [9:0] _meirotest_map_value_arg160;
  wire [9:0] _meirotest_map_value_arg161;
  wire [9:0] _meirotest_map_value_arg162;
  wire [9:0] _meirotest_map_value_arg163;
  wire [9:0] _meirotest_map_value_arg164;
  wire [9:0] _meirotest_map_value_arg165;
  wire [9:0] _meirotest_map_value_arg166;
  wire [9:0] _meirotest_map_value_arg167;
  wire [9:0] _meirotest_map_value_arg168;
  wire [9:0] _meirotest_map_value_arg169;
  wire [9:0] _meirotest_map_value_arg170;
  wire [9:0] _meirotest_map_value_arg171;
  wire [9:0] _meirotest_map_value_arg172;
  wire [9:0] _meirotest_map_value_arg173;
  wire [9:0] _meirotest_map_value_arg174;
  wire [9:0] _meirotest_map_value_arg175;
  wire [9:0] _meirotest_map_value_arg176;
  wire [9:0] _meirotest_map_value_arg177;
  wire [9:0] _meirotest_map_value_arg178;
  wire [9:0] _meirotest_map_value_arg179;
  wire [9:0] _meirotest_map_value_arg180;
  wire [9:0] _meirotest_map_value_arg181;
  wire [9:0] _meirotest_map_value_arg182;
  wire [9:0] _meirotest_map_value_arg183;
  wire [9:0] _meirotest_map_value_arg184;
  wire [9:0] _meirotest_map_value_arg185;
  wire [9:0] _meirotest_map_value_arg186;
  wire [9:0] _meirotest_map_value_arg187;
  wire [9:0] _meirotest_map_value_arg188;
  wire [9:0] _meirotest_map_value_arg189;
  wire [9:0] _meirotest_map_value_arg190;
  wire [9:0] _meirotest_map_value_arg191;
  wire [9:0] _meirotest_map_value_arg192;
  wire [9:0] _meirotest_map_value_arg193;
  wire [9:0] _meirotest_map_value_arg194;
  wire [9:0] _meirotest_map_value_arg195;
  wire [9:0] _meirotest_map_value_arg196;
  wire [9:0] _meirotest_map_value_arg197;
  wire [9:0] _meirotest_map_value_arg198;
  wire [9:0] _meirotest_map_value_arg199;
  wire [9:0] _meirotest_map_value_arg200;
  wire [9:0] _meirotest_map_value_arg201;
  wire [9:0] _meirotest_map_value_arg202;
  wire [9:0] _meirotest_map_value_arg203;
  wire [9:0] _meirotest_map_value_arg204;
  wire [9:0] _meirotest_map_value_arg205;
  wire [9:0] _meirotest_map_value_arg206;
  wire [9:0] _meirotest_map_value_arg207;
  wire [9:0] _meirotest_map_value_arg208;
  wire [9:0] _meirotest_map_value_arg209;
  wire [9:0] _meirotest_map_value_arg210;
  wire [9:0] _meirotest_map_value_arg211;
  wire [9:0] _meirotest_map_value_arg212;
  wire [9:0] _meirotest_map_value_arg213;
  wire [9:0] _meirotest_map_value_arg214;
  wire [9:0] _meirotest_map_value_arg215;
  wire [9:0] _meirotest_map_value_arg216;
  wire [9:0] _meirotest_map_value_arg217;
  wire [9:0] _meirotest_map_value_arg218;
  wire [9:0] _meirotest_map_value_arg219;
  wire [9:0] _meirotest_map_value_arg220;
  wire [9:0] _meirotest_map_value_arg221;
  wire [9:0] _meirotest_map_value_arg222;
  wire [9:0] _meirotest_map_value_arg223;
  wire [9:0] _meirotest_map_value_arg224;
  wire [9:0] _meirotest_map_value_arg225;
  wire [9:0] _meirotest_map_value_arg226;
  wire [9:0] _meirotest_map_value_arg227;
  wire [9:0] _meirotest_map_value_arg228;
  wire [9:0] _meirotest_map_value_arg229;
  wire [9:0] _meirotest_map_value_arg230;
  wire [9:0] _meirotest_map_value_arg231;
  wire [9:0] _meirotest_map_value_arg232;
  wire [9:0] _meirotest_map_value_arg233;
  wire [9:0] _meirotest_map_value_arg234;
  wire [9:0] _meirotest_map_value_arg235;
  wire [9:0] _meirotest_map_value_arg236;
  wire [9:0] _meirotest_map_value_arg237;
  wire [9:0] _meirotest_map_value_arg238;
  wire [9:0] _meirotest_map_value_arg239;
  wire [9:0] _meirotest_map_value_arg240;
  wire [9:0] _meirotest_map_value_arg241;
  wire [9:0] _meirotest_map_value_arg242;
  wire [9:0] _meirotest_map_value_arg243;
  wire [9:0] _meirotest_map_value_arg244;
  wire [9:0] _meirotest_map_value_arg245;
  wire [9:0] _meirotest_map_value_arg246;
  wire [9:0] _meirotest_map_value_arg247;
  wire [9:0] _meirotest_map_value_arg248;
  wire [9:0] _meirotest_map_value_arg249;
  wire [9:0] _meirotest_map_value_arg250;
  wire [9:0] _meirotest_map_value_arg251;
  wire [9:0] _meirotest_map_value_arg252;
  wire [9:0] _meirotest_map_value_arg253;
  wire [9:0] _meirotest_map_value_arg254;
  wire [9:0] _meirotest_map_value_arg255;
  wire [9:0] _meirotest_map_value_arg256;
  wire [9:0] _meirotest_map_value_arg257;
  wire [9:0] _meirotest_map_value_arg258;
  wire [9:0] _meirotest_map_value_arg259;
  wire [9:0] _meirotest_map_value_arg260;
  wire [9:0] _meirotest_map_value_arg261;
  wire [9:0] _meirotest_map_value_arg262;
  wire [9:0] _meirotest_map_value_arg263;
  wire [9:0] _meirotest_map_value_arg264;
  wire [9:0] _meirotest_map_value_arg265;
  wire [9:0] _meirotest_map_value_arg266;
  wire [9:0] _meirotest_map_value_arg267;
  wire [9:0] _meirotest_map_value_arg268;
  wire [9:0] _meirotest_map_value_arg269;
  wire [9:0] _meirotest_map_value_arg270;
  wire [9:0] _meirotest_map_value_arg271;
  wire [9:0] _meirotest_map_value_arg272;
  wire [9:0] _meirotest_map_value_arg273;
  wire [9:0] _meirotest_map_value_arg274;
  wire [9:0] _meirotest_map_value_arg275;
  wire [9:0] _meirotest_map_value_arg276;
  wire [9:0] _meirotest_map_value_arg277;
  wire [9:0] _meirotest_map_value_arg278;
  wire [9:0] _meirotest_map_value_arg279;
  wire [9:0] _meirotest_map_value_arg280;
  wire [9:0] _meirotest_map_value_arg281;
  wire [9:0] _meirotest_map_value_arg282;
  wire [9:0] _meirotest_map_value_arg283;
  wire [9:0] _meirotest_map_value_arg284;
  wire [9:0] _meirotest_map_value_arg285;
  wire [9:0] _meirotest_map_value_arg286;
  wire [9:0] _meirotest_map_value_arg287;
  wire [9:0] _meirotest_map_value_arg288;
  wire [9:0] _meirotest_map_value_arg289;
  wire [9:0] _meirotest_map_value_arg290;
  wire [9:0] _meirotest_map_value_arg291;
  wire [9:0] _meirotest_map_value_arg292;
  wire [9:0] _meirotest_map_value_arg293;
  wire [9:0] _meirotest_map_value_arg294;
  wire [9:0] _meirotest_map_value_arg295;
  wire [9:0] _meirotest_map_value_arg296;
  wire [9:0] _meirotest_map_value_arg297;
  wire [9:0] _meirotest_map_value_arg298;
  wire [9:0] _meirotest_map_value_arg299;
  wire [9:0] _meirotest_map_value_arg300;
  wire [9:0] _meirotest_map_value_arg301;
  wire [9:0] _meirotest_map_value_arg302;
  wire [9:0] _meirotest_map_value_arg303;
  wire [9:0] _meirotest_map_value_arg304;
  wire [9:0] _meirotest_map_value_arg305;
  wire [9:0] _meirotest_map_value_arg306;
  wire [9:0] _meirotest_map_value_arg307;
  wire [9:0] _meirotest_map_value_arg308;
  wire [9:0] _meirotest_map_value_arg309;
  wire [9:0] _meirotest_map_value_arg310;
  wire [9:0] _meirotest_map_value_arg311;
  wire [9:0] _meirotest_map_value_arg312;
  wire [9:0] _meirotest_map_value_arg313;
  wire [9:0] _meirotest_map_value_arg314;
  wire [9:0] _meirotest_map_value_arg315;
  wire [9:0] _meirotest_map_value_arg316;
  wire [9:0] _meirotest_map_value_arg317;
  wire [9:0] _meirotest_map_value_arg318;
  wire [9:0] _meirotest_map_value_arg319;
  wire [9:0] _meirotest_map_value_arg320;
  wire [9:0] _meirotest_map_value_arg321;
  wire [9:0] _meirotest_map_value_arg322;
  wire [9:0] _meirotest_map_value_arg323;
  wire [9:0] _meirotest_map_value_arg324;
  wire [9:0] _meirotest_map_value_arg325;
  wire [9:0] _meirotest_map_value_arg326;
  wire [9:0] _meirotest_map_value_arg327;
  wire [9:0] _meirotest_map_value_arg328;
  wire [9:0] _meirotest_map_value_arg329;
  wire [9:0] _meirotest_map_value_arg330;
  wire [9:0] _meirotest_map_value_arg331;
  wire [9:0] _meirotest_map_value_arg332;
  wire [9:0] _meirotest_map_value_arg333;
  wire [9:0] _meirotest_map_value_arg334;
  wire [9:0] _meirotest_map_value_arg335;
  wire [9:0] _meirotest_map_value_arg336;
  wire [9:0] _meirotest_map_value_arg337;
  wire [9:0] _meirotest_map_value_arg338;
  wire [9:0] _meirotest_map_value_arg339;
  wire [9:0] _meirotest_map_value_arg340;
  wire [9:0] _meirotest_map_value_arg341;
  wire [9:0] _meirotest_map_value_arg342;
  wire [9:0] _meirotest_map_value_arg343;
  wire [9:0] _meirotest_map_value_arg344;
  wire [9:0] _meirotest_map_value_arg345;
  wire [9:0] _meirotest_map_value_arg346;
  wire [9:0] _meirotest_map_value_arg347;
  wire [9:0] _meirotest_map_value_arg348;
  wire [9:0] _meirotest_map_value_arg349;
  wire [9:0] _meirotest_map_value_arg350;
  wire [9:0] _meirotest_map_value_arg351;
  wire [9:0] _meirotest_map_value_arg352;
  wire [9:0] _meirotest_map_value_arg353;
  wire [9:0] _meirotest_map_value_arg354;
  wire [9:0] _meirotest_map_value_arg355;
  wire [9:0] _meirotest_map_value_arg356;
  wire [9:0] _meirotest_map_value_arg357;
  wire [9:0] _meirotest_map_value_arg358;
  wire [9:0] _meirotest_map_value_arg359;
  wire [9:0] _meirotest_map_value_arg360;
  wire [9:0] _meirotest_map_value_arg361;
  wire [9:0] _meirotest_map_value_arg362;
  wire [9:0] _meirotest_map_value_arg363;
  wire [9:0] _meirotest_map_value_arg364;
  wire [9:0] _meirotest_map_value_arg365;
  wire [9:0] _meirotest_map_value_arg366;
  wire [9:0] _meirotest_map_value_arg367;
  wire [9:0] _meirotest_map_value_arg368;
  wire [9:0] _meirotest_map_value_arg369;
  wire [9:0] _meirotest_map_value_arg370;
  wire [9:0] _meirotest_map_value_arg371;
  wire [9:0] _meirotest_map_value_arg372;
  wire [9:0] _meirotest_map_value_arg373;
  wire [9:0] _meirotest_map_value_arg374;
  wire [9:0] _meirotest_map_value_arg375;
  wire [9:0] _meirotest_map_value_arg376;
  wire [9:0] _meirotest_map_value_arg377;
  wire [9:0] _meirotest_map_value_arg378;
  wire [9:0] _meirotest_map_value_arg379;
  wire [9:0] _meirotest_map_value_arg380;
  wire [9:0] _meirotest_map_value_arg381;
  wire [9:0] _meirotest_map_value_arg382;
  wire [9:0] _meirotest_map_value_arg383;
  wire [9:0] _meirotest_map_value_arg384;
  wire [9:0] _meirotest_map_value_arg385;
  wire [9:0] _meirotest_map_value_arg386;
  wire [9:0] _meirotest_map_value_arg387;
  wire [9:0] _meirotest_map_value_arg388;
  wire [9:0] _meirotest_map_value_arg389;
  wire [9:0] _meirotest_map_value_arg390;
  wire [9:0] _meirotest_map_value_arg391;
  wire [9:0] _meirotest_map_value_arg392;
  wire [9:0] _meirotest_map_value_arg393;
  wire [9:0] _meirotest_map_value_arg394;
  wire [9:0] _meirotest_map_value_arg395;
  wire [9:0] _meirotest_map_value_arg396;
  wire [9:0] _meirotest_map_value_arg397;
  wire [9:0] _meirotest_map_value_arg398;
  wire [9:0] _meirotest_map_value_arg399;
  wire [9:0] _meirotest_map_value_arg400;
  wire [9:0] _meirotest_map_value_arg401;
  wire [9:0] _meirotest_map_value_arg402;
  wire [9:0] _meirotest_map_value_arg403;
  wire [9:0] _meirotest_map_value_arg404;
  wire [9:0] _meirotest_map_value_arg405;
  wire [9:0] _meirotest_map_value_arg406;
  wire [9:0] _meirotest_map_value_arg407;
  wire [9:0] _meirotest_map_value_arg408;
  wire [9:0] _meirotest_map_value_arg409;
  wire [9:0] _meirotest_map_value_arg410;
  wire [9:0] _meirotest_map_value_arg411;
  wire [9:0] _meirotest_map_value_arg412;
  wire [9:0] _meirotest_map_value_arg413;
  wire [9:0] _meirotest_map_value_arg414;
  wire [9:0] _meirotest_map_value_arg415;
  wire [9:0] _meirotest_map_value_arg416;
  wire [9:0] _meirotest_map_value_arg417;
  wire [9:0] _meirotest_map_value_arg418;
  wire [9:0] _meirotest_map_value_arg419;
  wire [9:0] _meirotest_map_value_arg420;
  wire [9:0] _meirotest_map_value_arg421;
  wire [9:0] _meirotest_map_value_arg422;
  wire [9:0] _meirotest_map_value_arg423;
  wire [9:0] _meirotest_map_value_arg424;
  wire [9:0] _meirotest_map_value_arg425;
  wire [9:0] _meirotest_map_value_arg426;
  wire [9:0] _meirotest_map_value_arg427;
  wire [9:0] _meirotest_map_value_arg428;
  wire [9:0] _meirotest_map_value_arg429;
  wire [9:0] _meirotest_map_value_arg430;
  wire [9:0] _meirotest_map_value_arg431;
  wire [9:0] _meirotest_map_value_arg432;
  wire [9:0] _meirotest_map_value_arg433;
  wire [9:0] _meirotest_map_value_arg434;
  wire [9:0] _meirotest_map_value_arg435;
  wire [9:0] _meirotest_map_value_arg436;
  wire [9:0] _meirotest_map_value_arg437;
  wire [9:0] _meirotest_map_value_arg438;
  wire [9:0] _meirotest_map_value_arg439;
  wire [9:0] _meirotest_map_value_arg440;
  wire [9:0] _meirotest_map_value_arg441;
  wire [9:0] _meirotest_map_value_arg442;
  wire [9:0] _meirotest_map_value_arg443;
  wire [9:0] _meirotest_map_value_arg444;
  wire [9:0] _meirotest_map_value_arg445;
  wire [9:0] _meirotest_map_value_arg446;
  wire [9:0] _meirotest_map_value_arg447;
  wire [9:0] _meirotest_map_value_arg448;
  wire [9:0] _meirotest_map_value_arg449;
  wire [9:0] _meirotest_map_value_arg450;
  wire [9:0] _meirotest_map_value_arg451;
  wire [9:0] _meirotest_map_value_arg452;
  wire [9:0] _meirotest_map_value_arg453;
  wire [9:0] _meirotest_map_value_arg454;
  wire [9:0] _meirotest_map_value_arg455;
  wire [9:0] _meirotest_map_value_arg456;
  wire [9:0] _meirotest_map_value_arg457;
  wire [9:0] _meirotest_map_value_arg458;
  wire [9:0] _meirotest_map_value_arg459;
  wire [9:0] _meirotest_map_value_arg460;
  wire [9:0] _meirotest_map_value_arg461;
  wire [9:0] _meirotest_map_value_arg462;
  wire [9:0] _meirotest_map_value_arg463;
  wire [9:0] _meirotest_map_value_arg464;
  wire [9:0] _meirotest_map_value_arg465;
  wire [9:0] _meirotest_map_value_arg466;
  wire [9:0] _meirotest_map_value_arg467;
  wire [9:0] _meirotest_map_value_arg468;
  wire [9:0] _meirotest_map_value_arg469;
  wire [9:0] _meirotest_map_value_arg470;
  wire [9:0] _meirotest_map_value_arg471;
  wire [9:0] _meirotest_map_value_arg472;
  wire [9:0] _meirotest_map_value_arg473;
  wire [9:0] _meirotest_map_value_arg474;
  wire [9:0] _meirotest_map_value_arg475;
  wire [9:0] _meirotest_map_value_arg476;
  wire [9:0] _meirotest_map_value_arg477;
  wire [9:0] _meirotest_map_value_arg478;
  wire [9:0] _meirotest_map_value_arg479;
  wire [9:0] _meirotest_map_value_arg480;
  wire [9:0] _meirotest_map_value_arg481;
  wire [9:0] _meirotest_map_value_arg482;
  wire [9:0] _meirotest_map_value_arg483;
  wire [9:0] _meirotest_map_value_arg484;
  wire [9:0] _meirotest_map_value_arg485;
  wire [9:0] _meirotest_map_value_arg486;
  wire [9:0] _meirotest_map_value_arg487;
  wire [9:0] _meirotest_map_value_arg488;
  wire [9:0] _meirotest_map_value_arg489;
  wire [9:0] _meirotest_map_value_arg490;
  wire [9:0] _meirotest_map_value_arg491;
  wire [9:0] _meirotest_map_value_arg492;
  wire [9:0] _meirotest_map_value_arg493;
  wire [9:0] _meirotest_map_value_arg494;
  wire [9:0] _meirotest_map_value_arg495;
  wire [9:0] _meirotest_map_value_arg496;
  wire [9:0] _meirotest_map_value_arg497;
  wire [9:0] _meirotest_map_value_arg498;
  wire [9:0] _meirotest_map_value_arg499;
  wire [9:0] _meirotest_map_value_arg500;
  wire [9:0] _meirotest_map_value_arg501;
  wire [9:0] _meirotest_map_value_arg502;
  wire [9:0] _meirotest_map_value_arg503;
  wire [9:0] _meirotest_map_value_arg504;
  wire [9:0] _meirotest_map_value_arg505;
  wire [9:0] _meirotest_map_value_arg506;
  wire [9:0] _meirotest_map_value_arg507;
  wire [9:0] _meirotest_map_value_arg508;
  wire [9:0] _meirotest_map_value_arg509;
  wire [9:0] _meirotest_map_value_arg510;
  wire [9:0] _meirotest_map_value_arg511;
  wire [9:0] _meirotest_kekka_out0;
  wire [9:0] _meirotest_kekka_out1;
  wire [9:0] _meirotest_kekka_out2;
  wire [9:0] _meirotest_kekka_out3;
  wire [9:0] _meirotest_kekka_out4;
  wire [9:0] _meirotest_kekka_out5;
  wire [9:0] _meirotest_kekka_out6;
  wire [9:0] _meirotest_kekka_out7;
  wire [9:0] _meirotest_kekka_out8;
  wire [9:0] _meirotest_kekka_out9;
  wire [9:0] _meirotest_kekka_out10;
  wire [9:0] _meirotest_kekka_out11;
  wire [9:0] _meirotest_kekka_out12;
  wire [9:0] _meirotest_kekka_out13;
  wire [9:0] _meirotest_kekka_out14;
  wire [9:0] _meirotest_kekka_out15;
  wire [9:0] _meirotest_kekka_out16;
  wire [9:0] _meirotest_kekka_out17;
  wire [9:0] _meirotest_kekka_out18;
  wire [9:0] _meirotest_kekka_out19;
  wire [9:0] _meirotest_kekka_out20;
  wire [9:0] _meirotest_kekka_out21;
  wire [9:0] _meirotest_kekka_out22;
  wire [9:0] _meirotest_kekka_out23;
  wire [9:0] _meirotest_kekka_out24;
  wire [9:0] _meirotest_kekka_out25;
  wire [9:0] _meirotest_kekka_out26;
  wire [9:0] _meirotest_kekka_out27;
  wire [9:0] _meirotest_kekka_out28;
  wire [9:0] _meirotest_kekka_out29;
  wire [9:0] _meirotest_kekka_out30;
  wire [9:0] _meirotest_kekka_out31;
  wire [9:0] _meirotest_kekka_out32;
  wire [9:0] _meirotest_kekka_out33;
  wire [9:0] _meirotest_kekka_out34;
  wire [9:0] _meirotest_kekka_out35;
  wire [9:0] _meirotest_kekka_out36;
  wire [9:0] _meirotest_kekka_out37;
  wire [9:0] _meirotest_kekka_out38;
  wire [9:0] _meirotest_kekka_out39;
  wire [9:0] _meirotest_kekka_out40;
  wire [9:0] _meirotest_kekka_out41;
  wire [9:0] _meirotest_kekka_out42;
  wire [9:0] _meirotest_kekka_out43;
  wire [9:0] _meirotest_kekka_out44;
  wire [9:0] _meirotest_kekka_out45;
  wire [9:0] _meirotest_kekka_out46;
  wire [9:0] _meirotest_kekka_out47;
  wire [9:0] _meirotest_kekka_out48;
  wire [9:0] _meirotest_kekka_out49;
  wire [9:0] _meirotest_kekka_out50;
  wire [9:0] _meirotest_kekka_out51;
  wire [9:0] _meirotest_kekka_out52;
  wire [9:0] _meirotest_kekka_out53;
  wire [9:0] _meirotest_kekka_out54;
  wire [9:0] _meirotest_kekka_out55;
  wire [9:0] _meirotest_kekka_out56;
  wire [9:0] _meirotest_kekka_out57;
  wire [9:0] _meirotest_kekka_out58;
  wire [9:0] _meirotest_kekka_out59;
  wire [9:0] _meirotest_kekka_out60;
  wire [9:0] _meirotest_kekka_out61;
  wire [9:0] _meirotest_kekka_out62;
  wire [9:0] _meirotest_kekka_out63;
  wire [9:0] _meirotest_kekka_out64;
  wire [9:0] _meirotest_kekka_out65;
  wire [9:0] _meirotest_kekka_out66;
  wire [9:0] _meirotest_kekka_out67;
  wire [9:0] _meirotest_kekka_out68;
  wire [9:0] _meirotest_kekka_out69;
  wire [9:0] _meirotest_kekka_out70;
  wire [9:0] _meirotest_kekka_out71;
  wire [9:0] _meirotest_kekka_out72;
  wire [9:0] _meirotest_kekka_out73;
  wire [9:0] _meirotest_kekka_out74;
  wire [9:0] _meirotest_kekka_out75;
  wire [9:0] _meirotest_kekka_out76;
  wire [9:0] _meirotest_kekka_out77;
  wire [9:0] _meirotest_kekka_out78;
  wire [9:0] _meirotest_kekka_out79;
  wire [9:0] _meirotest_kekka_out80;
  wire [9:0] _meirotest_kekka_out81;
  wire [9:0] _meirotest_kekka_out82;
  wire [9:0] _meirotest_kekka_out83;
  wire [9:0] _meirotest_kekka_out84;
  wire [9:0] _meirotest_kekka_out85;
  wire [9:0] _meirotest_kekka_out86;
  wire [9:0] _meirotest_kekka_out87;
  wire [9:0] _meirotest_kekka_out88;
  wire [9:0] _meirotest_kekka_out89;
  wire [9:0] _meirotest_kekka_out90;
  wire [9:0] _meirotest_kekka_out91;
  wire [9:0] _meirotest_kekka_out92;
  wire [9:0] _meirotest_kekka_out93;
  wire [9:0] _meirotest_kekka_out94;
  wire [9:0] _meirotest_kekka_out95;
  wire [9:0] _meirotest_kekka_out96;
  wire [9:0] _meirotest_kekka_out97;
  wire [9:0] _meirotest_kekka_out98;
  wire [9:0] _meirotest_kekka_out99;
  wire [9:0] _meirotest_kekka_out100;
  wire [9:0] _meirotest_kekka_out101;
  wire [9:0] _meirotest_kekka_out102;
  wire [9:0] _meirotest_kekka_out103;
  wire [9:0] _meirotest_kekka_out104;
  wire [9:0] _meirotest_kekka_out105;
  wire [9:0] _meirotest_kekka_out106;
  wire [9:0] _meirotest_kekka_out107;
  wire [9:0] _meirotest_kekka_out108;
  wire [9:0] _meirotest_kekka_out109;
  wire [9:0] _meirotest_kekka_out110;
  wire [9:0] _meirotest_kekka_out111;
  wire [9:0] _meirotest_kekka_out112;
  wire [9:0] _meirotest_kekka_out113;
  wire [9:0] _meirotest_kekka_out114;
  wire [9:0] _meirotest_kekka_out115;
  wire [9:0] _meirotest_kekka_out116;
  wire [9:0] _meirotest_kekka_out117;
  wire [9:0] _meirotest_kekka_out118;
  wire [9:0] _meirotest_kekka_out119;
  wire [9:0] _meirotest_kekka_out120;
  wire [9:0] _meirotest_kekka_out121;
  wire [9:0] _meirotest_kekka_out122;
  wire [9:0] _meirotest_kekka_out123;
  wire [9:0] _meirotest_kekka_out124;
  wire [9:0] _meirotest_kekka_out125;
  wire [9:0] _meirotest_kekka_out126;
  wire [9:0] _meirotest_kekka_out127;
  wire [9:0] _meirotest_kekka_out128;
  wire [9:0] _meirotest_kekka_out129;
  wire [9:0] _meirotest_kekka_out130;
  wire [9:0] _meirotest_kekka_out131;
  wire [9:0] _meirotest_kekka_out132;
  wire [9:0] _meirotest_kekka_out133;
  wire [9:0] _meirotest_kekka_out134;
  wire [9:0] _meirotest_kekka_out135;
  wire [9:0] _meirotest_kekka_out136;
  wire [9:0] _meirotest_kekka_out137;
  wire [9:0] _meirotest_kekka_out138;
  wire [9:0] _meirotest_kekka_out139;
  wire [9:0] _meirotest_kekka_out140;
  wire [9:0] _meirotest_kekka_out141;
  wire [9:0] _meirotest_kekka_out142;
  wire [9:0] _meirotest_kekka_out143;
  wire [9:0] _meirotest_kekka_out144;
  wire [9:0] _meirotest_kekka_out145;
  wire [9:0] _meirotest_kekka_out146;
  wire [9:0] _meirotest_kekka_out147;
  wire [9:0] _meirotest_kekka_out148;
  wire [9:0] _meirotest_kekka_out149;
  wire [9:0] _meirotest_kekka_out150;
  wire [9:0] _meirotest_kekka_out151;
  wire [9:0] _meirotest_kekka_out152;
  wire [9:0] _meirotest_kekka_out153;
  wire [9:0] _meirotest_kekka_out154;
  wire [9:0] _meirotest_kekka_out155;
  wire [9:0] _meirotest_kekka_out156;
  wire [9:0] _meirotest_kekka_out157;
  wire [9:0] _meirotest_kekka_out158;
  wire [9:0] _meirotest_kekka_out159;
  wire [9:0] _meirotest_kekka_out160;
  wire [9:0] _meirotest_kekka_out161;
  wire [9:0] _meirotest_kekka_out162;
  wire [9:0] _meirotest_kekka_out163;
  wire [9:0] _meirotest_kekka_out164;
  wire [9:0] _meirotest_kekka_out165;
  wire [9:0] _meirotest_kekka_out166;
  wire [9:0] _meirotest_kekka_out167;
  wire [9:0] _meirotest_kekka_out168;
  wire [9:0] _meirotest_kekka_out169;
  wire [9:0] _meirotest_kekka_out170;
  wire [9:0] _meirotest_kekka_out171;
  wire [9:0] _meirotest_kekka_out172;
  wire [9:0] _meirotest_kekka_out173;
  wire [9:0] _meirotest_kekka_out174;
  wire [9:0] _meirotest_kekka_out175;
  wire [9:0] _meirotest_kekka_out176;
  wire [9:0] _meirotest_kekka_out177;
  wire [9:0] _meirotest_kekka_out178;
  wire [9:0] _meirotest_kekka_out179;
  wire [9:0] _meirotest_kekka_out180;
  wire [9:0] _meirotest_kekka_out181;
  wire [9:0] _meirotest_kekka_out182;
  wire [9:0] _meirotest_kekka_out183;
  wire [9:0] _meirotest_kekka_out184;
  wire [9:0] _meirotest_kekka_out185;
  wire [9:0] _meirotest_kekka_out186;
  wire [9:0] _meirotest_kekka_out187;
  wire [9:0] _meirotest_kekka_out188;
  wire [9:0] _meirotest_kekka_out189;
  wire [9:0] _meirotest_kekka_out190;
  wire [9:0] _meirotest_kekka_out191;
  wire [9:0] _meirotest_kekka_out192;
  wire [9:0] _meirotest_kekka_out193;
  wire [9:0] _meirotest_kekka_out194;
  wire [9:0] _meirotest_kekka_out195;
  wire [9:0] _meirotest_kekka_out196;
  wire [9:0] _meirotest_kekka_out197;
  wire [9:0] _meirotest_kekka_out198;
  wire [9:0] _meirotest_kekka_out199;
  wire [9:0] _meirotest_kekka_out200;
  wire [9:0] _meirotest_kekka_out201;
  wire [9:0] _meirotest_kekka_out202;
  wire [9:0] _meirotest_kekka_out203;
  wire [9:0] _meirotest_kekka_out204;
  wire [9:0] _meirotest_kekka_out205;
  wire [9:0] _meirotest_kekka_out206;
  wire [9:0] _meirotest_kekka_out207;
  wire [9:0] _meirotest_kekka_out208;
  wire [9:0] _meirotest_kekka_out209;
  wire [9:0] _meirotest_kekka_out210;
  wire [9:0] _meirotest_kekka_out211;
  wire [9:0] _meirotest_kekka_out212;
  wire [9:0] _meirotest_kekka_out213;
  wire [9:0] _meirotest_kekka_out214;
  wire [9:0] _meirotest_kekka_out215;
  wire [9:0] _meirotest_kekka_out216;
  wire [9:0] _meirotest_kekka_out217;
  wire [9:0] _meirotest_kekka_out218;
  wire [9:0] _meirotest_kekka_out219;
  wire [9:0] _meirotest_kekka_out220;
  wire [9:0] _meirotest_kekka_out221;
  wire [9:0] _meirotest_kekka_out222;
  wire _meirotest_in_do;
  wire _meirotest_end_meiro;
  wire _meirotest_p_reset;
  wire _meirotest_m_clock;
  wire _net_0;
  wire _net_1;
  wire _net_2;
  reg _reg_3;
  wire _net_4;
  wire _net_5;
  wire _net_6;
  wire _net_7;
  wire _net_8;
  wire _net_9;
  wire _net_10;
  wire _net_11;
  wire _net_12;
  wire _net_13;
  wire _net_14;
  wire _net_15;
  wire _net_16;
  wire _net_17;
  wire _net_18;
  wire _net_19;
  wire _net_20;
  wire _net_21;
  wire _net_22;
  wire _net_23;
  wire _net_24;
  wire _net_25;
  wire _net_26;
  wire _net_27;
  wire _net_28;
  wire _net_29;
  wire _net_30;
  wire _net_31;
  wire _net_32;
  wire _net_33;
  wire _net_34;
  wire _net_35;
  wire _net_36;
  wire _net_37;
  wire _net_38;
  wire _net_39;
  wire _net_40;
  wire _net_41;
  wire _net_42;
  wire _net_43;
  wire _net_44;
  wire _net_45;
  wire _net_46;
  wire _net_47;
  wire _net_48;
  wire _net_49;
  wire _net_50;
  wire _net_51;
  wire _net_52;
  wire _net_53;
  wire _net_54;
  wire _net_55;
  wire _net_56;
  wire _net_57;
  wire _net_58;
  wire _net_59;
  wire _net_60;
  wire _net_61;
  wire _net_62;
  wire _net_63;
  wire _net_64;
  wire _net_65;
  wire _net_66;
  wire _net_67;
  wire _net_68;
  wire _net_69;
  wire _net_70;
  wire _net_71;
  wire _net_72;
  wire _net_73;
  wire _net_74;
  wire _net_75;
  wire _net_76;
  wire _net_77;
  wire _net_78;
  wire _net_79;
  wire _net_80;
  wire _net_81;
  wire _net_82;
  wire _net_83;
  wire _net_84;
  wire _net_85;
  wire _net_86;
  wire _net_87;
  wire _net_88;
  wire _net_89;
  wire _net_90;
  wire _net_91;
  wire _net_92;
  wire _net_93;
  wire _net_94;
  wire _net_95;
  wire _net_96;
  wire _net_97;
  wire _net_98;
  wire _net_99;
  wire _net_100;
  wire _net_101;
  wire _net_102;
  wire _net_103;
  wire _net_104;
  wire _net_105;
  wire _net_106;
  wire _net_107;
  wire _net_108;
  wire _net_109;
  wire _net_110;
  wire _net_111;
  wire _net_112;
  wire _net_113;
  wire _net_114;
  wire _net_115;
  wire _net_116;
  wire _net_117;
  wire _net_118;
  wire _net_119;
  wire _net_120;
  wire _net_121;
  wire _net_122;
  wire _net_123;
  wire _net_124;
  wire _net_125;
  wire _net_126;
  wire _net_127;
  wire _net_128;
  wire _net_129;
  wire _net_130;
  wire _net_131;
  wire _net_132;
  wire _net_133;
  wire _net_134;
  wire _net_135;
  wire _net_136;
  wire _net_137;
  wire _net_138;
  wire _net_139;
  wire _net_140;
  wire _net_141;
  wire _net_142;
  wire _net_143;
  wire _net_144;
  wire _net_145;
  wire _net_146;
  wire _net_147;
  wire _net_148;
  wire _net_149;
  wire _net_150;
  wire _net_151;
  wire _net_152;
  wire _net_153;
  wire _net_154;
  wire _net_155;
  wire _net_156;
  wire _net_157;
  wire _net_158;
  wire _net_159;
  wire _net_160;
  wire _net_161;
  wire _net_162;
  wire _net_163;
  wire _net_164;
  wire _net_165;
  wire _net_166;
  wire _net_167;
  wire _net_168;
  wire _net_169;
  wire _net_170;
  wire _net_171;
  wire _net_172;
  wire _net_173;
  wire _net_174;
  wire _net_175;
  wire _net_176;
  wire _net_177;
  wire _net_178;
  wire _net_179;
  wire _net_180;
  wire _net_181;
  wire _net_182;
  wire _net_183;
  wire _net_184;
  wire _net_185;
  wire _net_186;
  wire _net_187;
  wire _net_188;
  wire _net_189;
  wire _net_190;
  wire _net_191;
  wire _net_192;
  wire _net_193;
  wire _net_194;
  wire _net_195;
  wire _net_196;
  wire _net_197;
  wire _net_198;
  wire _net_199;
  wire _net_200;
  wire _net_201;
  wire _net_202;
  wire _net_203;
  wire _net_204;
  wire _net_205;
  wire _net_206;
  wire _net_207;
  wire _net_208;
  wire _net_209;
  wire _net_210;
  wire _net_211;
  wire _net_212;
  wire _net_213;
  wire _net_214;
  wire _net_215;
  wire _net_216;
  wire _net_217;
  wire _net_218;
  wire _net_219;
  wire _net_220;
  wire _net_221;
  wire _net_222;
  wire _net_223;
  wire _net_224;
  wire _net_225;
  wire _net_226;
  wire _net_227;
  wire _net_228;
  wire _net_229;
  wire _net_230;
  wire _net_231;
  wire _net_232;
  wire _net_233;
  wire _net_234;
  wire _net_235;
  wire _net_236;
  wire _net_237;
  wire _net_238;
  wire _net_239;
  wire _net_240;
  wire _net_241;
  wire _net_242;
  wire _net_243;
  wire _net_244;
  wire _net_245;
  wire _net_246;
  wire _net_247;
  wire _net_248;
  wire _net_249;
  wire _net_250;
  wire _net_251;
  wire _net_252;
  wire _net_253;
  wire _net_254;
  wire _net_255;
  wire _net_256;
  wire _net_257;
  wire _net_258;
  wire _net_259;
  wire _net_260;
  wire _net_261;
  wire _net_262;
  wire _net_263;
  wire _net_264;
  wire _net_265;
  wire _net_266;
  wire _net_267;
  wire _net_268;
  wire _net_269;
  wire _net_270;
  wire _net_271;
  wire _net_272;
  wire _net_273;
  wire _net_274;
  wire _net_275;
  wire _net_276;
  wire _net_277;
  wire _net_278;
  wire _net_279;
  wire _net_280;
  wire _net_281;
  wire _net_282;
  wire _net_283;
  wire _net_284;
  wire _net_285;
  wire _net_286;
  wire _net_287;
  wire _net_288;
  wire _net_289;
  wire _net_290;
  wire _net_291;
  wire _net_292;
  wire _net_293;
  wire _net_294;
  wire _net_295;
  wire _net_296;
  wire _net_297;
  wire _net_298;
  wire _net_299;
  wire _net_300;
  wire _net_301;
  wire _net_302;
  wire _net_303;
  wire _net_304;
  wire _net_305;
  wire _net_306;
  wire _net_307;
  wire _net_308;
  wire _net_309;
  wire _net_310;
  wire _net_311;
  wire _net_312;
  wire _net_313;
  wire _net_314;
  wire _net_315;
  wire _net_316;
  wire _net_317;
  wire _net_318;
  wire _net_319;
  wire _net_320;
  wire _net_321;
  wire _net_322;
  wire _net_323;
  wire _net_324;
  wire _net_325;
  wire _net_326;
  wire _net_327;
  wire _net_328;
  wire _net_329;
  wire _net_330;
  wire _net_331;
  wire _net_332;
  wire _net_333;
  wire _net_334;
  wire _net_335;
  wire _net_336;
  wire _net_337;
  wire _net_338;
  wire _net_339;
  wire _net_340;
  wire _net_341;
  wire _net_342;
  wire _net_343;
  wire _net_344;
  wire _net_345;
  wire _net_346;
  wire _net_347;
  wire _net_348;
  wire _net_349;
  wire _net_350;
  wire _net_351;
  wire _net_352;
  wire _net_353;
  wire _net_354;
  wire _net_355;
  wire _net_356;
  wire _net_357;
  wire _net_358;
  wire _net_359;
  wire _net_360;
  wire _net_361;
  wire _net_362;
  wire _net_363;
  wire _net_364;
  wire _net_365;
  wire _net_366;
  wire _net_367;
  wire _net_368;
  wire _net_369;
  wire _net_370;
  wire _net_371;
  wire _net_372;
  wire _net_373;
  wire _net_374;
  wire _net_375;
  wire _net_376;
  wire _net_377;
  wire _net_378;
  wire _net_379;
  wire _net_380;
  wire _net_381;
  wire _net_382;
  wire _net_383;
  wire _net_384;
  wire _net_385;
  wire _net_386;
  wire _net_387;
  wire _net_388;
  wire _net_389;
  wire _net_390;
  wire _net_391;
  wire _net_392;
  wire _net_393;
  wire _net_394;
  wire _net_395;
  wire _net_396;
  wire _net_397;
  wire _net_398;
  wire _net_399;
  wire _net_400;
  wire _net_401;
  wire _net_402;
  wire _net_403;
  wire _net_404;
  wire _net_405;
  wire _net_406;
  wire _net_407;
  wire _net_408;
  wire _net_409;
  wire _net_410;
  wire _net_411;
  wire _net_412;
  wire _net_413;
  wire _net_414;
  wire _net_415;
  wire _net_416;
  wire _net_417;
  wire _net_418;
  wire _net_419;
  wire _net_420;
  wire _net_421;
  wire _net_422;
  wire _net_423;
  wire _net_424;
  wire _net_425;
  wire _net_426;
  wire _net_427;
  wire _net_428;
  wire _net_429;
  wire _net_430;
  wire _net_431;
  wire _net_432;
  wire _net_433;
  wire _net_434;
  wire _net_435;
  wire _net_436;
  wire _net_437;
  wire _net_438;
  wire _net_439;
  wire _net_440;
  wire _net_441;
  wire _net_442;
  wire _net_443;
  wire _net_444;
  wire _net_445;
  wire _net_446;
  wire _net_447;
  wire _net_448;
  wire _net_449;
  wire _net_450;
  wire _net_451;
  wire _net_452;
  wire _net_453;
  wire _net_454;
  wire _net_455;
  wire _net_456;
  wire _net_457;
  wire _net_458;
  wire _net_459;
  wire _net_460;
  wire _net_461;
  wire _net_462;
  wire _net_463;
  wire _net_464;
  wire _net_465;
  wire _net_466;
  wire _net_467;
  wire _net_468;
  wire _net_469;
  wire _net_470;
  wire _net_471;
  wire _net_472;
  wire _net_473;
  wire _net_474;
  wire _net_475;
  wire _net_476;
  wire _net_477;
  wire _net_478;
  wire _net_479;
  wire _net_480;
  wire _net_481;
  wire _net_482;
  wire _net_483;
  wire _net_484;
  wire _net_485;
  wire _net_486;
  wire _net_487;
  wire _net_488;
  wire _net_489;
  wire _net_490;
  wire _net_491;
  wire _net_492;
  wire _net_493;
  wire _net_494;
  wire _net_495;
  wire _net_496;
  wire _net_497;
  wire _net_498;
  wire _net_499;
  wire _net_500;
  wire _net_501;
  wire _net_502;
  wire _net_503;
  wire _net_504;
  wire _net_505;
  wire _net_506;
  wire _net_507;
  wire _net_508;
  wire _net_509;
  wire _net_510;
  wire _net_511;
  wire _net_512;
  wire _net_513;
  wire _net_514;
  wire _net_515;
  wire _net_516;
meiro meirotest (.m_clock(m_clock), .p_reset( p_reset), .end_meiro(_meirotest_end_meiro), .in_do(_meirotest_in_do), .kekka_out0(_meirotest_kekka_out0), .kekka_out1(_meirotest_kekka_out1), .kekka_out2(_meirotest_kekka_out2), .kekka_out3(_meirotest_kekka_out3), .kekka_out4(_meirotest_kekka_out4), .kekka_out5(_meirotest_kekka_out5), .kekka_out6(_meirotest_kekka_out6), .kekka_out7(_meirotest_kekka_out7), .kekka_out8(_meirotest_kekka_out8), .kekka_out9(_meirotest_kekka_out9), .kekka_out10(_meirotest_kekka_out10), .kekka_out11(_meirotest_kekka_out11), .kekka_out12(_meirotest_kekka_out12), .kekka_out13(_meirotest_kekka_out13), .kekka_out14(_meirotest_kekka_out14), .kekka_out15(_meirotest_kekka_out15), .kekka_out16(_meirotest_kekka_out16), .kekka_out17(_meirotest_kekka_out17), .kekka_out18(_meirotest_kekka_out18), .kekka_out19(_meirotest_kekka_out19), .kekka_out20(_meirotest_kekka_out20), .kekka_out21(_meirotest_kekka_out21), .kekka_out22(_meirotest_kekka_out22), .kekka_out23(_meirotest_kekka_out23), .kekka_out24(_meirotest_kekka_out24), .kekka_out25(_meirotest_kekka_out25), .kekka_out26(_meirotest_kekka_out26), .kekka_out27(_meirotest_kekka_out27), .kekka_out28(_meirotest_kekka_out28), .kekka_out29(_meirotest_kekka_out29), .kekka_out30(_meirotest_kekka_out30), .kekka_out31(_meirotest_kekka_out31), .kekka_out32(_meirotest_kekka_out32), .kekka_out33(_meirotest_kekka_out33), .kekka_out34(_meirotest_kekka_out34), .kekka_out35(_meirotest_kekka_out35), .kekka_out36(_meirotest_kekka_out36), .kekka_out37(_meirotest_kekka_out37), .kekka_out38(_meirotest_kekka_out38), .kekka_out39(_meirotest_kekka_out39), .kekka_out40(_meirotest_kekka_out40), .kekka_out41(_meirotest_kekka_out41), .kekka_out42(_meirotest_kekka_out42), .kekka_out43(_meirotest_kekka_out43), .kekka_out44(_meirotest_kekka_out44), .kekka_out45(_meirotest_kekka_out45), .kekka_out46(_meirotest_kekka_out46), .kekka_out47(_meirotest_kekka_out47), .kekka_out48(_meirotest_kekka_out48), .kekka_out49(_meirotest_kekka_out49), .kekka_out50(_meirotest_kekka_out50), .kekka_out51(_meirotest_kekka_out51), .kekka_out52(_meirotest_kekka_out52), .kekka_out53(_meirotest_kekka_out53), .kekka_out54(_meirotest_kekka_out54), .kekka_out55(_meirotest_kekka_out55), .kekka_out56(_meirotest_kekka_out56), .kekka_out57(_meirotest_kekka_out57), .kekka_out58(_meirotest_kekka_out58), .kekka_out59(_meirotest_kekka_out59), .kekka_out60(_meirotest_kekka_out60), .kekka_out61(_meirotest_kekka_out61), .kekka_out62(_meirotest_kekka_out62), .kekka_out63(_meirotest_kekka_out63), .kekka_out64(_meirotest_kekka_out64), .kekka_out65(_meirotest_kekka_out65), .kekka_out66(_meirotest_kekka_out66), .kekka_out67(_meirotest_kekka_out67), .kekka_out68(_meirotest_kekka_out68), .kekka_out69(_meirotest_kekka_out69), .kekka_out70(_meirotest_kekka_out70), .kekka_out71(_meirotest_kekka_out71), .kekka_out72(_meirotest_kekka_out72), .kekka_out73(_meirotest_kekka_out73), .kekka_out74(_meirotest_kekka_out74), .kekka_out75(_meirotest_kekka_out75), .kekka_out76(_meirotest_kekka_out76), .kekka_out77(_meirotest_kekka_out77), .kekka_out78(_meirotest_kekka_out78), .kekka_out79(_meirotest_kekka_out79), .kekka_out80(_meirotest_kekka_out80), .kekka_out81(_meirotest_kekka_out81), .kekka_out82(_meirotest_kekka_out82), .kekka_out83(_meirotest_kekka_out83), .kekka_out84(_meirotest_kekka_out84), .kekka_out85(_meirotest_kekka_out85), .kekka_out86(_meirotest_kekka_out86), .kekka_out87(_meirotest_kekka_out87), .kekka_out88(_meirotest_kekka_out88), .kekka_out89(_meirotest_kekka_out89), .kekka_out90(_meirotest_kekka_out90), .kekka_out91(_meirotest_kekka_out91), .kekka_out92(_meirotest_kekka_out92), .kekka_out93(_meirotest_kekka_out93), .kekka_out94(_meirotest_kekka_out94), .kekka_out95(_meirotest_kekka_out95), .kekka_out96(_meirotest_kekka_out96), .kekka_out97(_meirotest_kekka_out97), .kekka_out98(_meirotest_kekka_out98), .kekka_out99(_meirotest_kekka_out99), .kekka_out100(_meirotest_kekka_out100), .kekka_out101(_meirotest_kekka_out101), .kekka_out102(_meirotest_kekka_out102), .kekka_out103(_meirotest_kekka_out103), .kekka_out104(_meirotest_kekka_out104), .kekka_out105(_meirotest_kekka_out105), .kekka_out106(_meirotest_kekka_out106), .kekka_out107(_meirotest_kekka_out107), .kekka_out108(_meirotest_kekka_out108), .kekka_out109(_meirotest_kekka_out109), .kekka_out110(_meirotest_kekka_out110), .kekka_out111(_meirotest_kekka_out111), .kekka_out112(_meirotest_kekka_out112), .kekka_out113(_meirotest_kekka_out113), .kekka_out114(_meirotest_kekka_out114), .kekka_out115(_meirotest_kekka_out115), .kekka_out116(_meirotest_kekka_out116), .kekka_out117(_meirotest_kekka_out117), .kekka_out118(_meirotest_kekka_out118), .kekka_out119(_meirotest_kekka_out119), .kekka_out120(_meirotest_kekka_out120), .kekka_out121(_meirotest_kekka_out121), .kekka_out122(_meirotest_kekka_out122), .kekka_out123(_meirotest_kekka_out123), .kekka_out124(_meirotest_kekka_out124), .kekka_out125(_meirotest_kekka_out125), .kekka_out126(_meirotest_kekka_out126), .kekka_out127(_meirotest_kekka_out127), .kekka_out128(_meirotest_kekka_out128), .kekka_out129(_meirotest_kekka_out129), .kekka_out130(_meirotest_kekka_out130), .kekka_out131(_meirotest_kekka_out131), .kekka_out132(_meirotest_kekka_out132), .kekka_out133(_meirotest_kekka_out133), .kekka_out134(_meirotest_kekka_out134), .kekka_out135(_meirotest_kekka_out135), .kekka_out136(_meirotest_kekka_out136), .kekka_out137(_meirotest_kekka_out137), .kekka_out138(_meirotest_kekka_out138), .kekka_out139(_meirotest_kekka_out139), .kekka_out140(_meirotest_kekka_out140), .kekka_out141(_meirotest_kekka_out141), .kekka_out142(_meirotest_kekka_out142), .kekka_out143(_meirotest_kekka_out143), .kekka_out144(_meirotest_kekka_out144), .kekka_out145(_meirotest_kekka_out145), .kekka_out146(_meirotest_kekka_out146), .kekka_out147(_meirotest_kekka_out147), .kekka_out148(_meirotest_kekka_out148), .kekka_out149(_meirotest_kekka_out149), .kekka_out150(_meirotest_kekka_out150), .kekka_out151(_meirotest_kekka_out151), .kekka_out152(_meirotest_kekka_out152), .kekka_out153(_meirotest_kekka_out153), .kekka_out154(_meirotest_kekka_out154), .kekka_out155(_meirotest_kekka_out155), .kekka_out156(_meirotest_kekka_out156), .kekka_out157(_meirotest_kekka_out157), .kekka_out158(_meirotest_kekka_out158), .kekka_out159(_meirotest_kekka_out159), .kekka_out160(_meirotest_kekka_out160), .kekka_out161(_meirotest_kekka_out161), .kekka_out162(_meirotest_kekka_out162), .kekka_out163(_meirotest_kekka_out163), .kekka_out164(_meirotest_kekka_out164), .kekka_out165(_meirotest_kekka_out165), .kekka_out166(_meirotest_kekka_out166), .kekka_out167(_meirotest_kekka_out167), .kekka_out168(_meirotest_kekka_out168), .kekka_out169(_meirotest_kekka_out169), .kekka_out170(_meirotest_kekka_out170), .kekka_out171(_meirotest_kekka_out171), .kekka_out172(_meirotest_kekka_out172), .kekka_out173(_meirotest_kekka_out173), .kekka_out174(_meirotest_kekka_out174), .kekka_out175(_meirotest_kekka_out175), .kekka_out176(_meirotest_kekka_out176), .kekka_out177(_meirotest_kekka_out177), .kekka_out178(_meirotest_kekka_out178), .kekka_out179(_meirotest_kekka_out179), .kekka_out180(_meirotest_kekka_out180), .kekka_out181(_meirotest_kekka_out181), .kekka_out182(_meirotest_kekka_out182), .kekka_out183(_meirotest_kekka_out183), .kekka_out184(_meirotest_kekka_out184), .kekka_out185(_meirotest_kekka_out185), .kekka_out186(_meirotest_kekka_out186), .kekka_out187(_meirotest_kekka_out187), .kekka_out188(_meirotest_kekka_out188), .kekka_out189(_meirotest_kekka_out189), .kekka_out190(_meirotest_kekka_out190), .kekka_out191(_meirotest_kekka_out191), .kekka_out192(_meirotest_kekka_out192), .kekka_out193(_meirotest_kekka_out193), .kekka_out194(_meirotest_kekka_out194), .kekka_out195(_meirotest_kekka_out195), .kekka_out196(_meirotest_kekka_out196), .kekka_out197(_meirotest_kekka_out197), .kekka_out198(_meirotest_kekka_out198), .kekka_out199(_meirotest_kekka_out199), .kekka_out200(_meirotest_kekka_out200), .kekka_out201(_meirotest_kekka_out201), .kekka_out202(_meirotest_kekka_out202), .kekka_out203(_meirotest_kekka_out203), .kekka_out204(_meirotest_kekka_out204), .kekka_out205(_meirotest_kekka_out205), .kekka_out206(_meirotest_kekka_out206), .kekka_out207(_meirotest_kekka_out207), .kekka_out208(_meirotest_kekka_out208), .kekka_out209(_meirotest_kekka_out209), .kekka_out210(_meirotest_kekka_out210), .kekka_out211(_meirotest_kekka_out211), .kekka_out212(_meirotest_kekka_out212), .kekka_out213(_meirotest_kekka_out213), .kekka_out214(_meirotest_kekka_out214), .kekka_out215(_meirotest_kekka_out215), .kekka_out216(_meirotest_kekka_out216), .kekka_out217(_meirotest_kekka_out217), .kekka_out218(_meirotest_kekka_out218), .kekka_out219(_meirotest_kekka_out219), .kekka_out220(_meirotest_kekka_out220), .kekka_out221(_meirotest_kekka_out221), .kekka_out222(_meirotest_kekka_out222), .map_value_arg0(_meirotest_map_value_arg0), .map_value_arg1(_meirotest_map_value_arg1), .map_value_arg2(_meirotest_map_value_arg2), .map_value_arg3(_meirotest_map_value_arg3), .map_value_arg4(_meirotest_map_value_arg4), .map_value_arg5(_meirotest_map_value_arg5), .map_value_arg6(_meirotest_map_value_arg6), .map_value_arg7(_meirotest_map_value_arg7), .map_value_arg8(_meirotest_map_value_arg8), .map_value_arg9(_meirotest_map_value_arg9), .map_value_arg10(_meirotest_map_value_arg10), .map_value_arg11(_meirotest_map_value_arg11), .map_value_arg12(_meirotest_map_value_arg12), .map_value_arg13(_meirotest_map_value_arg13), .map_value_arg14(_meirotest_map_value_arg14), .map_value_arg15(_meirotest_map_value_arg15), .map_value_arg16(_meirotest_map_value_arg16), .map_value_arg17(_meirotest_map_value_arg17), .map_value_arg18(_meirotest_map_value_arg18), .map_value_arg19(_meirotest_map_value_arg19), .map_value_arg20(_meirotest_map_value_arg20), .map_value_arg21(_meirotest_map_value_arg21), .map_value_arg22(_meirotest_map_value_arg22), .map_value_arg23(_meirotest_map_value_arg23), .map_value_arg24(_meirotest_map_value_arg24), .map_value_arg25(_meirotest_map_value_arg25), .map_value_arg26(_meirotest_map_value_arg26), .map_value_arg27(_meirotest_map_value_arg27), .map_value_arg28(_meirotest_map_value_arg28), .map_value_arg29(_meirotest_map_value_arg29), .map_value_arg30(_meirotest_map_value_arg30), .map_value_arg31(_meirotest_map_value_arg31), .map_value_arg32(_meirotest_map_value_arg32), .map_value_arg33(_meirotest_map_value_arg33), .map_value_arg34(_meirotest_map_value_arg34), .map_value_arg35(_meirotest_map_value_arg35), .map_value_arg36(_meirotest_map_value_arg36), .map_value_arg37(_meirotest_map_value_arg37), .map_value_arg38(_meirotest_map_value_arg38), .map_value_arg39(_meirotest_map_value_arg39), .map_value_arg40(_meirotest_map_value_arg40), .map_value_arg41(_meirotest_map_value_arg41), .map_value_arg42(_meirotest_map_value_arg42), .map_value_arg43(_meirotest_map_value_arg43), .map_value_arg44(_meirotest_map_value_arg44), .map_value_arg45(_meirotest_map_value_arg45), .map_value_arg46(_meirotest_map_value_arg46), .map_value_arg47(_meirotest_map_value_arg47), .map_value_arg48(_meirotest_map_value_arg48), .map_value_arg49(_meirotest_map_value_arg49), .map_value_arg50(_meirotest_map_value_arg50), .map_value_arg51(_meirotest_map_value_arg51), .map_value_arg52(_meirotest_map_value_arg52), .map_value_arg53(_meirotest_map_value_arg53), .map_value_arg54(_meirotest_map_value_arg54), .map_value_arg55(_meirotest_map_value_arg55), .map_value_arg56(_meirotest_map_value_arg56), .map_value_arg57(_meirotest_map_value_arg57), .map_value_arg58(_meirotest_map_value_arg58), .map_value_arg59(_meirotest_map_value_arg59), .map_value_arg60(_meirotest_map_value_arg60), .map_value_arg61(_meirotest_map_value_arg61), .map_value_arg62(_meirotest_map_value_arg62), .map_value_arg63(_meirotest_map_value_arg63), .map_value_arg64(_meirotest_map_value_arg64), .map_value_arg65(_meirotest_map_value_arg65), .map_value_arg66(_meirotest_map_value_arg66), .map_value_arg67(_meirotest_map_value_arg67), .map_value_arg68(_meirotest_map_value_arg68), .map_value_arg69(_meirotest_map_value_arg69), .map_value_arg70(_meirotest_map_value_arg70), .map_value_arg71(_meirotest_map_value_arg71), .map_value_arg72(_meirotest_map_value_arg72), .map_value_arg73(_meirotest_map_value_arg73), .map_value_arg74(_meirotest_map_value_arg74), .map_value_arg75(_meirotest_map_value_arg75), .map_value_arg76(_meirotest_map_value_arg76), .map_value_arg77(_meirotest_map_value_arg77), .map_value_arg78(_meirotest_map_value_arg78), .map_value_arg79(_meirotest_map_value_arg79), .map_value_arg80(_meirotest_map_value_arg80), .map_value_arg81(_meirotest_map_value_arg81), .map_value_arg82(_meirotest_map_value_arg82), .map_value_arg83(_meirotest_map_value_arg83), .map_value_arg84(_meirotest_map_value_arg84), .map_value_arg85(_meirotest_map_value_arg85), .map_value_arg86(_meirotest_map_value_arg86), .map_value_arg87(_meirotest_map_value_arg87), .map_value_arg88(_meirotest_map_value_arg88), .map_value_arg89(_meirotest_map_value_arg89), .map_value_arg90(_meirotest_map_value_arg90), .map_value_arg91(_meirotest_map_value_arg91), .map_value_arg92(_meirotest_map_value_arg92), .map_value_arg93(_meirotest_map_value_arg93), .map_value_arg94(_meirotest_map_value_arg94), .map_value_arg95(_meirotest_map_value_arg95), .map_value_arg96(_meirotest_map_value_arg96), .map_value_arg97(_meirotest_map_value_arg97), .map_value_arg98(_meirotest_map_value_arg98), .map_value_arg99(_meirotest_map_value_arg99), .map_value_arg100(_meirotest_map_value_arg100), .map_value_arg101(_meirotest_map_value_arg101), .map_value_arg102(_meirotest_map_value_arg102), .map_value_arg103(_meirotest_map_value_arg103), .map_value_arg104(_meirotest_map_value_arg104), .map_value_arg105(_meirotest_map_value_arg105), .map_value_arg106(_meirotest_map_value_arg106), .map_value_arg107(_meirotest_map_value_arg107), .map_value_arg108(_meirotest_map_value_arg108), .map_value_arg109(_meirotest_map_value_arg109), .map_value_arg110(_meirotest_map_value_arg110), .map_value_arg111(_meirotest_map_value_arg111), .map_value_arg112(_meirotest_map_value_arg112), .map_value_arg113(_meirotest_map_value_arg113), .map_value_arg114(_meirotest_map_value_arg114), .map_value_arg115(_meirotest_map_value_arg115), .map_value_arg116(_meirotest_map_value_arg116), .map_value_arg117(_meirotest_map_value_arg117), .map_value_arg118(_meirotest_map_value_arg118), .map_value_arg119(_meirotest_map_value_arg119), .map_value_arg120(_meirotest_map_value_arg120), .map_value_arg121(_meirotest_map_value_arg121), .map_value_arg122(_meirotest_map_value_arg122), .map_value_arg123(_meirotest_map_value_arg123), .map_value_arg124(_meirotest_map_value_arg124), .map_value_arg125(_meirotest_map_value_arg125), .map_value_arg126(_meirotest_map_value_arg126), .map_value_arg127(_meirotest_map_value_arg127), .map_value_arg128(_meirotest_map_value_arg128), .map_value_arg129(_meirotest_map_value_arg129), .map_value_arg130(_meirotest_map_value_arg130), .map_value_arg131(_meirotest_map_value_arg131), .map_value_arg132(_meirotest_map_value_arg132), .map_value_arg133(_meirotest_map_value_arg133), .map_value_arg134(_meirotest_map_value_arg134), .map_value_arg135(_meirotest_map_value_arg135), .map_value_arg136(_meirotest_map_value_arg136), .map_value_arg137(_meirotest_map_value_arg137), .map_value_arg138(_meirotest_map_value_arg138), .map_value_arg139(_meirotest_map_value_arg139), .map_value_arg140(_meirotest_map_value_arg140), .map_value_arg141(_meirotest_map_value_arg141), .map_value_arg142(_meirotest_map_value_arg142), .map_value_arg143(_meirotest_map_value_arg143), .map_value_arg144(_meirotest_map_value_arg144), .map_value_arg145(_meirotest_map_value_arg145), .map_value_arg146(_meirotest_map_value_arg146), .map_value_arg147(_meirotest_map_value_arg147), .map_value_arg148(_meirotest_map_value_arg148), .map_value_arg149(_meirotest_map_value_arg149), .map_value_arg150(_meirotest_map_value_arg150), .map_value_arg151(_meirotest_map_value_arg151), .map_value_arg152(_meirotest_map_value_arg152), .map_value_arg153(_meirotest_map_value_arg153), .map_value_arg154(_meirotest_map_value_arg154), .map_value_arg155(_meirotest_map_value_arg155), .map_value_arg156(_meirotest_map_value_arg156), .map_value_arg157(_meirotest_map_value_arg157), .map_value_arg158(_meirotest_map_value_arg158), .map_value_arg159(_meirotest_map_value_arg159), .map_value_arg160(_meirotest_map_value_arg160), .map_value_arg161(_meirotest_map_value_arg161), .map_value_arg162(_meirotest_map_value_arg162), .map_value_arg163(_meirotest_map_value_arg163), .map_value_arg164(_meirotest_map_value_arg164), .map_value_arg165(_meirotest_map_value_arg165), .map_value_arg166(_meirotest_map_value_arg166), .map_value_arg167(_meirotest_map_value_arg167), .map_value_arg168(_meirotest_map_value_arg168), .map_value_arg169(_meirotest_map_value_arg169), .map_value_arg170(_meirotest_map_value_arg170), .map_value_arg171(_meirotest_map_value_arg171), .map_value_arg172(_meirotest_map_value_arg172), .map_value_arg173(_meirotest_map_value_arg173), .map_value_arg174(_meirotest_map_value_arg174), .map_value_arg175(_meirotest_map_value_arg175), .map_value_arg176(_meirotest_map_value_arg176), .map_value_arg177(_meirotest_map_value_arg177), .map_value_arg178(_meirotest_map_value_arg178), .map_value_arg179(_meirotest_map_value_arg179), .map_value_arg180(_meirotest_map_value_arg180), .map_value_arg181(_meirotest_map_value_arg181), .map_value_arg182(_meirotest_map_value_arg182), .map_value_arg183(_meirotest_map_value_arg183), .map_value_arg184(_meirotest_map_value_arg184), .map_value_arg185(_meirotest_map_value_arg185), .map_value_arg186(_meirotest_map_value_arg186), .map_value_arg187(_meirotest_map_value_arg187), .map_value_arg188(_meirotest_map_value_arg188), .map_value_arg189(_meirotest_map_value_arg189), .map_value_arg190(_meirotest_map_value_arg190), .map_value_arg191(_meirotest_map_value_arg191), .map_value_arg192(_meirotest_map_value_arg192), .map_value_arg193(_meirotest_map_value_arg193), .map_value_arg194(_meirotest_map_value_arg194), .map_value_arg195(_meirotest_map_value_arg195), .map_value_arg196(_meirotest_map_value_arg196), .map_value_arg197(_meirotest_map_value_arg197), .map_value_arg198(_meirotest_map_value_arg198), .map_value_arg199(_meirotest_map_value_arg199), .map_value_arg200(_meirotest_map_value_arg200), .map_value_arg201(_meirotest_map_value_arg201), .map_value_arg202(_meirotest_map_value_arg202), .map_value_arg203(_meirotest_map_value_arg203), .map_value_arg204(_meirotest_map_value_arg204), .map_value_arg205(_meirotest_map_value_arg205), .map_value_arg206(_meirotest_map_value_arg206), .map_value_arg207(_meirotest_map_value_arg207), .map_value_arg208(_meirotest_map_value_arg208), .map_value_arg209(_meirotest_map_value_arg209), .map_value_arg210(_meirotest_map_value_arg210), .map_value_arg211(_meirotest_map_value_arg211), .map_value_arg212(_meirotest_map_value_arg212), .map_value_arg213(_meirotest_map_value_arg213), .map_value_arg214(_meirotest_map_value_arg214), .map_value_arg215(_meirotest_map_value_arg215), .map_value_arg216(_meirotest_map_value_arg216), .map_value_arg217(_meirotest_map_value_arg217), .map_value_arg218(_meirotest_map_value_arg218), .map_value_arg219(_meirotest_map_value_arg219), .map_value_arg220(_meirotest_map_value_arg220), .map_value_arg221(_meirotest_map_value_arg221), .map_value_arg222(_meirotest_map_value_arg222), .map_value_arg223(_meirotest_map_value_arg223), .map_value_arg224(_meirotest_map_value_arg224), .map_value_arg225(_meirotest_map_value_arg225), .map_value_arg226(_meirotest_map_value_arg226), .map_value_arg227(_meirotest_map_value_arg227), .map_value_arg228(_meirotest_map_value_arg228), .map_value_arg229(_meirotest_map_value_arg229), .map_value_arg230(_meirotest_map_value_arg230), .map_value_arg231(_meirotest_map_value_arg231), .map_value_arg232(_meirotest_map_value_arg232), .map_value_arg233(_meirotest_map_value_arg233), .map_value_arg234(_meirotest_map_value_arg234), .map_value_arg235(_meirotest_map_value_arg235), .map_value_arg236(_meirotest_map_value_arg236), .map_value_arg237(_meirotest_map_value_arg237), .map_value_arg238(_meirotest_map_value_arg238), .map_value_arg239(_meirotest_map_value_arg239), .map_value_arg240(_meirotest_map_value_arg240), .map_value_arg241(_meirotest_map_value_arg241), .map_value_arg242(_meirotest_map_value_arg242), .map_value_arg243(_meirotest_map_value_arg243), .map_value_arg244(_meirotest_map_value_arg244), .map_value_arg245(_meirotest_map_value_arg245), .map_value_arg246(_meirotest_map_value_arg246), .map_value_arg247(_meirotest_map_value_arg247), .map_value_arg248(_meirotest_map_value_arg248), .map_value_arg249(_meirotest_map_value_arg249), .map_value_arg250(_meirotest_map_value_arg250), .map_value_arg251(_meirotest_map_value_arg251), .map_value_arg252(_meirotest_map_value_arg252), .map_value_arg253(_meirotest_map_value_arg253), .map_value_arg254(_meirotest_map_value_arg254), .map_value_arg255(_meirotest_map_value_arg255), .map_value_arg256(_meirotest_map_value_arg256), .map_value_arg257(_meirotest_map_value_arg257), .map_value_arg258(_meirotest_map_value_arg258), .map_value_arg259(_meirotest_map_value_arg259), .map_value_arg260(_meirotest_map_value_arg260), .map_value_arg261(_meirotest_map_value_arg261), .map_value_arg262(_meirotest_map_value_arg262), .map_value_arg263(_meirotest_map_value_arg263), .map_value_arg264(_meirotest_map_value_arg264), .map_value_arg265(_meirotest_map_value_arg265), .map_value_arg266(_meirotest_map_value_arg266), .map_value_arg267(_meirotest_map_value_arg267), .map_value_arg268(_meirotest_map_value_arg268), .map_value_arg269(_meirotest_map_value_arg269), .map_value_arg270(_meirotest_map_value_arg270), .map_value_arg271(_meirotest_map_value_arg271), .map_value_arg272(_meirotest_map_value_arg272), .map_value_arg273(_meirotest_map_value_arg273), .map_value_arg274(_meirotest_map_value_arg274), .map_value_arg275(_meirotest_map_value_arg275), .map_value_arg276(_meirotest_map_value_arg276), .map_value_arg277(_meirotest_map_value_arg277), .map_value_arg278(_meirotest_map_value_arg278), .map_value_arg279(_meirotest_map_value_arg279), .map_value_arg280(_meirotest_map_value_arg280), .map_value_arg281(_meirotest_map_value_arg281), .map_value_arg282(_meirotest_map_value_arg282), .map_value_arg283(_meirotest_map_value_arg283), .map_value_arg284(_meirotest_map_value_arg284), .map_value_arg285(_meirotest_map_value_arg285), .map_value_arg286(_meirotest_map_value_arg286), .map_value_arg287(_meirotest_map_value_arg287), .map_value_arg288(_meirotest_map_value_arg288), .map_value_arg289(_meirotest_map_value_arg289), .map_value_arg290(_meirotest_map_value_arg290), .map_value_arg291(_meirotest_map_value_arg291), .map_value_arg292(_meirotest_map_value_arg292), .map_value_arg293(_meirotest_map_value_arg293), .map_value_arg294(_meirotest_map_value_arg294), .map_value_arg295(_meirotest_map_value_arg295), .map_value_arg296(_meirotest_map_value_arg296), .map_value_arg297(_meirotest_map_value_arg297), .map_value_arg298(_meirotest_map_value_arg298), .map_value_arg299(_meirotest_map_value_arg299), .map_value_arg300(_meirotest_map_value_arg300), .map_value_arg301(_meirotest_map_value_arg301), .map_value_arg302(_meirotest_map_value_arg302), .map_value_arg303(_meirotest_map_value_arg303), .map_value_arg304(_meirotest_map_value_arg304), .map_value_arg305(_meirotest_map_value_arg305), .map_value_arg306(_meirotest_map_value_arg306), .map_value_arg307(_meirotest_map_value_arg307), .map_value_arg308(_meirotest_map_value_arg308), .map_value_arg309(_meirotest_map_value_arg309), .map_value_arg310(_meirotest_map_value_arg310), .map_value_arg311(_meirotest_map_value_arg311), .map_value_arg312(_meirotest_map_value_arg312), .map_value_arg313(_meirotest_map_value_arg313), .map_value_arg314(_meirotest_map_value_arg314), .map_value_arg315(_meirotest_map_value_arg315), .map_value_arg316(_meirotest_map_value_arg316), .map_value_arg317(_meirotest_map_value_arg317), .map_value_arg318(_meirotest_map_value_arg318), .map_value_arg319(_meirotest_map_value_arg319), .map_value_arg320(_meirotest_map_value_arg320), .map_value_arg321(_meirotest_map_value_arg321), .map_value_arg322(_meirotest_map_value_arg322), .map_value_arg323(_meirotest_map_value_arg323), .map_value_arg324(_meirotest_map_value_arg324), .map_value_arg325(_meirotest_map_value_arg325), .map_value_arg326(_meirotest_map_value_arg326), .map_value_arg327(_meirotest_map_value_arg327), .map_value_arg328(_meirotest_map_value_arg328), .map_value_arg329(_meirotest_map_value_arg329), .map_value_arg330(_meirotest_map_value_arg330), .map_value_arg331(_meirotest_map_value_arg331), .map_value_arg332(_meirotest_map_value_arg332), .map_value_arg333(_meirotest_map_value_arg333), .map_value_arg334(_meirotest_map_value_arg334), .map_value_arg335(_meirotest_map_value_arg335), .map_value_arg336(_meirotest_map_value_arg336), .map_value_arg337(_meirotest_map_value_arg337), .map_value_arg338(_meirotest_map_value_arg338), .map_value_arg339(_meirotest_map_value_arg339), .map_value_arg340(_meirotest_map_value_arg340), .map_value_arg341(_meirotest_map_value_arg341), .map_value_arg342(_meirotest_map_value_arg342), .map_value_arg343(_meirotest_map_value_arg343), .map_value_arg344(_meirotest_map_value_arg344), .map_value_arg345(_meirotest_map_value_arg345), .map_value_arg346(_meirotest_map_value_arg346), .map_value_arg347(_meirotest_map_value_arg347), .map_value_arg348(_meirotest_map_value_arg348), .map_value_arg349(_meirotest_map_value_arg349), .map_value_arg350(_meirotest_map_value_arg350), .map_value_arg351(_meirotest_map_value_arg351), .map_value_arg352(_meirotest_map_value_arg352), .map_value_arg353(_meirotest_map_value_arg353), .map_value_arg354(_meirotest_map_value_arg354), .map_value_arg355(_meirotest_map_value_arg355), .map_value_arg356(_meirotest_map_value_arg356), .map_value_arg357(_meirotest_map_value_arg357), .map_value_arg358(_meirotest_map_value_arg358), .map_value_arg359(_meirotest_map_value_arg359), .map_value_arg360(_meirotest_map_value_arg360), .map_value_arg361(_meirotest_map_value_arg361), .map_value_arg362(_meirotest_map_value_arg362), .map_value_arg363(_meirotest_map_value_arg363), .map_value_arg364(_meirotest_map_value_arg364), .map_value_arg365(_meirotest_map_value_arg365), .map_value_arg366(_meirotest_map_value_arg366), .map_value_arg367(_meirotest_map_value_arg367), .map_value_arg368(_meirotest_map_value_arg368), .map_value_arg369(_meirotest_map_value_arg369), .map_value_arg370(_meirotest_map_value_arg370), .map_value_arg371(_meirotest_map_value_arg371), .map_value_arg372(_meirotest_map_value_arg372), .map_value_arg373(_meirotest_map_value_arg373), .map_value_arg374(_meirotest_map_value_arg374), .map_value_arg375(_meirotest_map_value_arg375), .map_value_arg376(_meirotest_map_value_arg376), .map_value_arg377(_meirotest_map_value_arg377), .map_value_arg378(_meirotest_map_value_arg378), .map_value_arg379(_meirotest_map_value_arg379), .map_value_arg380(_meirotest_map_value_arg380), .map_value_arg381(_meirotest_map_value_arg381), .map_value_arg382(_meirotest_map_value_arg382), .map_value_arg383(_meirotest_map_value_arg383), .map_value_arg384(_meirotest_map_value_arg384), .map_value_arg385(_meirotest_map_value_arg385), .map_value_arg386(_meirotest_map_value_arg386), .map_value_arg387(_meirotest_map_value_arg387), .map_value_arg388(_meirotest_map_value_arg388), .map_value_arg389(_meirotest_map_value_arg389), .map_value_arg390(_meirotest_map_value_arg390), .map_value_arg391(_meirotest_map_value_arg391), .map_value_arg392(_meirotest_map_value_arg392), .map_value_arg393(_meirotest_map_value_arg393), .map_value_arg394(_meirotest_map_value_arg394), .map_value_arg395(_meirotest_map_value_arg395), .map_value_arg396(_meirotest_map_value_arg396), .map_value_arg397(_meirotest_map_value_arg397), .map_value_arg398(_meirotest_map_value_arg398), .map_value_arg399(_meirotest_map_value_arg399), .map_value_arg400(_meirotest_map_value_arg400), .map_value_arg401(_meirotest_map_value_arg401), .map_value_arg402(_meirotest_map_value_arg402), .map_value_arg403(_meirotest_map_value_arg403), .map_value_arg404(_meirotest_map_value_arg404), .map_value_arg405(_meirotest_map_value_arg405), .map_value_arg406(_meirotest_map_value_arg406), .map_value_arg407(_meirotest_map_value_arg407), .map_value_arg408(_meirotest_map_value_arg408), .map_value_arg409(_meirotest_map_value_arg409), .map_value_arg410(_meirotest_map_value_arg410), .map_value_arg411(_meirotest_map_value_arg411), .map_value_arg412(_meirotest_map_value_arg412), .map_value_arg413(_meirotest_map_value_arg413), .map_value_arg414(_meirotest_map_value_arg414), .map_value_arg415(_meirotest_map_value_arg415), .map_value_arg416(_meirotest_map_value_arg416), .map_value_arg417(_meirotest_map_value_arg417), .map_value_arg418(_meirotest_map_value_arg418), .map_value_arg419(_meirotest_map_value_arg419), .map_value_arg420(_meirotest_map_value_arg420), .map_value_arg421(_meirotest_map_value_arg421), .map_value_arg422(_meirotest_map_value_arg422), .map_value_arg423(_meirotest_map_value_arg423), .map_value_arg424(_meirotest_map_value_arg424), .map_value_arg425(_meirotest_map_value_arg425), .map_value_arg426(_meirotest_map_value_arg426), .map_value_arg427(_meirotest_map_value_arg427), .map_value_arg428(_meirotest_map_value_arg428), .map_value_arg429(_meirotest_map_value_arg429), .map_value_arg430(_meirotest_map_value_arg430), .map_value_arg431(_meirotest_map_value_arg431), .map_value_arg432(_meirotest_map_value_arg432), .map_value_arg433(_meirotest_map_value_arg433), .map_value_arg434(_meirotest_map_value_arg434), .map_value_arg435(_meirotest_map_value_arg435), .map_value_arg436(_meirotest_map_value_arg436), .map_value_arg437(_meirotest_map_value_arg437), .map_value_arg438(_meirotest_map_value_arg438), .map_value_arg439(_meirotest_map_value_arg439), .map_value_arg440(_meirotest_map_value_arg440), .map_value_arg441(_meirotest_map_value_arg441), .map_value_arg442(_meirotest_map_value_arg442), .map_value_arg443(_meirotest_map_value_arg443), .map_value_arg444(_meirotest_map_value_arg444), .map_value_arg445(_meirotest_map_value_arg445), .map_value_arg446(_meirotest_map_value_arg446), .map_value_arg447(_meirotest_map_value_arg447), .map_value_arg448(_meirotest_map_value_arg448), .map_value_arg449(_meirotest_map_value_arg449), .map_value_arg450(_meirotest_map_value_arg450), .map_value_arg451(_meirotest_map_value_arg451), .map_value_arg452(_meirotest_map_value_arg452), .map_value_arg453(_meirotest_map_value_arg453), .map_value_arg454(_meirotest_map_value_arg454), .map_value_arg455(_meirotest_map_value_arg455), .map_value_arg456(_meirotest_map_value_arg456), .map_value_arg457(_meirotest_map_value_arg457), .map_value_arg458(_meirotest_map_value_arg458), .map_value_arg459(_meirotest_map_value_arg459), .map_value_arg460(_meirotest_map_value_arg460), .map_value_arg461(_meirotest_map_value_arg461), .map_value_arg462(_meirotest_map_value_arg462), .map_value_arg463(_meirotest_map_value_arg463), .map_value_arg464(_meirotest_map_value_arg464), .map_value_arg465(_meirotest_map_value_arg465), .map_value_arg466(_meirotest_map_value_arg466), .map_value_arg467(_meirotest_map_value_arg467), .map_value_arg468(_meirotest_map_value_arg468), .map_value_arg469(_meirotest_map_value_arg469), .map_value_arg470(_meirotest_map_value_arg470), .map_value_arg471(_meirotest_map_value_arg471), .map_value_arg472(_meirotest_map_value_arg472), .map_value_arg473(_meirotest_map_value_arg473), .map_value_arg474(_meirotest_map_value_arg474), .map_value_arg475(_meirotest_map_value_arg475), .map_value_arg476(_meirotest_map_value_arg476), .map_value_arg477(_meirotest_map_value_arg477), .map_value_arg478(_meirotest_map_value_arg478), .map_value_arg479(_meirotest_map_value_arg479), .map_value_arg480(_meirotest_map_value_arg480), .map_value_arg481(_meirotest_map_value_arg481), .map_value_arg482(_meirotest_map_value_arg482), .map_value_arg483(_meirotest_map_value_arg483), .map_value_arg484(_meirotest_map_value_arg484), .map_value_arg485(_meirotest_map_value_arg485), .map_value_arg486(_meirotest_map_value_arg486), .map_value_arg487(_meirotest_map_value_arg487), .map_value_arg488(_meirotest_map_value_arg488), .map_value_arg489(_meirotest_map_value_arg489), .map_value_arg490(_meirotest_map_value_arg490), .map_value_arg491(_meirotest_map_value_arg491), .map_value_arg492(_meirotest_map_value_arg492), .map_value_arg493(_meirotest_map_value_arg493), .map_value_arg494(_meirotest_map_value_arg494), .map_value_arg495(_meirotest_map_value_arg495), .map_value_arg496(_meirotest_map_value_arg496), .map_value_arg497(_meirotest_map_value_arg497), .map_value_arg498(_meirotest_map_value_arg498), .map_value_arg499(_meirotest_map_value_arg499), .map_value_arg500(_meirotest_map_value_arg500), .map_value_arg501(_meirotest_map_value_arg501), .map_value_arg502(_meirotest_map_value_arg502), .map_value_arg503(_meirotest_map_value_arg503), .map_value_arg504(_meirotest_map_value_arg504), .map_value_arg505(_meirotest_map_value_arg505), .map_value_arg506(_meirotest_map_value_arg506), .map_value_arg507(_meirotest_map_value_arg507), .map_value_arg508(_meirotest_map_value_arg508), .map_value_arg509(_meirotest_map_value_arg509), .map_value_arg510(_meirotest_map_value_arg510), .map_value_arg511(_meirotest_map_value_arg511));
mul_bit mul_bit_x (.m_clock(m_clock), .p_reset( p_reset), .mul_bit_exe(_mul_bit_x_mul_bit_exe), .mul_bit_result(_mul_bit_x_mul_bit_result), .mul_bit1(_mul_bit_x_mul_bit1), .mul_bit2(_mul_bit_x_mul_bit2));
mul_bit mul_bit_x_1 (.m_clock(m_clock), .p_reset( p_reset), .mul_bit_exe(_mul_bit_x_1_mul_bit_exe), .mul_bit_result(_mul_bit_x_1_mul_bit_result), .mul_bit1(_mul_bit_x_1_mul_bit1), .mul_bit2(_mul_bit_x_1_mul_bit2));

   assign  fpga_512_start = _net_2;
   assign  out_put = 1'b0;
   assign  _mul_bit_x_mul_bit_exe = 1'b0;
   assign  _mul_bit_x_p_reset = p_reset;
   assign  _mul_bit_x_m_clock = m_clock;
   assign  _mul_bit_x_1_mul_bit_exe = 1'b0;
   assign  _mul_bit_x_1_p_reset = p_reset;
   assign  _mul_bit_x_1_m_clock = m_clock;
   assign  _meirotest_map_value_arg0 = ((_net_516)?(map_test[9'b000000000]):10'b0);
   assign  _meirotest_map_value_arg1 = ((_net_515)?(map_test[9'b000000001]):10'b0);
   assign  _meirotest_map_value_arg2 = ((_net_514)?(map_test[9'b000000010]):10'b0);
   assign  _meirotest_map_value_arg3 = ((_net_513)?(map_test[9'b000000011]):10'b0);
   assign  _meirotest_map_value_arg4 = ((_net_512)?(map_test[9'b000000100]):10'b0);
   assign  _meirotest_map_value_arg5 = ((_net_511)?(map_test[9'b000000101]):10'b0);
   assign  _meirotest_map_value_arg6 = ((_net_510)?(map_test[9'b000000110]):10'b0);
   assign  _meirotest_map_value_arg7 = ((_net_509)?(map_test[9'b000000111]):10'b0);
   assign  _meirotest_map_value_arg8 = ((_net_508)?(map_test[9'b000001000]):10'b0);
   assign  _meirotest_map_value_arg9 = ((_net_507)?(map_test[9'b000001001]):10'b0);
   assign  _meirotest_map_value_arg10 = ((_net_506)?(map_test[9'b000001010]):10'b0);
   assign  _meirotest_map_value_arg11 = ((_net_505)?(map_test[9'b000001011]):10'b0);
   assign  _meirotest_map_value_arg12 = ((_net_504)?(map_test[9'b000001100]):10'b0);
   assign  _meirotest_map_value_arg13 = ((_net_503)?(map_test[9'b000001101]):10'b0);
   assign  _meirotest_map_value_arg14 = ((_net_502)?(map_test[9'b000001110]):10'b0);
   assign  _meirotest_map_value_arg15 = ((_net_501)?(map_test[9'b000001111]):10'b0);
   assign  _meirotest_map_value_arg16 = ((_net_500)?(map_test[9'b000010000]):10'b0);
   assign  _meirotest_map_value_arg17 = ((_net_499)?(map_test[9'b000010001]):10'b0);
   assign  _meirotest_map_value_arg18 = ((_net_498)?(map_test[9'b000010010]):10'b0);
   assign  _meirotest_map_value_arg19 = ((_net_497)?(map_test[9'b000010011]):10'b0);
   assign  _meirotest_map_value_arg20 = ((_net_496)?(map_test[9'b000010100]):10'b0);
   assign  _meirotest_map_value_arg21 = ((_net_495)?(map_test[9'b000010101]):10'b0);
   assign  _meirotest_map_value_arg22 = ((_net_494)?(map_test[9'b000010110]):10'b0);
   assign  _meirotest_map_value_arg23 = ((_net_493)?(map_test[9'b000010111]):10'b0);
   assign  _meirotest_map_value_arg24 = ((_net_492)?(map_test[9'b000011000]):10'b0);
   assign  _meirotest_map_value_arg25 = ((_net_491)?(map_test[9'b000011001]):10'b0);
   assign  _meirotest_map_value_arg26 = ((_net_490)?(map_test[9'b000011010]):10'b0);
   assign  _meirotest_map_value_arg27 = ((_net_489)?(map_test[9'b000011011]):10'b0);
   assign  _meirotest_map_value_arg28 = ((_net_488)?(map_test[9'b000011100]):10'b0);
   assign  _meirotest_map_value_arg29 = ((_net_487)?(map_test[9'b000011101]):10'b0);
   assign  _meirotest_map_value_arg30 = ((_net_486)?(map_test[9'b000011110]):10'b0);
   assign  _meirotest_map_value_arg31 = ((_net_485)?(map_test[9'b000011111]):10'b0);
   assign  _meirotest_map_value_arg32 = ((_net_484)?(map_test[9'b000100000]):10'b0);
   assign  _meirotest_map_value_arg33 = ((_net_483)?(map_test[9'b000100001]):10'b0);
   assign  _meirotest_map_value_arg34 = ((_net_482)?(map_test[9'b000100010]):10'b0);
   assign  _meirotest_map_value_arg35 = ((_net_481)?(map_test[9'b000100011]):10'b0);
   assign  _meirotest_map_value_arg36 = ((_net_480)?(map_test[9'b000100100]):10'b0);
   assign  _meirotest_map_value_arg37 = ((_net_479)?(map_test[9'b000100101]):10'b0);
   assign  _meirotest_map_value_arg38 = ((_net_478)?(map_test[9'b000100110]):10'b0);
   assign  _meirotest_map_value_arg39 = ((_net_477)?(map_test[9'b000100111]):10'b0);
   assign  _meirotest_map_value_arg40 = ((_net_476)?(map_test[9'b000101000]):10'b0);
   assign  _meirotest_map_value_arg41 = ((_net_475)?(map_test[9'b000101001]):10'b0);
   assign  _meirotest_map_value_arg42 = ((_net_474)?(map_test[9'b000101010]):10'b0);
   assign  _meirotest_map_value_arg43 = ((_net_473)?(map_test[9'b000101011]):10'b0);
   assign  _meirotest_map_value_arg44 = ((_net_472)?(map_test[9'b000101100]):10'b0);
   assign  _meirotest_map_value_arg45 = ((_net_471)?(map_test[9'b000101101]):10'b0);
   assign  _meirotest_map_value_arg46 = ((_net_470)?(map_test[9'b000101110]):10'b0);
   assign  _meirotest_map_value_arg47 = ((_net_469)?(map_test[9'b000101111]):10'b0);
   assign  _meirotest_map_value_arg48 = ((_net_468)?(map_test[9'b000110000]):10'b0);
   assign  _meirotest_map_value_arg49 = ((_net_467)?(map_test[9'b000110001]):10'b0);
   assign  _meirotest_map_value_arg50 = ((_net_466)?(map_test[9'b000110010]):10'b0);
   assign  _meirotest_map_value_arg51 = ((_net_465)?(map_test[9'b000110011]):10'b0);
   assign  _meirotest_map_value_arg52 = ((_net_464)?(map_test[9'b000110100]):10'b0);
   assign  _meirotest_map_value_arg53 = ((_net_463)?(map_test[9'b000110101]):10'b0);
   assign  _meirotest_map_value_arg54 = ((_net_462)?(map_test[9'b000110110]):10'b0);
   assign  _meirotest_map_value_arg55 = ((_net_461)?(map_test[9'b000110111]):10'b0);
   assign  _meirotest_map_value_arg56 = ((_net_460)?(map_test[9'b000111000]):10'b0);
   assign  _meirotest_map_value_arg57 = ((_net_459)?(map_test[9'b000111001]):10'b0);
   assign  _meirotest_map_value_arg58 = ((_net_458)?(map_test[9'b000111010]):10'b0);
   assign  _meirotest_map_value_arg59 = ((_net_457)?(map_test[9'b000111011]):10'b0);
   assign  _meirotest_map_value_arg60 = ((_net_456)?(map_test[9'b000111100]):10'b0);
   assign  _meirotest_map_value_arg61 = ((_net_455)?(map_test[9'b000111101]):10'b0);
   assign  _meirotest_map_value_arg62 = ((_net_454)?(map_test[9'b000111110]):10'b0);
   assign  _meirotest_map_value_arg63 = ((_net_453)?(map_test[9'b000111111]):10'b0);
   assign  _meirotest_map_value_arg64 = ((_net_452)?(map_test[9'b001000000]):10'b0);
   assign  _meirotest_map_value_arg65 = ((_net_451)?(map_test[9'b001000001]):10'b0);
   assign  _meirotest_map_value_arg66 = ((_net_450)?(map_test[9'b001000010]):10'b0);
   assign  _meirotest_map_value_arg67 = ((_net_449)?(map_test[9'b001000011]):10'b0);
   assign  _meirotest_map_value_arg68 = ((_net_448)?(map_test[9'b001000100]):10'b0);
   assign  _meirotest_map_value_arg69 = ((_net_447)?(map_test[9'b001000101]):10'b0);
   assign  _meirotest_map_value_arg70 = ((_net_446)?(map_test[9'b001000110]):10'b0);
   assign  _meirotest_map_value_arg71 = ((_net_445)?(map_test[9'b001000111]):10'b0);
   assign  _meirotest_map_value_arg72 = ((_net_444)?(map_test[9'b001001000]):10'b0);
   assign  _meirotest_map_value_arg73 = ((_net_443)?(map_test[9'b001001001]):10'b0);
   assign  _meirotest_map_value_arg74 = ((_net_442)?(map_test[9'b001001010]):10'b0);
   assign  _meirotest_map_value_arg75 = ((_net_441)?(map_test[9'b001001011]):10'b0);
   assign  _meirotest_map_value_arg76 = ((_net_440)?(map_test[9'b001001100]):10'b0);
   assign  _meirotest_map_value_arg77 = ((_net_439)?(map_test[9'b001001101]):10'b0);
   assign  _meirotest_map_value_arg78 = ((_net_438)?(map_test[9'b001001110]):10'b0);
   assign  _meirotest_map_value_arg79 = ((_net_437)?(map_test[9'b001001111]):10'b0);
   assign  _meirotest_map_value_arg80 = ((_net_436)?(map_test[9'b001010000]):10'b0);
   assign  _meirotest_map_value_arg81 = ((_net_435)?(map_test[9'b001010001]):10'b0);
   assign  _meirotest_map_value_arg82 = ((_net_434)?(map_test[9'b001010010]):10'b0);
   assign  _meirotest_map_value_arg83 = ((_net_433)?(map_test[9'b001010011]):10'b0);
   assign  _meirotest_map_value_arg84 = ((_net_432)?(map_test[9'b001010100]):10'b0);
   assign  _meirotest_map_value_arg85 = ((_net_431)?(map_test[9'b001010101]):10'b0);
   assign  _meirotest_map_value_arg86 = ((_net_430)?(map_test[9'b001010110]):10'b0);
   assign  _meirotest_map_value_arg87 = ((_net_429)?(map_test[9'b001010111]):10'b0);
   assign  _meirotest_map_value_arg88 = ((_net_428)?(map_test[9'b001011000]):10'b0);
   assign  _meirotest_map_value_arg89 = ((_net_427)?(map_test[9'b001011001]):10'b0);
   assign  _meirotest_map_value_arg90 = ((_net_426)?(map_test[9'b001011010]):10'b0);
   assign  _meirotest_map_value_arg91 = ((_net_425)?(map_test[9'b001011011]):10'b0);
   assign  _meirotest_map_value_arg92 = ((_net_424)?(map_test[9'b001011100]):10'b0);
   assign  _meirotest_map_value_arg93 = ((_net_423)?(map_test[9'b001011101]):10'b0);
   assign  _meirotest_map_value_arg94 = ((_net_422)?(map_test[9'b001011110]):10'b0);
   assign  _meirotest_map_value_arg95 = ((_net_421)?(map_test[9'b001011111]):10'b0);
   assign  _meirotest_map_value_arg96 = ((_net_420)?(map_test[9'b001100000]):10'b0);
   assign  _meirotest_map_value_arg97 = ((_net_419)?(map_test[9'b001100001]):10'b0);
   assign  _meirotest_map_value_arg98 = ((_net_418)?(map_test[9'b001100010]):10'b0);
   assign  _meirotest_map_value_arg99 = ((_net_417)?(map_test[9'b001100011]):10'b0);
   assign  _meirotest_map_value_arg100 = ((_net_416)?(map_test[9'b001100100]):10'b0);
   assign  _meirotest_map_value_arg101 = ((_net_415)?(map_test[9'b001100101]):10'b0);
   assign  _meirotest_map_value_arg102 = ((_net_414)?(map_test[9'b001100110]):10'b0);
   assign  _meirotest_map_value_arg103 = ((_net_413)?(map_test[9'b001100111]):10'b0);
   assign  _meirotest_map_value_arg104 = ((_net_412)?(map_test[9'b001101000]):10'b0);
   assign  _meirotest_map_value_arg105 = ((_net_411)?(map_test[9'b001101001]):10'b0);
   assign  _meirotest_map_value_arg106 = ((_net_410)?(map_test[9'b001101010]):10'b0);
   assign  _meirotest_map_value_arg107 = ((_net_409)?(map_test[9'b001101011]):10'b0);
   assign  _meirotest_map_value_arg108 = ((_net_408)?(map_test[9'b001101100]):10'b0);
   assign  _meirotest_map_value_arg109 = ((_net_407)?(map_test[9'b001101101]):10'b0);
   assign  _meirotest_map_value_arg110 = ((_net_406)?(map_test[9'b001101110]):10'b0);
   assign  _meirotest_map_value_arg111 = ((_net_405)?(map_test[9'b001101111]):10'b0);
   assign  _meirotest_map_value_arg112 = ((_net_404)?(map_test[9'b001110000]):10'b0);
   assign  _meirotest_map_value_arg113 = ((_net_403)?(map_test[9'b001110001]):10'b0);
   assign  _meirotest_map_value_arg114 = ((_net_402)?(map_test[9'b001110010]):10'b0);
   assign  _meirotest_map_value_arg115 = ((_net_401)?(map_test[9'b001110011]):10'b0);
   assign  _meirotest_map_value_arg116 = ((_net_400)?(map_test[9'b001110100]):10'b0);
   assign  _meirotest_map_value_arg117 = ((_net_399)?(map_test[9'b001110101]):10'b0);
   assign  _meirotest_map_value_arg118 = ((_net_398)?(map_test[9'b001110110]):10'b0);
   assign  _meirotest_map_value_arg119 = ((_net_397)?(map_test[9'b001110111]):10'b0);
   assign  _meirotest_map_value_arg120 = ((_net_396)?(map_test[9'b001111000]):10'b0);
   assign  _meirotest_map_value_arg121 = ((_net_395)?(map_test[9'b001111001]):10'b0);
   assign  _meirotest_map_value_arg122 = ((_net_394)?(map_test[9'b001111010]):10'b0);
   assign  _meirotest_map_value_arg123 = ((_net_393)?(map_test[9'b001111011]):10'b0);
   assign  _meirotest_map_value_arg124 = ((_net_392)?(map_test[9'b001111100]):10'b0);
   assign  _meirotest_map_value_arg125 = ((_net_391)?(map_test[9'b001111101]):10'b0);
   assign  _meirotest_map_value_arg126 = ((_net_390)?(map_test[9'b001111110]):10'b0);
   assign  _meirotest_map_value_arg127 = ((_net_389)?(map_test[9'b001111111]):10'b0);
   assign  _meirotest_map_value_arg128 = ((_net_388)?(map_test[9'b010000000]):10'b0);
   assign  _meirotest_map_value_arg129 = ((_net_387)?(map_test[9'b010000001]):10'b0);
   assign  _meirotest_map_value_arg130 = ((_net_386)?(map_test[9'b010000010]):10'b0);
   assign  _meirotest_map_value_arg131 = ((_net_385)?(map_test[9'b010000011]):10'b0);
   assign  _meirotest_map_value_arg132 = ((_net_384)?(map_test[9'b010000100]):10'b0);
   assign  _meirotest_map_value_arg133 = ((_net_383)?(map_test[9'b010000101]):10'b0);
   assign  _meirotest_map_value_arg134 = ((_net_382)?(map_test[9'b010000110]):10'b0);
   assign  _meirotest_map_value_arg135 = ((_net_381)?(map_test[9'b010000111]):10'b0);
   assign  _meirotest_map_value_arg136 = ((_net_380)?(map_test[9'b010001000]):10'b0);
   assign  _meirotest_map_value_arg137 = ((_net_379)?(map_test[9'b010001001]):10'b0);
   assign  _meirotest_map_value_arg138 = ((_net_378)?(map_test[9'b010001010]):10'b0);
   assign  _meirotest_map_value_arg139 = ((_net_377)?(map_test[9'b010001011]):10'b0);
   assign  _meirotest_map_value_arg140 = ((_net_376)?(map_test[9'b010001100]):10'b0);
   assign  _meirotest_map_value_arg141 = ((_net_375)?(map_test[9'b010001101]):10'b0);
   assign  _meirotest_map_value_arg142 = ((_net_374)?(map_test[9'b010001110]):10'b0);
   assign  _meirotest_map_value_arg143 = ((_net_373)?(map_test[9'b010001111]):10'b0);
   assign  _meirotest_map_value_arg144 = ((_net_372)?(map_test[9'b010010000]):10'b0);
   assign  _meirotest_map_value_arg145 = ((_net_371)?(map_test[9'b010010001]):10'b0);
   assign  _meirotest_map_value_arg146 = ((_net_370)?(map_test[9'b010010010]):10'b0);
   assign  _meirotest_map_value_arg147 = ((_net_369)?(map_test[9'b010010011]):10'b0);
   assign  _meirotest_map_value_arg148 = ((_net_368)?(map_test[9'b010010100]):10'b0);
   assign  _meirotest_map_value_arg149 = ((_net_367)?(map_test[9'b010010101]):10'b0);
   assign  _meirotest_map_value_arg150 = ((_net_366)?(map_test[9'b010010110]):10'b0);
   assign  _meirotest_map_value_arg151 = ((_net_365)?(map_test[9'b010010111]):10'b0);
   assign  _meirotest_map_value_arg152 = ((_net_364)?(map_test[9'b010011000]):10'b0);
   assign  _meirotest_map_value_arg153 = ((_net_363)?(map_test[9'b010011001]):10'b0);
   assign  _meirotest_map_value_arg154 = ((_net_362)?(map_test[9'b010011010]):10'b0);
   assign  _meirotest_map_value_arg155 = ((_net_361)?(map_test[9'b010011011]):10'b0);
   assign  _meirotest_map_value_arg156 = ((_net_360)?(map_test[9'b010011100]):10'b0);
   assign  _meirotest_map_value_arg157 = ((_net_359)?(map_test[9'b010011101]):10'b0);
   assign  _meirotest_map_value_arg158 = ((_net_358)?(map_test[9'b010011110]):10'b0);
   assign  _meirotest_map_value_arg159 = ((_net_357)?(map_test[9'b010011111]):10'b0);
   assign  _meirotest_map_value_arg160 = ((_net_356)?(map_test[9'b010100000]):10'b0);
   assign  _meirotest_map_value_arg161 = ((_net_355)?(map_test[9'b010100001]):10'b0);
   assign  _meirotest_map_value_arg162 = ((_net_354)?(map_test[9'b010100010]):10'b0);
   assign  _meirotest_map_value_arg163 = ((_net_353)?(map_test[9'b010100011]):10'b0);
   assign  _meirotest_map_value_arg164 = ((_net_352)?(map_test[9'b010100100]):10'b0);
   assign  _meirotest_map_value_arg165 = ((_net_351)?(map_test[9'b010100101]):10'b0);
   assign  _meirotest_map_value_arg166 = ((_net_350)?(map_test[9'b010100110]):10'b0);
   assign  _meirotest_map_value_arg167 = ((_net_349)?(map_test[9'b010100111]):10'b0);
   assign  _meirotest_map_value_arg168 = ((_net_348)?(map_test[9'b010101000]):10'b0);
   assign  _meirotest_map_value_arg169 = ((_net_347)?(map_test[9'b010101001]):10'b0);
   assign  _meirotest_map_value_arg170 = ((_net_346)?(map_test[9'b010101010]):10'b0);
   assign  _meirotest_map_value_arg171 = ((_net_345)?(map_test[9'b010101011]):10'b0);
   assign  _meirotest_map_value_arg172 = ((_net_344)?(map_test[9'b010101100]):10'b0);
   assign  _meirotest_map_value_arg173 = ((_net_343)?(map_test[9'b010101101]):10'b0);
   assign  _meirotest_map_value_arg174 = ((_net_342)?(map_test[9'b010101110]):10'b0);
   assign  _meirotest_map_value_arg175 = ((_net_341)?(map_test[9'b010101111]):10'b0);
   assign  _meirotest_map_value_arg176 = ((_net_340)?(map_test[9'b010110000]):10'b0);
   assign  _meirotest_map_value_arg177 = ((_net_339)?(map_test[9'b010110001]):10'b0);
   assign  _meirotest_map_value_arg178 = ((_net_338)?(map_test[9'b010110010]):10'b0);
   assign  _meirotest_map_value_arg179 = ((_net_337)?(map_test[9'b010110011]):10'b0);
   assign  _meirotest_map_value_arg180 = ((_net_336)?(map_test[9'b010110100]):10'b0);
   assign  _meirotest_map_value_arg181 = ((_net_335)?(map_test[9'b010110101]):10'b0);
   assign  _meirotest_map_value_arg182 = ((_net_334)?(map_test[9'b010110110]):10'b0);
   assign  _meirotest_map_value_arg183 = ((_net_333)?(map_test[9'b010110111]):10'b0);
   assign  _meirotest_map_value_arg184 = ((_net_332)?(map_test[9'b010111000]):10'b0);
   assign  _meirotest_map_value_arg185 = ((_net_331)?(map_test[9'b010111001]):10'b0);
   assign  _meirotest_map_value_arg186 = ((_net_330)?(map_test[9'b010111010]):10'b0);
   assign  _meirotest_map_value_arg187 = ((_net_329)?(map_test[9'b010111011]):10'b0);
   assign  _meirotest_map_value_arg188 = ((_net_328)?(map_test[9'b010111100]):10'b0);
   assign  _meirotest_map_value_arg189 = ((_net_327)?(map_test[9'b010111101]):10'b0);
   assign  _meirotest_map_value_arg190 = ((_net_326)?(map_test[9'b010111110]):10'b0);
   assign  _meirotest_map_value_arg191 = ((_net_325)?(map_test[9'b010111111]):10'b0);
   assign  _meirotest_map_value_arg192 = ((_net_324)?(map_test[9'b011000000]):10'b0);
   assign  _meirotest_map_value_arg193 = ((_net_323)?(map_test[9'b011000001]):10'b0);
   assign  _meirotest_map_value_arg194 = ((_net_322)?(map_test[9'b011000010]):10'b0);
   assign  _meirotest_map_value_arg195 = ((_net_321)?(map_test[9'b011000011]):10'b0);
   assign  _meirotest_map_value_arg196 = ((_net_320)?(map_test[9'b011000100]):10'b0);
   assign  _meirotest_map_value_arg197 = ((_net_319)?(map_test[9'b011000101]):10'b0);
   assign  _meirotest_map_value_arg198 = ((_net_318)?(map_test[9'b011000110]):10'b0);
   assign  _meirotest_map_value_arg199 = ((_net_317)?(map_test[9'b011000111]):10'b0);
   assign  _meirotest_map_value_arg200 = ((_net_316)?(map_test[9'b011001000]):10'b0);
   assign  _meirotest_map_value_arg201 = ((_net_315)?(map_test[9'b011001001]):10'b0);
   assign  _meirotest_map_value_arg202 = ((_net_314)?(map_test[9'b011001010]):10'b0);
   assign  _meirotest_map_value_arg203 = ((_net_313)?(map_test[9'b011001011]):10'b0);
   assign  _meirotest_map_value_arg204 = ((_net_312)?(map_test[9'b011001100]):10'b0);
   assign  _meirotest_map_value_arg205 = ((_net_311)?(map_test[9'b011001101]):10'b0);
   assign  _meirotest_map_value_arg206 = ((_net_310)?(map_test[9'b011001110]):10'b0);
   assign  _meirotest_map_value_arg207 = ((_net_309)?(map_test[9'b011001111]):10'b0);
   assign  _meirotest_map_value_arg208 = ((_net_308)?(map_test[9'b011010000]):10'b0);
   assign  _meirotest_map_value_arg209 = ((_net_307)?(map_test[9'b011010001]):10'b0);
   assign  _meirotest_map_value_arg210 = ((_net_306)?(map_test[9'b011010010]):10'b0);
   assign  _meirotest_map_value_arg211 = ((_net_305)?(map_test[9'b011010011]):10'b0);
   assign  _meirotest_map_value_arg212 = ((_net_304)?(map_test[9'b011010100]):10'b0);
   assign  _meirotest_map_value_arg213 = ((_net_303)?(map_test[9'b011010101]):10'b0);
   assign  _meirotest_map_value_arg214 = ((_net_302)?(map_test[9'b011010110]):10'b0);
   assign  _meirotest_map_value_arg215 = ((_net_301)?(map_test[9'b011010111]):10'b0);
   assign  _meirotest_map_value_arg216 = ((_net_300)?(map_test[9'b011011000]):10'b0);
   assign  _meirotest_map_value_arg217 = ((_net_299)?(map_test[9'b011011001]):10'b0);
   assign  _meirotest_map_value_arg218 = ((_net_298)?(map_test[9'b011011010]):10'b0);
   assign  _meirotest_map_value_arg219 = ((_net_297)?(map_test[9'b011011011]):10'b0);
   assign  _meirotest_map_value_arg220 = ((_net_296)?(map_test[9'b011011100]):10'b0);
   assign  _meirotest_map_value_arg221 = ((_net_295)?(map_test[9'b011011101]):10'b0);
   assign  _meirotest_map_value_arg222 = ((_net_294)?(map_test[9'b011011110]):10'b0);
   assign  _meirotest_map_value_arg223 = ((_net_293)?(map_test[9'b011011111]):10'b0);
   assign  _meirotest_map_value_arg224 = ((_net_292)?(map_test[9'b011100000]):10'b0);
   assign  _meirotest_map_value_arg225 = ((_net_291)?(map_test[9'b011100001]):10'b0);
   assign  _meirotest_map_value_arg226 = ((_net_290)?(map_test[9'b011100010]):10'b0);
   assign  _meirotest_map_value_arg227 = ((_net_289)?(map_test[9'b011100011]):10'b0);
   assign  _meirotest_map_value_arg228 = ((_net_288)?(map_test[9'b011100100]):10'b0);
   assign  _meirotest_map_value_arg229 = ((_net_287)?(map_test[9'b011100101]):10'b0);
   assign  _meirotest_map_value_arg230 = ((_net_286)?(map_test[9'b011100110]):10'b0);
   assign  _meirotest_map_value_arg231 = ((_net_285)?(map_test[9'b011100111]):10'b0);
   assign  _meirotest_map_value_arg232 = ((_net_284)?(map_test[9'b011101000]):10'b0);
   assign  _meirotest_map_value_arg233 = ((_net_283)?(map_test[9'b011101001]):10'b0);
   assign  _meirotest_map_value_arg234 = ((_net_282)?(map_test[9'b011101010]):10'b0);
   assign  _meirotest_map_value_arg235 = ((_net_281)?(map_test[9'b011101011]):10'b0);
   assign  _meirotest_map_value_arg236 = ((_net_280)?(map_test[9'b011101100]):10'b0);
   assign  _meirotest_map_value_arg237 = ((_net_279)?(map_test[9'b011101101]):10'b0);
   assign  _meirotest_map_value_arg238 = ((_net_278)?(map_test[9'b011101110]):10'b0);
   assign  _meirotest_map_value_arg239 = ((_net_277)?(map_test[9'b011101111]):10'b0);
   assign  _meirotest_map_value_arg240 = ((_net_276)?(map_test[9'b011110000]):10'b0);
   assign  _meirotest_map_value_arg241 = ((_net_275)?(map_test[9'b011110001]):10'b0);
   assign  _meirotest_map_value_arg242 = ((_net_274)?(map_test[9'b011110010]):10'b0);
   assign  _meirotest_map_value_arg243 = ((_net_273)?(map_test[9'b011110011]):10'b0);
   assign  _meirotest_map_value_arg244 = ((_net_272)?(map_test[9'b011110100]):10'b0);
   assign  _meirotest_map_value_arg245 = ((_net_271)?(map_test[9'b011110101]):10'b0);
   assign  _meirotest_map_value_arg246 = ((_net_270)?(map_test[9'b011110110]):10'b0);
   assign  _meirotest_map_value_arg247 = ((_net_269)?(map_test[9'b011110111]):10'b0);
   assign  _meirotest_map_value_arg248 = ((_net_268)?(map_test[9'b011111000]):10'b0);
   assign  _meirotest_map_value_arg249 = ((_net_267)?(map_test[9'b011111001]):10'b0);
   assign  _meirotest_map_value_arg250 = ((_net_266)?(map_test[9'b011111010]):10'b0);
   assign  _meirotest_map_value_arg251 = ((_net_265)?(map_test[9'b011111011]):10'b0);
   assign  _meirotest_map_value_arg252 = ((_net_264)?(map_test[9'b011111100]):10'b0);
   assign  _meirotest_map_value_arg253 = ((_net_263)?(map_test[9'b011111101]):10'b0);
   assign  _meirotest_map_value_arg254 = ((_net_262)?(map_test[9'b011111110]):10'b0);
   assign  _meirotest_map_value_arg255 = ((_net_261)?(map_test[9'b011111111]):10'b0);
   assign  _meirotest_map_value_arg256 = ((_net_260)?(map_test[9'b100000000]):10'b0);
   assign  _meirotest_map_value_arg257 = ((_net_259)?(map_test[9'b100000001]):10'b0);
   assign  _meirotest_map_value_arg258 = ((_net_258)?(map_test[9'b100000010]):10'b0);
   assign  _meirotest_map_value_arg259 = ((_net_257)?(map_test[9'b100000011]):10'b0);
   assign  _meirotest_map_value_arg260 = ((_net_256)?(map_test[9'b100000100]):10'b0);
   assign  _meirotest_map_value_arg261 = ((_net_255)?(map_test[9'b100000101]):10'b0);
   assign  _meirotest_map_value_arg262 = ((_net_254)?(map_test[9'b100000110]):10'b0);
   assign  _meirotest_map_value_arg263 = ((_net_253)?(map_test[9'b100000111]):10'b0);
   assign  _meirotest_map_value_arg264 = ((_net_252)?(map_test[9'b100001000]):10'b0);
   assign  _meirotest_map_value_arg265 = ((_net_251)?(map_test[9'b100001001]):10'b0);
   assign  _meirotest_map_value_arg266 = ((_net_250)?(map_test[9'b100001010]):10'b0);
   assign  _meirotest_map_value_arg267 = ((_net_249)?(map_test[9'b100001011]):10'b0);
   assign  _meirotest_map_value_arg268 = ((_net_248)?(map_test[9'b100001100]):10'b0);
   assign  _meirotest_map_value_arg269 = ((_net_247)?(map_test[9'b100001101]):10'b0);
   assign  _meirotest_map_value_arg270 = ((_net_246)?(map_test[9'b100001110]):10'b0);
   assign  _meirotest_map_value_arg271 = ((_net_245)?(map_test[9'b100001111]):10'b0);
   assign  _meirotest_map_value_arg272 = ((_net_244)?(map_test[9'b100010000]):10'b0);
   assign  _meirotest_map_value_arg273 = ((_net_243)?(map_test[9'b100010001]):10'b0);
   assign  _meirotest_map_value_arg274 = ((_net_242)?(map_test[9'b100010010]):10'b0);
   assign  _meirotest_map_value_arg275 = ((_net_241)?(map_test[9'b100010011]):10'b0);
   assign  _meirotest_map_value_arg276 = ((_net_240)?(map_test[9'b100010100]):10'b0);
   assign  _meirotest_map_value_arg277 = ((_net_239)?(map_test[9'b100010101]):10'b0);
   assign  _meirotest_map_value_arg278 = ((_net_238)?(map_test[9'b100010110]):10'b0);
   assign  _meirotest_map_value_arg279 = ((_net_237)?(map_test[9'b100010111]):10'b0);
   assign  _meirotest_map_value_arg280 = ((_net_236)?(map_test[9'b100011000]):10'b0);
   assign  _meirotest_map_value_arg281 = ((_net_235)?(map_test[9'b100011001]):10'b0);
   assign  _meirotest_map_value_arg282 = ((_net_234)?(map_test[9'b100011010]):10'b0);
   assign  _meirotest_map_value_arg283 = ((_net_233)?(map_test[9'b100011011]):10'b0);
   assign  _meirotest_map_value_arg284 = ((_net_232)?(map_test[9'b100011100]):10'b0);
   assign  _meirotest_map_value_arg285 = ((_net_231)?(map_test[9'b100011101]):10'b0);
   assign  _meirotest_map_value_arg286 = ((_net_230)?(map_test[9'b100011110]):10'b0);
   assign  _meirotest_map_value_arg287 = ((_net_229)?(map_test[9'b100011111]):10'b0);
   assign  _meirotest_map_value_arg288 = ((_net_228)?(map_test[9'b100100000]):10'b0);
   assign  _meirotest_map_value_arg289 = ((_net_227)?(map_test[9'b100100001]):10'b0);
   assign  _meirotest_map_value_arg290 = ((_net_226)?(map_test[9'b100100010]):10'b0);
   assign  _meirotest_map_value_arg291 = ((_net_225)?(map_test[9'b100100011]):10'b0);
   assign  _meirotest_map_value_arg292 = ((_net_224)?(map_test[9'b100100100]):10'b0);
   assign  _meirotest_map_value_arg293 = ((_net_223)?(map_test[9'b100100101]):10'b0);
   assign  _meirotest_map_value_arg294 = ((_net_222)?(map_test[9'b100100110]):10'b0);
   assign  _meirotest_map_value_arg295 = ((_net_221)?(map_test[9'b100100111]):10'b0);
   assign  _meirotest_map_value_arg296 = ((_net_220)?(map_test[9'b100101000]):10'b0);
   assign  _meirotest_map_value_arg297 = ((_net_219)?(map_test[9'b100101001]):10'b0);
   assign  _meirotest_map_value_arg298 = ((_net_218)?(map_test[9'b100101010]):10'b0);
   assign  _meirotest_map_value_arg299 = ((_net_217)?(map_test[9'b100101011]):10'b0);
   assign  _meirotest_map_value_arg300 = ((_net_216)?(map_test[9'b100101100]):10'b0);
   assign  _meirotest_map_value_arg301 = ((_net_215)?(map_test[9'b100101101]):10'b0);
   assign  _meirotest_map_value_arg302 = ((_net_214)?(map_test[9'b100101110]):10'b0);
   assign  _meirotest_map_value_arg303 = ((_net_213)?(map_test[9'b100101111]):10'b0);
   assign  _meirotest_map_value_arg304 = ((_net_212)?(map_test[9'b100110000]):10'b0);
   assign  _meirotest_map_value_arg305 = ((_net_211)?(map_test[9'b100110001]):10'b0);
   assign  _meirotest_map_value_arg306 = ((_net_210)?(map_test[9'b100110010]):10'b0);
   assign  _meirotest_map_value_arg307 = ((_net_209)?(map_test[9'b100110011]):10'b0);
   assign  _meirotest_map_value_arg308 = ((_net_208)?(map_test[9'b100110100]):10'b0);
   assign  _meirotest_map_value_arg309 = ((_net_207)?(map_test[9'b100110101]):10'b0);
   assign  _meirotest_map_value_arg310 = ((_net_206)?(map_test[9'b100110110]):10'b0);
   assign  _meirotest_map_value_arg311 = ((_net_205)?(map_test[9'b100110111]):10'b0);
   assign  _meirotest_map_value_arg312 = ((_net_204)?(map_test[9'b100111000]):10'b0);
   assign  _meirotest_map_value_arg313 = ((_net_203)?(map_test[9'b100111001]):10'b0);
   assign  _meirotest_map_value_arg314 = ((_net_202)?(map_test[9'b100111010]):10'b0);
   assign  _meirotest_map_value_arg315 = ((_net_201)?(map_test[9'b100111011]):10'b0);
   assign  _meirotest_map_value_arg316 = ((_net_200)?(map_test[9'b100111100]):10'b0);
   assign  _meirotest_map_value_arg317 = ((_net_199)?(map_test[9'b100111101]):10'b0);
   assign  _meirotest_map_value_arg318 = ((_net_198)?(map_test[9'b100111110]):10'b0);
   assign  _meirotest_map_value_arg319 = ((_net_197)?(map_test[9'b100111111]):10'b0);
   assign  _meirotest_map_value_arg320 = ((_net_196)?(map_test[9'b101000000]):10'b0);
   assign  _meirotest_map_value_arg321 = ((_net_195)?(map_test[9'b101000001]):10'b0);
   assign  _meirotest_map_value_arg322 = ((_net_194)?(map_test[9'b101000010]):10'b0);
   assign  _meirotest_map_value_arg323 = ((_net_193)?(map_test[9'b101000011]):10'b0);
   assign  _meirotest_map_value_arg324 = ((_net_192)?(map_test[9'b101000100]):10'b0);
   assign  _meirotest_map_value_arg325 = ((_net_191)?(map_test[9'b101000101]):10'b0);
   assign  _meirotest_map_value_arg326 = ((_net_190)?(map_test[9'b101000110]):10'b0);
   assign  _meirotest_map_value_arg327 = ((_net_189)?(map_test[9'b101000111]):10'b0);
   assign  _meirotest_map_value_arg328 = ((_net_188)?(map_test[9'b101001000]):10'b0);
   assign  _meirotest_map_value_arg329 = ((_net_187)?(map_test[9'b101001001]):10'b0);
   assign  _meirotest_map_value_arg330 = ((_net_186)?(map_test[9'b101001010]):10'b0);
   assign  _meirotest_map_value_arg331 = ((_net_185)?(map_test[9'b101001011]):10'b0);
   assign  _meirotest_map_value_arg332 = ((_net_184)?(map_test[9'b101001100]):10'b0);
   assign  _meirotest_map_value_arg333 = ((_net_183)?(map_test[9'b101001101]):10'b0);
   assign  _meirotest_map_value_arg334 = ((_net_182)?(map_test[9'b101001110]):10'b0);
   assign  _meirotest_map_value_arg335 = ((_net_181)?(map_test[9'b101001111]):10'b0);
   assign  _meirotest_map_value_arg336 = ((_net_180)?(map_test[9'b101010000]):10'b0);
   assign  _meirotest_map_value_arg337 = ((_net_179)?(map_test[9'b101010001]):10'b0);
   assign  _meirotest_map_value_arg338 = ((_net_178)?(map_test[9'b101010010]):10'b0);
   assign  _meirotest_map_value_arg339 = ((_net_177)?(map_test[9'b101010011]):10'b0);
   assign  _meirotest_map_value_arg340 = ((_net_176)?(map_test[9'b101010100]):10'b0);
   assign  _meirotest_map_value_arg341 = ((_net_175)?(map_test[9'b101010101]):10'b0);
   assign  _meirotest_map_value_arg342 = ((_net_174)?(map_test[9'b101010110]):10'b0);
   assign  _meirotest_map_value_arg343 = ((_net_173)?(map_test[9'b101010111]):10'b0);
   assign  _meirotest_map_value_arg344 = ((_net_172)?(map_test[9'b101011000]):10'b0);
   assign  _meirotest_map_value_arg345 = ((_net_171)?(map_test[9'b101011001]):10'b0);
   assign  _meirotest_map_value_arg346 = ((_net_170)?(map_test[9'b101011010]):10'b0);
   assign  _meirotest_map_value_arg347 = ((_net_169)?(map_test[9'b101011011]):10'b0);
   assign  _meirotest_map_value_arg348 = ((_net_168)?(map_test[9'b101011100]):10'b0);
   assign  _meirotest_map_value_arg349 = ((_net_167)?(map_test[9'b101011101]):10'b0);
   assign  _meirotest_map_value_arg350 = ((_net_166)?(map_test[9'b101011110]):10'b0);
   assign  _meirotest_map_value_arg351 = ((_net_165)?(map_test[9'b101011111]):10'b0);
   assign  _meirotest_map_value_arg352 = ((_net_164)?(map_test[9'b101100000]):10'b0);
   assign  _meirotest_map_value_arg353 = ((_net_163)?(map_test[9'b101100001]):10'b0);
   assign  _meirotest_map_value_arg354 = ((_net_162)?(map_test[9'b101100010]):10'b0);
   assign  _meirotest_map_value_arg355 = ((_net_161)?(map_test[9'b101100011]):10'b0);
   assign  _meirotest_map_value_arg356 = ((_net_160)?(map_test[9'b101100100]):10'b0);
   assign  _meirotest_map_value_arg357 = ((_net_159)?(map_test[9'b101100101]):10'b0);
   assign  _meirotest_map_value_arg358 = ((_net_158)?(map_test[9'b101100110]):10'b0);
   assign  _meirotest_map_value_arg359 = ((_net_157)?(map_test[9'b101100111]):10'b0);
   assign  _meirotest_map_value_arg360 = ((_net_156)?(map_test[9'b101101000]):10'b0);
   assign  _meirotest_map_value_arg361 = ((_net_155)?(map_test[9'b101101001]):10'b0);
   assign  _meirotest_map_value_arg362 = ((_net_154)?(map_test[9'b101101010]):10'b0);
   assign  _meirotest_map_value_arg363 = ((_net_153)?(map_test[9'b101101011]):10'b0);
   assign  _meirotest_map_value_arg364 = ((_net_152)?(map_test[9'b101101100]):10'b0);
   assign  _meirotest_map_value_arg365 = ((_net_151)?(map_test[9'b101101101]):10'b0);
   assign  _meirotest_map_value_arg366 = ((_net_150)?(map_test[9'b101101110]):10'b0);
   assign  _meirotest_map_value_arg367 = ((_net_149)?(map_test[9'b101101111]):10'b0);
   assign  _meirotest_map_value_arg368 = ((_net_148)?(map_test[9'b101110000]):10'b0);
   assign  _meirotest_map_value_arg369 = ((_net_147)?(map_test[9'b101110001]):10'b0);
   assign  _meirotest_map_value_arg370 = ((_net_146)?(map_test[9'b101110010]):10'b0);
   assign  _meirotest_map_value_arg371 = ((_net_145)?(map_test[9'b101110011]):10'b0);
   assign  _meirotest_map_value_arg372 = ((_net_144)?(map_test[9'b101110100]):10'b0);
   assign  _meirotest_map_value_arg373 = ((_net_143)?(map_test[9'b101110101]):10'b0);
   assign  _meirotest_map_value_arg374 = ((_net_142)?(map_test[9'b101110110]):10'b0);
   assign  _meirotest_map_value_arg375 = ((_net_141)?(map_test[9'b101110111]):10'b0);
   assign  _meirotest_map_value_arg376 = ((_net_140)?(map_test[9'b101111000]):10'b0);
   assign  _meirotest_map_value_arg377 = ((_net_139)?(map_test[9'b101111001]):10'b0);
   assign  _meirotest_map_value_arg378 = ((_net_138)?(map_test[9'b101111010]):10'b0);
   assign  _meirotest_map_value_arg379 = ((_net_137)?(map_test[9'b101111011]):10'b0);
   assign  _meirotest_map_value_arg380 = ((_net_136)?(map_test[9'b101111100]):10'b0);
   assign  _meirotest_map_value_arg381 = ((_net_135)?(map_test[9'b101111101]):10'b0);
   assign  _meirotest_map_value_arg382 = ((_net_134)?(map_test[9'b101111110]):10'b0);
   assign  _meirotest_map_value_arg383 = ((_net_133)?(map_test[9'b101111111]):10'b0);
   assign  _meirotest_map_value_arg384 = ((_net_132)?(map_test[9'b110000000]):10'b0);
   assign  _meirotest_map_value_arg385 = ((_net_131)?(map_test[9'b110000001]):10'b0);
   assign  _meirotest_map_value_arg386 = ((_net_130)?(map_test[9'b110000010]):10'b0);
   assign  _meirotest_map_value_arg387 = ((_net_129)?(map_test[9'b110000011]):10'b0);
   assign  _meirotest_map_value_arg388 = ((_net_128)?(map_test[9'b110000100]):10'b0);
   assign  _meirotest_map_value_arg389 = ((_net_127)?(map_test[9'b110000101]):10'b0);
   assign  _meirotest_map_value_arg390 = ((_net_126)?(map_test[9'b110000110]):10'b0);
   assign  _meirotest_map_value_arg391 = ((_net_125)?(map_test[9'b110000111]):10'b0);
   assign  _meirotest_map_value_arg392 = ((_net_124)?(map_test[9'b110001000]):10'b0);
   assign  _meirotest_map_value_arg393 = ((_net_123)?(map_test[9'b110001001]):10'b0);
   assign  _meirotest_map_value_arg394 = ((_net_122)?(map_test[9'b110001010]):10'b0);
   assign  _meirotest_map_value_arg395 = ((_net_121)?(map_test[9'b110001011]):10'b0);
   assign  _meirotest_map_value_arg396 = ((_net_120)?(map_test[9'b110001100]):10'b0);
   assign  _meirotest_map_value_arg397 = ((_net_119)?(map_test[9'b110001101]):10'b0);
   assign  _meirotest_map_value_arg398 = ((_net_118)?(map_test[9'b110001110]):10'b0);
   assign  _meirotest_map_value_arg399 = ((_net_117)?(map_test[9'b110001111]):10'b0);
   assign  _meirotest_map_value_arg400 = ((_net_116)?(map_test[9'b110010000]):10'b0);
   assign  _meirotest_map_value_arg401 = ((_net_115)?(map_test[9'b110010001]):10'b0);
   assign  _meirotest_map_value_arg402 = ((_net_114)?(map_test[9'b110010010]):10'b0);
   assign  _meirotest_map_value_arg403 = ((_net_113)?(map_test[9'b110010011]):10'b0);
   assign  _meirotest_map_value_arg404 = ((_net_112)?(map_test[9'b110010100]):10'b0);
   assign  _meirotest_map_value_arg405 = ((_net_111)?(map_test[9'b110010101]):10'b0);
   assign  _meirotest_map_value_arg406 = ((_net_110)?(map_test[9'b110010110]):10'b0);
   assign  _meirotest_map_value_arg407 = ((_net_109)?(map_test[9'b110010111]):10'b0);
   assign  _meirotest_map_value_arg408 = ((_net_108)?(map_test[9'b110011000]):10'b0);
   assign  _meirotest_map_value_arg409 = ((_net_107)?(map_test[9'b110011001]):10'b0);
   assign  _meirotest_map_value_arg410 = ((_net_106)?(map_test[9'b110011010]):10'b0);
   assign  _meirotest_map_value_arg411 = ((_net_105)?(map_test[9'b110011011]):10'b0);
   assign  _meirotest_map_value_arg412 = ((_net_104)?(map_test[9'b110011100]):10'b0);
   assign  _meirotest_map_value_arg413 = ((_net_103)?(map_test[9'b110011101]):10'b0);
   assign  _meirotest_map_value_arg414 = ((_net_102)?(map_test[9'b110011110]):10'b0);
   assign  _meirotest_map_value_arg415 = ((_net_101)?(map_test[9'b110011111]):10'b0);
   assign  _meirotest_map_value_arg416 = ((_net_100)?(map_test[9'b110100000]):10'b0);
   assign  _meirotest_map_value_arg417 = ((_net_99)?(map_test[9'b110100001]):10'b0);
   assign  _meirotest_map_value_arg418 = ((_net_98)?(map_test[9'b110100010]):10'b0);
   assign  _meirotest_map_value_arg419 = ((_net_97)?(map_test[9'b110100011]):10'b0);
   assign  _meirotest_map_value_arg420 = ((_net_96)?(map_test[9'b110100100]):10'b0);
   assign  _meirotest_map_value_arg421 = ((_net_95)?(map_test[9'b110100101]):10'b0);
   assign  _meirotest_map_value_arg422 = ((_net_94)?(map_test[9'b110100110]):10'b0);
   assign  _meirotest_map_value_arg423 = ((_net_93)?(map_test[9'b110100111]):10'b0);
   assign  _meirotest_map_value_arg424 = ((_net_92)?(map_test[9'b110101000]):10'b0);
   assign  _meirotest_map_value_arg425 = ((_net_91)?(map_test[9'b110101001]):10'b0);
   assign  _meirotest_map_value_arg426 = ((_net_90)?(map_test[9'b110101010]):10'b0);
   assign  _meirotest_map_value_arg427 = ((_net_89)?(map_test[9'b110101011]):10'b0);
   assign  _meirotest_map_value_arg428 = ((_net_88)?(map_test[9'b110101100]):10'b0);
   assign  _meirotest_map_value_arg429 = ((_net_87)?(map_test[9'b110101101]):10'b0);
   assign  _meirotest_map_value_arg430 = ((_net_86)?(map_test[9'b110101110]):10'b0);
   assign  _meirotest_map_value_arg431 = ((_net_85)?(map_test[9'b110101111]):10'b0);
   assign  _meirotest_map_value_arg432 = ((_net_84)?(map_test[9'b110110000]):10'b0);
   assign  _meirotest_map_value_arg433 = ((_net_83)?(map_test[9'b110110001]):10'b0);
   assign  _meirotest_map_value_arg434 = ((_net_82)?(map_test[9'b110110010]):10'b0);
   assign  _meirotest_map_value_arg435 = ((_net_81)?(map_test[9'b110110011]):10'b0);
   assign  _meirotest_map_value_arg436 = ((_net_80)?(map_test[9'b110110100]):10'b0);
   assign  _meirotest_map_value_arg437 = ((_net_79)?(map_test[9'b110110101]):10'b0);
   assign  _meirotest_map_value_arg438 = ((_net_78)?(map_test[9'b110110110]):10'b0);
   assign  _meirotest_map_value_arg439 = ((_net_77)?(map_test[9'b110110111]):10'b0);
   assign  _meirotest_map_value_arg440 = ((_net_76)?(map_test[9'b110111000]):10'b0);
   assign  _meirotest_map_value_arg441 = ((_net_75)?(map_test[9'b110111001]):10'b0);
   assign  _meirotest_map_value_arg442 = ((_net_74)?(map_test[9'b110111010]):10'b0);
   assign  _meirotest_map_value_arg443 = ((_net_73)?(map_test[9'b110111011]):10'b0);
   assign  _meirotest_map_value_arg444 = ((_net_72)?(map_test[9'b110111100]):10'b0);
   assign  _meirotest_map_value_arg445 = ((_net_71)?(map_test[9'b110111101]):10'b0);
   assign  _meirotest_map_value_arg446 = ((_net_70)?(map_test[9'b110111110]):10'b0);
   assign  _meirotest_map_value_arg447 = ((_net_69)?(map_test[9'b110111111]):10'b0);
   assign  _meirotest_map_value_arg448 = ((_net_68)?(map_test[9'b111000000]):10'b0);
   assign  _meirotest_map_value_arg449 = ((_net_67)?(map_test[9'b111000001]):10'b0);
   assign  _meirotest_map_value_arg450 = ((_net_66)?(map_test[9'b111000010]):10'b0);
   assign  _meirotest_map_value_arg451 = ((_net_65)?(map_test[9'b111000011]):10'b0);
   assign  _meirotest_map_value_arg452 = ((_net_64)?(map_test[9'b111000100]):10'b0);
   assign  _meirotest_map_value_arg453 = ((_net_63)?(map_test[9'b111000101]):10'b0);
   assign  _meirotest_map_value_arg454 = ((_net_62)?(map_test[9'b111000110]):10'b0);
   assign  _meirotest_map_value_arg455 = ((_net_61)?(map_test[9'b111000111]):10'b0);
   assign  _meirotest_map_value_arg456 = ((_net_60)?(map_test[9'b111001000]):10'b0);
   assign  _meirotest_map_value_arg457 = ((_net_59)?(map_test[9'b111001001]):10'b0);
   assign  _meirotest_map_value_arg458 = ((_net_58)?(map_test[9'b111001010]):10'b0);
   assign  _meirotest_map_value_arg459 = ((_net_57)?(map_test[9'b111001011]):10'b0);
   assign  _meirotest_map_value_arg460 = ((_net_56)?(map_test[9'b111001100]):10'b0);
   assign  _meirotest_map_value_arg461 = ((_net_55)?(map_test[9'b111001101]):10'b0);
   assign  _meirotest_map_value_arg462 = ((_net_54)?(map_test[9'b111001110]):10'b0);
   assign  _meirotest_map_value_arg463 = ((_net_53)?(map_test[9'b111001111]):10'b0);
   assign  _meirotest_map_value_arg464 = ((_net_52)?(map_test[9'b111010000]):10'b0);
   assign  _meirotest_map_value_arg465 = ((_net_51)?(map_test[9'b111010001]):10'b0);
   assign  _meirotest_map_value_arg466 = ((_net_50)?(map_test[9'b111010010]):10'b0);
   assign  _meirotest_map_value_arg467 = ((_net_49)?(map_test[9'b111010011]):10'b0);
   assign  _meirotest_map_value_arg468 = ((_net_48)?(map_test[9'b111010100]):10'b0);
   assign  _meirotest_map_value_arg469 = ((_net_47)?(map_test[9'b111010101]):10'b0);
   assign  _meirotest_map_value_arg470 = ((_net_46)?(map_test[9'b111010110]):10'b0);
   assign  _meirotest_map_value_arg471 = ((_net_45)?(map_test[9'b111010111]):10'b0);
   assign  _meirotest_map_value_arg472 = ((_net_44)?(map_test[9'b111011000]):10'b0);
   assign  _meirotest_map_value_arg473 = ((_net_43)?(map_test[9'b111011001]):10'b0);
   assign  _meirotest_map_value_arg474 = ((_net_42)?(map_test[9'b111011010]):10'b0);
   assign  _meirotest_map_value_arg475 = ((_net_41)?(map_test[9'b111011011]):10'b0);
   assign  _meirotest_map_value_arg476 = ((_net_40)?(map_test[9'b111011100]):10'b0);
   assign  _meirotest_map_value_arg477 = ((_net_39)?(map_test[9'b111011101]):10'b0);
   assign  _meirotest_map_value_arg478 = ((_net_38)?(map_test[9'b111011110]):10'b0);
   assign  _meirotest_map_value_arg479 = ((_net_37)?(map_test[9'b111011111]):10'b0);
   assign  _meirotest_map_value_arg480 = ((_net_36)?(map_test[9'b111100000]):10'b0);
   assign  _meirotest_map_value_arg481 = ((_net_35)?(map_test[9'b111100001]):10'b0);
   assign  _meirotest_map_value_arg482 = ((_net_34)?(map_test[9'b111100010]):10'b0);
   assign  _meirotest_map_value_arg483 = ((_net_33)?(map_test[9'b111100011]):10'b0);
   assign  _meirotest_map_value_arg484 = ((_net_32)?(map_test[9'b111100100]):10'b0);
   assign  _meirotest_map_value_arg485 = ((_net_31)?(map_test[9'b111100101]):10'b0);
   assign  _meirotest_map_value_arg486 = ((_net_30)?(map_test[9'b111100110]):10'b0);
   assign  _meirotest_map_value_arg487 = ((_net_29)?(map_test[9'b111100111]):10'b0);
   assign  _meirotest_map_value_arg488 = ((_net_28)?(map_test[9'b111101000]):10'b0);
   assign  _meirotest_map_value_arg489 = ((_net_27)?(map_test[9'b111101001]):10'b0);
   assign  _meirotest_map_value_arg490 = ((_net_26)?(map_test[9'b111101010]):10'b0);
   assign  _meirotest_map_value_arg491 = ((_net_25)?(map_test[9'b111101011]):10'b0);
   assign  _meirotest_map_value_arg492 = ((_net_24)?(map_test[9'b111101100]):10'b0);
   assign  _meirotest_map_value_arg493 = ((_net_23)?(map_test[9'b111101101]):10'b0);
   assign  _meirotest_map_value_arg494 = ((_net_22)?(map_test[9'b111101110]):10'b0);
   assign  _meirotest_map_value_arg495 = ((_net_21)?(map_test[9'b111101111]):10'b0);
   assign  _meirotest_map_value_arg496 = ((_net_20)?(map_test[9'b111110000]):10'b0);
   assign  _meirotest_map_value_arg497 = ((_net_19)?(map_test[9'b111110001]):10'b0);
   assign  _meirotest_map_value_arg498 = ((_net_18)?(map_test[9'b111110010]):10'b0);
   assign  _meirotest_map_value_arg499 = ((_net_17)?(map_test[9'b111110011]):10'b0);
   assign  _meirotest_map_value_arg500 = ((_net_16)?(map_test[9'b111110100]):10'b0);
   assign  _meirotest_map_value_arg501 = ((_net_15)?(map_test[9'b111110101]):10'b0);
   assign  _meirotest_map_value_arg502 = ((_net_14)?(map_test[9'b111110110]):10'b0);
   assign  _meirotest_map_value_arg503 = ((_net_13)?(map_test[9'b111110111]):10'b0);
   assign  _meirotest_map_value_arg504 = ((_net_12)?(map_test[9'b111111000]):10'b0);
   assign  _meirotest_map_value_arg505 = ((_net_11)?(map_test[9'b111111001]):10'b0);
   assign  _meirotest_map_value_arg506 = ((_net_10)?(map_test[9'b111111010]):10'b0);
   assign  _meirotest_map_value_arg507 = ((_net_9)?(map_test[9'b111111011]):10'b0);
   assign  _meirotest_map_value_arg508 = ((_net_8)?(map_test[9'b111111100]):10'b0);
   assign  _meirotest_map_value_arg509 = ((_net_7)?(map_test[9'b111111101]):10'b0);
   assign  _meirotest_map_value_arg510 = ((_net_6)?(map_test[9'b111111110]):10'b0);
   assign  _meirotest_map_value_arg511 = ((_net_5)?(map_test[9'b111111111]):10'b0);
   assign  _meirotest_in_do = _net_4;
   assign  _meirotest_p_reset = p_reset;
   assign  _meirotest_m_clock = m_clock;
   assign  _net_0 = (end_reg==2'b11);
   assign  _net_1 = (~_net_0);
   assign  _net_2 = (end_reg==2'b01);
   assign  _net_4 = (fpga_512_start|_reg_3);
   assign  _net_5 = (fpga_512_start|_reg_3);
   assign  _net_6 = (fpga_512_start|_reg_3);
   assign  _net_7 = (fpga_512_start|_reg_3);
   assign  _net_8 = (fpga_512_start|_reg_3);
   assign  _net_9 = (fpga_512_start|_reg_3);
   assign  _net_10 = (fpga_512_start|_reg_3);
   assign  _net_11 = (fpga_512_start|_reg_3);
   assign  _net_12 = (fpga_512_start|_reg_3);
   assign  _net_13 = (fpga_512_start|_reg_3);
   assign  _net_14 = (fpga_512_start|_reg_3);
   assign  _net_15 = (fpga_512_start|_reg_3);
   assign  _net_16 = (fpga_512_start|_reg_3);
   assign  _net_17 = (fpga_512_start|_reg_3);
   assign  _net_18 = (fpga_512_start|_reg_3);
   assign  _net_19 = (fpga_512_start|_reg_3);
   assign  _net_20 = (fpga_512_start|_reg_3);
   assign  _net_21 = (fpga_512_start|_reg_3);
   assign  _net_22 = (fpga_512_start|_reg_3);
   assign  _net_23 = (fpga_512_start|_reg_3);
   assign  _net_24 = (fpga_512_start|_reg_3);
   assign  _net_25 = (fpga_512_start|_reg_3);
   assign  _net_26 = (fpga_512_start|_reg_3);
   assign  _net_27 = (fpga_512_start|_reg_3);
   assign  _net_28 = (fpga_512_start|_reg_3);
   assign  _net_29 = (fpga_512_start|_reg_3);
   assign  _net_30 = (fpga_512_start|_reg_3);
   assign  _net_31 = (fpga_512_start|_reg_3);
   assign  _net_32 = (fpga_512_start|_reg_3);
   assign  _net_33 = (fpga_512_start|_reg_3);
   assign  _net_34 = (fpga_512_start|_reg_3);
   assign  _net_35 = (fpga_512_start|_reg_3);
   assign  _net_36 = (fpga_512_start|_reg_3);
   assign  _net_37 = (fpga_512_start|_reg_3);
   assign  _net_38 = (fpga_512_start|_reg_3);
   assign  _net_39 = (fpga_512_start|_reg_3);
   assign  _net_40 = (fpga_512_start|_reg_3);
   assign  _net_41 = (fpga_512_start|_reg_3);
   assign  _net_42 = (fpga_512_start|_reg_3);
   assign  _net_43 = (fpga_512_start|_reg_3);
   assign  _net_44 = (fpga_512_start|_reg_3);
   assign  _net_45 = (fpga_512_start|_reg_3);
   assign  _net_46 = (fpga_512_start|_reg_3);
   assign  _net_47 = (fpga_512_start|_reg_3);
   assign  _net_48 = (fpga_512_start|_reg_3);
   assign  _net_49 = (fpga_512_start|_reg_3);
   assign  _net_50 = (fpga_512_start|_reg_3);
   assign  _net_51 = (fpga_512_start|_reg_3);
   assign  _net_52 = (fpga_512_start|_reg_3);
   assign  _net_53 = (fpga_512_start|_reg_3);
   assign  _net_54 = (fpga_512_start|_reg_3);
   assign  _net_55 = (fpga_512_start|_reg_3);
   assign  _net_56 = (fpga_512_start|_reg_3);
   assign  _net_57 = (fpga_512_start|_reg_3);
   assign  _net_58 = (fpga_512_start|_reg_3);
   assign  _net_59 = (fpga_512_start|_reg_3);
   assign  _net_60 = (fpga_512_start|_reg_3);
   assign  _net_61 = (fpga_512_start|_reg_3);
   assign  _net_62 = (fpga_512_start|_reg_3);
   assign  _net_63 = (fpga_512_start|_reg_3);
   assign  _net_64 = (fpga_512_start|_reg_3);
   assign  _net_65 = (fpga_512_start|_reg_3);
   assign  _net_66 = (fpga_512_start|_reg_3);
   assign  _net_67 = (fpga_512_start|_reg_3);
   assign  _net_68 = (fpga_512_start|_reg_3);
   assign  _net_69 = (fpga_512_start|_reg_3);
   assign  _net_70 = (fpga_512_start|_reg_3);
   assign  _net_71 = (fpga_512_start|_reg_3);
   assign  _net_72 = (fpga_512_start|_reg_3);
   assign  _net_73 = (fpga_512_start|_reg_3);
   assign  _net_74 = (fpga_512_start|_reg_3);
   assign  _net_75 = (fpga_512_start|_reg_3);
   assign  _net_76 = (fpga_512_start|_reg_3);
   assign  _net_77 = (fpga_512_start|_reg_3);
   assign  _net_78 = (fpga_512_start|_reg_3);
   assign  _net_79 = (fpga_512_start|_reg_3);
   assign  _net_80 = (fpga_512_start|_reg_3);
   assign  _net_81 = (fpga_512_start|_reg_3);
   assign  _net_82 = (fpga_512_start|_reg_3);
   assign  _net_83 = (fpga_512_start|_reg_3);
   assign  _net_84 = (fpga_512_start|_reg_3);
   assign  _net_85 = (fpga_512_start|_reg_3);
   assign  _net_86 = (fpga_512_start|_reg_3);
   assign  _net_87 = (fpga_512_start|_reg_3);
   assign  _net_88 = (fpga_512_start|_reg_3);
   assign  _net_89 = (fpga_512_start|_reg_3);
   assign  _net_90 = (fpga_512_start|_reg_3);
   assign  _net_91 = (fpga_512_start|_reg_3);
   assign  _net_92 = (fpga_512_start|_reg_3);
   assign  _net_93 = (fpga_512_start|_reg_3);
   assign  _net_94 = (fpga_512_start|_reg_3);
   assign  _net_95 = (fpga_512_start|_reg_3);
   assign  _net_96 = (fpga_512_start|_reg_3);
   assign  _net_97 = (fpga_512_start|_reg_3);
   assign  _net_98 = (fpga_512_start|_reg_3);
   assign  _net_99 = (fpga_512_start|_reg_3);
   assign  _net_100 = (fpga_512_start|_reg_3);
   assign  _net_101 = (fpga_512_start|_reg_3);
   assign  _net_102 = (fpga_512_start|_reg_3);
   assign  _net_103 = (fpga_512_start|_reg_3);
   assign  _net_104 = (fpga_512_start|_reg_3);
   assign  _net_105 = (fpga_512_start|_reg_3);
   assign  _net_106 = (fpga_512_start|_reg_3);
   assign  _net_107 = (fpga_512_start|_reg_3);
   assign  _net_108 = (fpga_512_start|_reg_3);
   assign  _net_109 = (fpga_512_start|_reg_3);
   assign  _net_110 = (fpga_512_start|_reg_3);
   assign  _net_111 = (fpga_512_start|_reg_3);
   assign  _net_112 = (fpga_512_start|_reg_3);
   assign  _net_113 = (fpga_512_start|_reg_3);
   assign  _net_114 = (fpga_512_start|_reg_3);
   assign  _net_115 = (fpga_512_start|_reg_3);
   assign  _net_116 = (fpga_512_start|_reg_3);
   assign  _net_117 = (fpga_512_start|_reg_3);
   assign  _net_118 = (fpga_512_start|_reg_3);
   assign  _net_119 = (fpga_512_start|_reg_3);
   assign  _net_120 = (fpga_512_start|_reg_3);
   assign  _net_121 = (fpga_512_start|_reg_3);
   assign  _net_122 = (fpga_512_start|_reg_3);
   assign  _net_123 = (fpga_512_start|_reg_3);
   assign  _net_124 = (fpga_512_start|_reg_3);
   assign  _net_125 = (fpga_512_start|_reg_3);
   assign  _net_126 = (fpga_512_start|_reg_3);
   assign  _net_127 = (fpga_512_start|_reg_3);
   assign  _net_128 = (fpga_512_start|_reg_3);
   assign  _net_129 = (fpga_512_start|_reg_3);
   assign  _net_130 = (fpga_512_start|_reg_3);
   assign  _net_131 = (fpga_512_start|_reg_3);
   assign  _net_132 = (fpga_512_start|_reg_3);
   assign  _net_133 = (fpga_512_start|_reg_3);
   assign  _net_134 = (fpga_512_start|_reg_3);
   assign  _net_135 = (fpga_512_start|_reg_3);
   assign  _net_136 = (fpga_512_start|_reg_3);
   assign  _net_137 = (fpga_512_start|_reg_3);
   assign  _net_138 = (fpga_512_start|_reg_3);
   assign  _net_139 = (fpga_512_start|_reg_3);
   assign  _net_140 = (fpga_512_start|_reg_3);
   assign  _net_141 = (fpga_512_start|_reg_3);
   assign  _net_142 = (fpga_512_start|_reg_3);
   assign  _net_143 = (fpga_512_start|_reg_3);
   assign  _net_144 = (fpga_512_start|_reg_3);
   assign  _net_145 = (fpga_512_start|_reg_3);
   assign  _net_146 = (fpga_512_start|_reg_3);
   assign  _net_147 = (fpga_512_start|_reg_3);
   assign  _net_148 = (fpga_512_start|_reg_3);
   assign  _net_149 = (fpga_512_start|_reg_3);
   assign  _net_150 = (fpga_512_start|_reg_3);
   assign  _net_151 = (fpga_512_start|_reg_3);
   assign  _net_152 = (fpga_512_start|_reg_3);
   assign  _net_153 = (fpga_512_start|_reg_3);
   assign  _net_154 = (fpga_512_start|_reg_3);
   assign  _net_155 = (fpga_512_start|_reg_3);
   assign  _net_156 = (fpga_512_start|_reg_3);
   assign  _net_157 = (fpga_512_start|_reg_3);
   assign  _net_158 = (fpga_512_start|_reg_3);
   assign  _net_159 = (fpga_512_start|_reg_3);
   assign  _net_160 = (fpga_512_start|_reg_3);
   assign  _net_161 = (fpga_512_start|_reg_3);
   assign  _net_162 = (fpga_512_start|_reg_3);
   assign  _net_163 = (fpga_512_start|_reg_3);
   assign  _net_164 = (fpga_512_start|_reg_3);
   assign  _net_165 = (fpga_512_start|_reg_3);
   assign  _net_166 = (fpga_512_start|_reg_3);
   assign  _net_167 = (fpga_512_start|_reg_3);
   assign  _net_168 = (fpga_512_start|_reg_3);
   assign  _net_169 = (fpga_512_start|_reg_3);
   assign  _net_170 = (fpga_512_start|_reg_3);
   assign  _net_171 = (fpga_512_start|_reg_3);
   assign  _net_172 = (fpga_512_start|_reg_3);
   assign  _net_173 = (fpga_512_start|_reg_3);
   assign  _net_174 = (fpga_512_start|_reg_3);
   assign  _net_175 = (fpga_512_start|_reg_3);
   assign  _net_176 = (fpga_512_start|_reg_3);
   assign  _net_177 = (fpga_512_start|_reg_3);
   assign  _net_178 = (fpga_512_start|_reg_3);
   assign  _net_179 = (fpga_512_start|_reg_3);
   assign  _net_180 = (fpga_512_start|_reg_3);
   assign  _net_181 = (fpga_512_start|_reg_3);
   assign  _net_182 = (fpga_512_start|_reg_3);
   assign  _net_183 = (fpga_512_start|_reg_3);
   assign  _net_184 = (fpga_512_start|_reg_3);
   assign  _net_185 = (fpga_512_start|_reg_3);
   assign  _net_186 = (fpga_512_start|_reg_3);
   assign  _net_187 = (fpga_512_start|_reg_3);
   assign  _net_188 = (fpga_512_start|_reg_3);
   assign  _net_189 = (fpga_512_start|_reg_3);
   assign  _net_190 = (fpga_512_start|_reg_3);
   assign  _net_191 = (fpga_512_start|_reg_3);
   assign  _net_192 = (fpga_512_start|_reg_3);
   assign  _net_193 = (fpga_512_start|_reg_3);
   assign  _net_194 = (fpga_512_start|_reg_3);
   assign  _net_195 = (fpga_512_start|_reg_3);
   assign  _net_196 = (fpga_512_start|_reg_3);
   assign  _net_197 = (fpga_512_start|_reg_3);
   assign  _net_198 = (fpga_512_start|_reg_3);
   assign  _net_199 = (fpga_512_start|_reg_3);
   assign  _net_200 = (fpga_512_start|_reg_3);
   assign  _net_201 = (fpga_512_start|_reg_3);
   assign  _net_202 = (fpga_512_start|_reg_3);
   assign  _net_203 = (fpga_512_start|_reg_3);
   assign  _net_204 = (fpga_512_start|_reg_3);
   assign  _net_205 = (fpga_512_start|_reg_3);
   assign  _net_206 = (fpga_512_start|_reg_3);
   assign  _net_207 = (fpga_512_start|_reg_3);
   assign  _net_208 = (fpga_512_start|_reg_3);
   assign  _net_209 = (fpga_512_start|_reg_3);
   assign  _net_210 = (fpga_512_start|_reg_3);
   assign  _net_211 = (fpga_512_start|_reg_3);
   assign  _net_212 = (fpga_512_start|_reg_3);
   assign  _net_213 = (fpga_512_start|_reg_3);
   assign  _net_214 = (fpga_512_start|_reg_3);
   assign  _net_215 = (fpga_512_start|_reg_3);
   assign  _net_216 = (fpga_512_start|_reg_3);
   assign  _net_217 = (fpga_512_start|_reg_3);
   assign  _net_218 = (fpga_512_start|_reg_3);
   assign  _net_219 = (fpga_512_start|_reg_3);
   assign  _net_220 = (fpga_512_start|_reg_3);
   assign  _net_221 = (fpga_512_start|_reg_3);
   assign  _net_222 = (fpga_512_start|_reg_3);
   assign  _net_223 = (fpga_512_start|_reg_3);
   assign  _net_224 = (fpga_512_start|_reg_3);
   assign  _net_225 = (fpga_512_start|_reg_3);
   assign  _net_226 = (fpga_512_start|_reg_3);
   assign  _net_227 = (fpga_512_start|_reg_3);
   assign  _net_228 = (fpga_512_start|_reg_3);
   assign  _net_229 = (fpga_512_start|_reg_3);
   assign  _net_230 = (fpga_512_start|_reg_3);
   assign  _net_231 = (fpga_512_start|_reg_3);
   assign  _net_232 = (fpga_512_start|_reg_3);
   assign  _net_233 = (fpga_512_start|_reg_3);
   assign  _net_234 = (fpga_512_start|_reg_3);
   assign  _net_235 = (fpga_512_start|_reg_3);
   assign  _net_236 = (fpga_512_start|_reg_3);
   assign  _net_237 = (fpga_512_start|_reg_3);
   assign  _net_238 = (fpga_512_start|_reg_3);
   assign  _net_239 = (fpga_512_start|_reg_3);
   assign  _net_240 = (fpga_512_start|_reg_3);
   assign  _net_241 = (fpga_512_start|_reg_3);
   assign  _net_242 = (fpga_512_start|_reg_3);
   assign  _net_243 = (fpga_512_start|_reg_3);
   assign  _net_244 = (fpga_512_start|_reg_3);
   assign  _net_245 = (fpga_512_start|_reg_3);
   assign  _net_246 = (fpga_512_start|_reg_3);
   assign  _net_247 = (fpga_512_start|_reg_3);
   assign  _net_248 = (fpga_512_start|_reg_3);
   assign  _net_249 = (fpga_512_start|_reg_3);
   assign  _net_250 = (fpga_512_start|_reg_3);
   assign  _net_251 = (fpga_512_start|_reg_3);
   assign  _net_252 = (fpga_512_start|_reg_3);
   assign  _net_253 = (fpga_512_start|_reg_3);
   assign  _net_254 = (fpga_512_start|_reg_3);
   assign  _net_255 = (fpga_512_start|_reg_3);
   assign  _net_256 = (fpga_512_start|_reg_3);
   assign  _net_257 = (fpga_512_start|_reg_3);
   assign  _net_258 = (fpga_512_start|_reg_3);
   assign  _net_259 = (fpga_512_start|_reg_3);
   assign  _net_260 = (fpga_512_start|_reg_3);
   assign  _net_261 = (fpga_512_start|_reg_3);
   assign  _net_262 = (fpga_512_start|_reg_3);
   assign  _net_263 = (fpga_512_start|_reg_3);
   assign  _net_264 = (fpga_512_start|_reg_3);
   assign  _net_265 = (fpga_512_start|_reg_3);
   assign  _net_266 = (fpga_512_start|_reg_3);
   assign  _net_267 = (fpga_512_start|_reg_3);
   assign  _net_268 = (fpga_512_start|_reg_3);
   assign  _net_269 = (fpga_512_start|_reg_3);
   assign  _net_270 = (fpga_512_start|_reg_3);
   assign  _net_271 = (fpga_512_start|_reg_3);
   assign  _net_272 = (fpga_512_start|_reg_3);
   assign  _net_273 = (fpga_512_start|_reg_3);
   assign  _net_274 = (fpga_512_start|_reg_3);
   assign  _net_275 = (fpga_512_start|_reg_3);
   assign  _net_276 = (fpga_512_start|_reg_3);
   assign  _net_277 = (fpga_512_start|_reg_3);
   assign  _net_278 = (fpga_512_start|_reg_3);
   assign  _net_279 = (fpga_512_start|_reg_3);
   assign  _net_280 = (fpga_512_start|_reg_3);
   assign  _net_281 = (fpga_512_start|_reg_3);
   assign  _net_282 = (fpga_512_start|_reg_3);
   assign  _net_283 = (fpga_512_start|_reg_3);
   assign  _net_284 = (fpga_512_start|_reg_3);
   assign  _net_285 = (fpga_512_start|_reg_3);
   assign  _net_286 = (fpga_512_start|_reg_3);
   assign  _net_287 = (fpga_512_start|_reg_3);
   assign  _net_288 = (fpga_512_start|_reg_3);
   assign  _net_289 = (fpga_512_start|_reg_3);
   assign  _net_290 = (fpga_512_start|_reg_3);
   assign  _net_291 = (fpga_512_start|_reg_3);
   assign  _net_292 = (fpga_512_start|_reg_3);
   assign  _net_293 = (fpga_512_start|_reg_3);
   assign  _net_294 = (fpga_512_start|_reg_3);
   assign  _net_295 = (fpga_512_start|_reg_3);
   assign  _net_296 = (fpga_512_start|_reg_3);
   assign  _net_297 = (fpga_512_start|_reg_3);
   assign  _net_298 = (fpga_512_start|_reg_3);
   assign  _net_299 = (fpga_512_start|_reg_3);
   assign  _net_300 = (fpga_512_start|_reg_3);
   assign  _net_301 = (fpga_512_start|_reg_3);
   assign  _net_302 = (fpga_512_start|_reg_3);
   assign  _net_303 = (fpga_512_start|_reg_3);
   assign  _net_304 = (fpga_512_start|_reg_3);
   assign  _net_305 = (fpga_512_start|_reg_3);
   assign  _net_306 = (fpga_512_start|_reg_3);
   assign  _net_307 = (fpga_512_start|_reg_3);
   assign  _net_308 = (fpga_512_start|_reg_3);
   assign  _net_309 = (fpga_512_start|_reg_3);
   assign  _net_310 = (fpga_512_start|_reg_3);
   assign  _net_311 = (fpga_512_start|_reg_3);
   assign  _net_312 = (fpga_512_start|_reg_3);
   assign  _net_313 = (fpga_512_start|_reg_3);
   assign  _net_314 = (fpga_512_start|_reg_3);
   assign  _net_315 = (fpga_512_start|_reg_3);
   assign  _net_316 = (fpga_512_start|_reg_3);
   assign  _net_317 = (fpga_512_start|_reg_3);
   assign  _net_318 = (fpga_512_start|_reg_3);
   assign  _net_319 = (fpga_512_start|_reg_3);
   assign  _net_320 = (fpga_512_start|_reg_3);
   assign  _net_321 = (fpga_512_start|_reg_3);
   assign  _net_322 = (fpga_512_start|_reg_3);
   assign  _net_323 = (fpga_512_start|_reg_3);
   assign  _net_324 = (fpga_512_start|_reg_3);
   assign  _net_325 = (fpga_512_start|_reg_3);
   assign  _net_326 = (fpga_512_start|_reg_3);
   assign  _net_327 = (fpga_512_start|_reg_3);
   assign  _net_328 = (fpga_512_start|_reg_3);
   assign  _net_329 = (fpga_512_start|_reg_3);
   assign  _net_330 = (fpga_512_start|_reg_3);
   assign  _net_331 = (fpga_512_start|_reg_3);
   assign  _net_332 = (fpga_512_start|_reg_3);
   assign  _net_333 = (fpga_512_start|_reg_3);
   assign  _net_334 = (fpga_512_start|_reg_3);
   assign  _net_335 = (fpga_512_start|_reg_3);
   assign  _net_336 = (fpga_512_start|_reg_3);
   assign  _net_337 = (fpga_512_start|_reg_3);
   assign  _net_338 = (fpga_512_start|_reg_3);
   assign  _net_339 = (fpga_512_start|_reg_3);
   assign  _net_340 = (fpga_512_start|_reg_3);
   assign  _net_341 = (fpga_512_start|_reg_3);
   assign  _net_342 = (fpga_512_start|_reg_3);
   assign  _net_343 = (fpga_512_start|_reg_3);
   assign  _net_344 = (fpga_512_start|_reg_3);
   assign  _net_345 = (fpga_512_start|_reg_3);
   assign  _net_346 = (fpga_512_start|_reg_3);
   assign  _net_347 = (fpga_512_start|_reg_3);
   assign  _net_348 = (fpga_512_start|_reg_3);
   assign  _net_349 = (fpga_512_start|_reg_3);
   assign  _net_350 = (fpga_512_start|_reg_3);
   assign  _net_351 = (fpga_512_start|_reg_3);
   assign  _net_352 = (fpga_512_start|_reg_3);
   assign  _net_353 = (fpga_512_start|_reg_3);
   assign  _net_354 = (fpga_512_start|_reg_3);
   assign  _net_355 = (fpga_512_start|_reg_3);
   assign  _net_356 = (fpga_512_start|_reg_3);
   assign  _net_357 = (fpga_512_start|_reg_3);
   assign  _net_358 = (fpga_512_start|_reg_3);
   assign  _net_359 = (fpga_512_start|_reg_3);
   assign  _net_360 = (fpga_512_start|_reg_3);
   assign  _net_361 = (fpga_512_start|_reg_3);
   assign  _net_362 = (fpga_512_start|_reg_3);
   assign  _net_363 = (fpga_512_start|_reg_3);
   assign  _net_364 = (fpga_512_start|_reg_3);
   assign  _net_365 = (fpga_512_start|_reg_3);
   assign  _net_366 = (fpga_512_start|_reg_3);
   assign  _net_367 = (fpga_512_start|_reg_3);
   assign  _net_368 = (fpga_512_start|_reg_3);
   assign  _net_369 = (fpga_512_start|_reg_3);
   assign  _net_370 = (fpga_512_start|_reg_3);
   assign  _net_371 = (fpga_512_start|_reg_3);
   assign  _net_372 = (fpga_512_start|_reg_3);
   assign  _net_373 = (fpga_512_start|_reg_3);
   assign  _net_374 = (fpga_512_start|_reg_3);
   assign  _net_375 = (fpga_512_start|_reg_3);
   assign  _net_376 = (fpga_512_start|_reg_3);
   assign  _net_377 = (fpga_512_start|_reg_3);
   assign  _net_378 = (fpga_512_start|_reg_3);
   assign  _net_379 = (fpga_512_start|_reg_3);
   assign  _net_380 = (fpga_512_start|_reg_3);
   assign  _net_381 = (fpga_512_start|_reg_3);
   assign  _net_382 = (fpga_512_start|_reg_3);
   assign  _net_383 = (fpga_512_start|_reg_3);
   assign  _net_384 = (fpga_512_start|_reg_3);
   assign  _net_385 = (fpga_512_start|_reg_3);
   assign  _net_386 = (fpga_512_start|_reg_3);
   assign  _net_387 = (fpga_512_start|_reg_3);
   assign  _net_388 = (fpga_512_start|_reg_3);
   assign  _net_389 = (fpga_512_start|_reg_3);
   assign  _net_390 = (fpga_512_start|_reg_3);
   assign  _net_391 = (fpga_512_start|_reg_3);
   assign  _net_392 = (fpga_512_start|_reg_3);
   assign  _net_393 = (fpga_512_start|_reg_3);
   assign  _net_394 = (fpga_512_start|_reg_3);
   assign  _net_395 = (fpga_512_start|_reg_3);
   assign  _net_396 = (fpga_512_start|_reg_3);
   assign  _net_397 = (fpga_512_start|_reg_3);
   assign  _net_398 = (fpga_512_start|_reg_3);
   assign  _net_399 = (fpga_512_start|_reg_3);
   assign  _net_400 = (fpga_512_start|_reg_3);
   assign  _net_401 = (fpga_512_start|_reg_3);
   assign  _net_402 = (fpga_512_start|_reg_3);
   assign  _net_403 = (fpga_512_start|_reg_3);
   assign  _net_404 = (fpga_512_start|_reg_3);
   assign  _net_405 = (fpga_512_start|_reg_3);
   assign  _net_406 = (fpga_512_start|_reg_3);
   assign  _net_407 = (fpga_512_start|_reg_3);
   assign  _net_408 = (fpga_512_start|_reg_3);
   assign  _net_409 = (fpga_512_start|_reg_3);
   assign  _net_410 = (fpga_512_start|_reg_3);
   assign  _net_411 = (fpga_512_start|_reg_3);
   assign  _net_412 = (fpga_512_start|_reg_3);
   assign  _net_413 = (fpga_512_start|_reg_3);
   assign  _net_414 = (fpga_512_start|_reg_3);
   assign  _net_415 = (fpga_512_start|_reg_3);
   assign  _net_416 = (fpga_512_start|_reg_3);
   assign  _net_417 = (fpga_512_start|_reg_3);
   assign  _net_418 = (fpga_512_start|_reg_3);
   assign  _net_419 = (fpga_512_start|_reg_3);
   assign  _net_420 = (fpga_512_start|_reg_3);
   assign  _net_421 = (fpga_512_start|_reg_3);
   assign  _net_422 = (fpga_512_start|_reg_3);
   assign  _net_423 = (fpga_512_start|_reg_3);
   assign  _net_424 = (fpga_512_start|_reg_3);
   assign  _net_425 = (fpga_512_start|_reg_3);
   assign  _net_426 = (fpga_512_start|_reg_3);
   assign  _net_427 = (fpga_512_start|_reg_3);
   assign  _net_428 = (fpga_512_start|_reg_3);
   assign  _net_429 = (fpga_512_start|_reg_3);
   assign  _net_430 = (fpga_512_start|_reg_3);
   assign  _net_431 = (fpga_512_start|_reg_3);
   assign  _net_432 = (fpga_512_start|_reg_3);
   assign  _net_433 = (fpga_512_start|_reg_3);
   assign  _net_434 = (fpga_512_start|_reg_3);
   assign  _net_435 = (fpga_512_start|_reg_3);
   assign  _net_436 = (fpga_512_start|_reg_3);
   assign  _net_437 = (fpga_512_start|_reg_3);
   assign  _net_438 = (fpga_512_start|_reg_3);
   assign  _net_439 = (fpga_512_start|_reg_3);
   assign  _net_440 = (fpga_512_start|_reg_3);
   assign  _net_441 = (fpga_512_start|_reg_3);
   assign  _net_442 = (fpga_512_start|_reg_3);
   assign  _net_443 = (fpga_512_start|_reg_3);
   assign  _net_444 = (fpga_512_start|_reg_3);
   assign  _net_445 = (fpga_512_start|_reg_3);
   assign  _net_446 = (fpga_512_start|_reg_3);
   assign  _net_447 = (fpga_512_start|_reg_3);
   assign  _net_448 = (fpga_512_start|_reg_3);
   assign  _net_449 = (fpga_512_start|_reg_3);
   assign  _net_450 = (fpga_512_start|_reg_3);
   assign  _net_451 = (fpga_512_start|_reg_3);
   assign  _net_452 = (fpga_512_start|_reg_3);
   assign  _net_453 = (fpga_512_start|_reg_3);
   assign  _net_454 = (fpga_512_start|_reg_3);
   assign  _net_455 = (fpga_512_start|_reg_3);
   assign  _net_456 = (fpga_512_start|_reg_3);
   assign  _net_457 = (fpga_512_start|_reg_3);
   assign  _net_458 = (fpga_512_start|_reg_3);
   assign  _net_459 = (fpga_512_start|_reg_3);
   assign  _net_460 = (fpga_512_start|_reg_3);
   assign  _net_461 = (fpga_512_start|_reg_3);
   assign  _net_462 = (fpga_512_start|_reg_3);
   assign  _net_463 = (fpga_512_start|_reg_3);
   assign  _net_464 = (fpga_512_start|_reg_3);
   assign  _net_465 = (fpga_512_start|_reg_3);
   assign  _net_466 = (fpga_512_start|_reg_3);
   assign  _net_467 = (fpga_512_start|_reg_3);
   assign  _net_468 = (fpga_512_start|_reg_3);
   assign  _net_469 = (fpga_512_start|_reg_3);
   assign  _net_470 = (fpga_512_start|_reg_3);
   assign  _net_471 = (fpga_512_start|_reg_3);
   assign  _net_472 = (fpga_512_start|_reg_3);
   assign  _net_473 = (fpga_512_start|_reg_3);
   assign  _net_474 = (fpga_512_start|_reg_3);
   assign  _net_475 = (fpga_512_start|_reg_3);
   assign  _net_476 = (fpga_512_start|_reg_3);
   assign  _net_477 = (fpga_512_start|_reg_3);
   assign  _net_478 = (fpga_512_start|_reg_3);
   assign  _net_479 = (fpga_512_start|_reg_3);
   assign  _net_480 = (fpga_512_start|_reg_3);
   assign  _net_481 = (fpga_512_start|_reg_3);
   assign  _net_482 = (fpga_512_start|_reg_3);
   assign  _net_483 = (fpga_512_start|_reg_3);
   assign  _net_484 = (fpga_512_start|_reg_3);
   assign  _net_485 = (fpga_512_start|_reg_3);
   assign  _net_486 = (fpga_512_start|_reg_3);
   assign  _net_487 = (fpga_512_start|_reg_3);
   assign  _net_488 = (fpga_512_start|_reg_3);
   assign  _net_489 = (fpga_512_start|_reg_3);
   assign  _net_490 = (fpga_512_start|_reg_3);
   assign  _net_491 = (fpga_512_start|_reg_3);
   assign  _net_492 = (fpga_512_start|_reg_3);
   assign  _net_493 = (fpga_512_start|_reg_3);
   assign  _net_494 = (fpga_512_start|_reg_3);
   assign  _net_495 = (fpga_512_start|_reg_3);
   assign  _net_496 = (fpga_512_start|_reg_3);
   assign  _net_497 = (fpga_512_start|_reg_3);
   assign  _net_498 = (fpga_512_start|_reg_3);
   assign  _net_499 = (fpga_512_start|_reg_3);
   assign  _net_500 = (fpga_512_start|_reg_3);
   assign  _net_501 = (fpga_512_start|_reg_3);
   assign  _net_502 = (fpga_512_start|_reg_3);
   assign  _net_503 = (fpga_512_start|_reg_3);
   assign  _net_504 = (fpga_512_start|_reg_3);
   assign  _net_505 = (fpga_512_start|_reg_3);
   assign  _net_506 = (fpga_512_start|_reg_3);
   assign  _net_507 = (fpga_512_start|_reg_3);
   assign  _net_508 = (fpga_512_start|_reg_3);
   assign  _net_509 = (fpga_512_start|_reg_3);
   assign  _net_510 = (fpga_512_start|_reg_3);
   assign  _net_511 = (fpga_512_start|_reg_3);
   assign  _net_512 = (fpga_512_start|_reg_3);
   assign  _net_513 = (fpga_512_start|_reg_3);
   assign  _net_514 = (fpga_512_start|_reg_3);
   assign  _net_515 = (fpga_512_start|_reg_3);
   assign  _net_516 = (fpga_512_start|_reg_3);

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_meirotest_end_meiro)
    begin
    $finish;
    end
  end

// synthesis translate_on
// synopsys translate_on
   assign  HEX0 = _meirotest_end_meiro;
initial begin
    map_test[0] = 10'b1111111111;
    map_test[1] = 10'b1111111111;
    map_test[2] = 10'b1111111111;
    map_test[3] = 10'b1111111111;
    map_test[4] = 10'b1111111111;
    map_test[5] = 10'b1111111111;
    map_test[6] = 10'b1111111111;
    map_test[7] = 10'b1111111111;
    map_test[8] = 10'b1111111111;
    map_test[9] = 10'b1111111111;
    map_test[10] = 10'b1111111111;
    map_test[11] = 10'b1111111111;
    map_test[12] = 10'b1111111111;
    map_test[13] = 10'b1111111111;
    map_test[14] = 10'b1111111111;
    map_test[15] = 10'b1111111111;
    map_test[16] = 10'b1111111111;
    map_test[17] = 10'b1111111111;
    map_test[18] = 10'b1111111111;
    map_test[19] = 10'b1111111111;
    map_test[20] = 10'b1111111111;
    map_test[21] = 10'b1111111111;
    map_test[22] = 10'b1111111111;
    map_test[23] = 10'b1111111111;
    map_test[24] = 10'b1111111111;
    map_test[25] = 10'b1111111111;
    map_test[26] = 10'b1111111111;
    map_test[27] = 10'b1111111111;
    map_test[28] = 10'b1111111111;
    map_test[29] = 10'b1111111111;
    map_test[30] = 10'b1111111111;
    map_test[31] = 10'b1111111111;
    map_test[32] = 10'b1111111111;
    map_test[33] = 10'b0100000000;
    map_test[34] = 10'b0111111111;
    map_test[35] = 10'b0100000000;
    map_test[36] = 10'b0100000000;
    map_test[37] = 10'b0100000000;
    map_test[38] = 10'b0000000000;
    map_test[39] = 10'b0100000000;
    map_test[40] = 10'b1111111111;
    map_test[41] = 10'b0100000000;
    map_test[42] = 10'b0100000000;
    map_test[43] = 10'b0100000000;
    map_test[44] = 10'b0100000000;
    map_test[45] = 10'b0100000000;
    map_test[46] = 10'b0100000000;
    map_test[47] = 10'b0100000000;
    map_test[48] = 10'b1111111111;
    map_test[49] = 10'b0100000000;
    map_test[50] = 10'b0100000000;
    map_test[51] = 10'b0100000000;
    map_test[52] = 10'b0100000000;
    map_test[53] = 10'b0100000000;
    map_test[54] = 10'b0100000000;
    map_test[55] = 10'b0100000000;
    map_test[56] = 10'b1111111111;
    map_test[57] = 10'b0100000000;
    map_test[58] = 10'b0100000000;
    map_test[59] = 10'b0100000000;
    map_test[60] = 10'b1111111111;
    map_test[61] = 10'b0100000000;
    map_test[62] = 10'b0100000000;
    map_test[63] = 10'b1111111111;
    map_test[64] = 10'b1111111111;
    map_test[65] = 10'b0100000000;
    map_test[66] = 10'b1111111111;
    map_test[67] = 10'b0100000000;
    map_test[68] = 10'b1111111111;
    map_test[69] = 10'b1111111111;
    map_test[70] = 10'b1111111111;
    map_test[71] = 10'b0100000000;
    map_test[72] = 10'b1111111111;
    map_test[73] = 10'b0100000000;
    map_test[74] = 10'b1111111111;
    map_test[75] = 10'b1111111111;
    map_test[76] = 10'b1111111111;
    map_test[77] = 10'b0100000000;
    map_test[78] = 10'b1111111111;
    map_test[79] = 10'b0100000000;
    map_test[80] = 10'b1111111111;
    map_test[81] = 10'b0100000000;
    map_test[82] = 10'b1111111111;
    map_test[83] = 10'b1111111111;
    map_test[84] = 10'b1111111111;
    map_test[85] = 10'b0100000000;
    map_test[86] = 10'b1111111111;
    map_test[87] = 10'b0100000000;
    map_test[88] = 10'b1111111111;
    map_test[89] = 10'b0100000000;
    map_test[90] = 10'b1111111111;
    map_test[91] = 10'b0100000000;
    map_test[92] = 10'b1111111111;
    map_test[93] = 10'b0100000000;
    map_test[94] = 10'b1111111111;
    map_test[95] = 10'b1111111111;
    map_test[96] = 10'b1111111111;
    map_test[97] = 10'b0100000000;
    map_test[98] = 10'b1111111111;
    map_test[99] = 10'b0100000000;
    map_test[100] = 10'b1111111111;
    map_test[101] = 10'b0100000000;
    map_test[102] = 10'b1111111111;
    map_test[103] = 10'b0100000000;
    map_test[104] = 10'b1111111111;
    map_test[105] = 10'b0100000000;
    map_test[106] = 10'b0100000000;
    map_test[107] = 10'b0100000000;
    map_test[108] = 10'b1111111111;
    map_test[109] = 10'b0100000000;
    map_test[110] = 10'b1111111111;
    map_test[111] = 10'b0100000000;
    map_test[112] = 10'b1111111111;
    map_test[113] = 10'b0100000000;
    map_test[114] = 10'b1111111111;
    map_test[115] = 10'b0100000000;
    map_test[116] = 10'b0100000000;
    map_test[117] = 10'b0100000000;
    map_test[118] = 10'b1111111111;
    map_test[119] = 10'b0100000000;
    map_test[120] = 10'b1111111111;
    map_test[121] = 10'b0100000000;
    map_test[122] = 10'b1111111111;
    map_test[123] = 10'b0100000000;
    map_test[124] = 10'b1111111111;
    map_test[125] = 10'b0100000000;
    map_test[126] = 10'b1111111111;
    map_test[127] = 10'b1111111111;
    map_test[128] = 10'b1111111111;
    map_test[129] = 10'b1111111111;
    map_test[130] = 10'b1111111111;
    map_test[131] = 10'b0100000000;
    map_test[132] = 10'b1111111111;
    map_test[133] = 10'b0100000000;
    map_test[134] = 10'b1111111111;
    map_test[135] = 10'b0100000000;
    map_test[136] = 10'b1111111111;
    map_test[137] = 10'b1111111111;
    map_test[138] = 10'b1111111111;
    map_test[139] = 10'b0100000000;
    map_test[140] = 10'b1111111111;
    map_test[141] = 10'b0100000000;
    map_test[142] = 10'b1111111111;
    map_test[143] = 10'b0100000000;
    map_test[144] = 10'b1111111111;
    map_test[145] = 10'b1111111111;
    map_test[146] = 10'b1111111111;
    map_test[147] = 10'b0100000000;
    map_test[148] = 10'b1111111111;
    map_test[149] = 10'b1111111111;
    map_test[150] = 10'b1111111111;
    map_test[151] = 10'b0100000000;
    map_test[152] = 10'b1111111111;
    map_test[153] = 10'b0100000000;
    map_test[154] = 10'b1111111111;
    map_test[155] = 10'b0100000000;
    map_test[156] = 10'b1111111111;
    map_test[157] = 10'b0100000000;
    map_test[158] = 10'b1111111111;
    map_test[159] = 10'b1111111111;
    map_test[160] = 10'b1111111111;
    map_test[161] = 10'b0100000000;
    map_test[162] = 10'b0100000000;
    map_test[163] = 10'b0100000000;
    map_test[164] = 10'b1111111111;
    map_test[165] = 10'b0100000000;
    map_test[166] = 10'b1111111111;
    map_test[167] = 10'b0100000000;
    map_test[168] = 10'b0100000000;
    map_test[169] = 10'b0100000000;
    map_test[170] = 10'b1111111111;
    map_test[171] = 10'b0100000000;
    map_test[172] = 10'b1111111111;
    map_test[173] = 10'b0100000000;
    map_test[174] = 10'b1111111111;
    map_test[175] = 10'b0100000000;
    map_test[176] = 10'b0100000000;
    map_test[177] = 10'b0100000000;
    map_test[178] = 10'b1111111111;
    map_test[179] = 10'b0100000000;
    map_test[180] = 10'b0100000000;
    map_test[181] = 10'b0100000000;
    map_test[182] = 10'b1111111111;
    map_test[183] = 10'b0100000000;
    map_test[184] = 10'b1111111111;
    map_test[185] = 10'b0100000000;
    map_test[186] = 10'b1111111111;
    map_test[187] = 10'b0100000000;
    map_test[188] = 10'b0100000000;
    map_test[189] = 10'b0100000000;
    map_test[190] = 10'b1111111111;
    map_test[191] = 10'b1111111111;
    map_test[192] = 10'b1111111111;
    map_test[193] = 10'b0100000000;
    map_test[194] = 10'b1111111111;
    map_test[195] = 10'b1111111111;
    map_test[196] = 10'b1111111111;
    map_test[197] = 10'b0100000000;
    map_test[198] = 10'b1111111111;
    map_test[199] = 10'b0100000000;
    map_test[200] = 10'b1111111111;
    map_test[201] = 10'b1111111111;
    map_test[202] = 10'b1111111111;
    map_test[203] = 10'b0100000000;
    map_test[204] = 10'b1111111111;
    map_test[205] = 10'b0100000000;
    map_test[206] = 10'b1111111111;
    map_test[207] = 10'b1111111111;
    map_test[208] = 10'b1111111111;
    map_test[209] = 10'b0100000000;
    map_test[210] = 10'b1111111111;
    map_test[211] = 10'b0100000000;
    map_test[212] = 10'b1111111111;
    map_test[213] = 10'b0100000000;
    map_test[214] = 10'b1111111111;
    map_test[215] = 10'b1111111111;
    map_test[216] = 10'b1111111111;
    map_test[217] = 10'b1111111111;
    map_test[218] = 10'b1111111111;
    map_test[219] = 10'b1111111111;
    map_test[220] = 10'b1111111111;
    map_test[221] = 10'b0100000000;
    map_test[222] = 10'b1111111111;
    map_test[223] = 10'b1111111111;
    map_test[224] = 10'b1111111111;
    map_test[225] = 10'b0100000000;
    map_test[226] = 10'b0100000000;
    map_test[227] = 10'b0100000000;
    map_test[228] = 10'b1111111111;
    map_test[229] = 10'b0100000000;
    map_test[230] = 10'b0100000000;
    map_test[231] = 10'b0100000000;
    map_test[232] = 10'b1111111111;
    map_test[233] = 10'b0100000000;
    map_test[234] = 10'b0100000000;
    map_test[235] = 10'b0100000000;
    map_test[236] = 10'b1111111111;
    map_test[237] = 10'b0100000000;
    map_test[238] = 10'b1111111111;
    map_test[239] = 10'b0100000000;
    map_test[240] = 10'b0100000000;
    map_test[241] = 10'b0100000000;
    map_test[242] = 10'b1111111111;
    map_test[243] = 10'b0100000000;
    map_test[244] = 10'b1111111111;
    map_test[245] = 10'b0100000000;
    map_test[246] = 10'b0100000000;
    map_test[247] = 10'b0100000000;
    map_test[248] = 10'b0100000000;
    map_test[249] = 10'b0100000000;
    map_test[250] = 10'b0100000000;
    map_test[251] = 10'b0100000000;
    map_test[252] = 10'b1111111111;
    map_test[253] = 10'b0100000000;
    map_test[254] = 10'b0100000000;
    map_test[255] = 10'b1111111111;
    map_test[256] = 10'b1111111111;
    map_test[257] = 10'b0100000000;
    map_test[258] = 10'b1111111111;
    map_test[259] = 10'b0100000000;
    map_test[260] = 10'b1111111111;
    map_test[261] = 10'b0100000000;
    map_test[262] = 10'b1111111111;
    map_test[263] = 10'b1111111111;
    map_test[264] = 10'b1111111111;
    map_test[265] = 10'b0100000000;
    map_test[266] = 10'b1111111111;
    map_test[267] = 10'b1111111111;
    map_test[268] = 10'b1111111111;
    map_test[269] = 10'b0100000000;
    map_test[270] = 10'b1111111111;
    map_test[271] = 10'b0100000000;
    map_test[272] = 10'b1111111111;
    map_test[273] = 10'b1111111111;
    map_test[274] = 10'b1111111111;
    map_test[275] = 10'b1111111111;
    map_test[276] = 10'b1111111111;
    map_test[277] = 10'b1111111111;
    map_test[278] = 10'b1111111111;
    map_test[279] = 10'b0100000000;
    map_test[280] = 10'b1111111111;
    map_test[281] = 10'b1111111111;
    map_test[282] = 10'b1111111111;
    map_test[283] = 10'b1111111111;
    map_test[284] = 10'b1111111111;
    map_test[285] = 10'b0100000000;
    map_test[286] = 10'b1111111111;
    map_test[287] = 10'b1111111111;
    map_test[288] = 10'b1111111111;
    map_test[289] = 10'b0100000000;
    map_test[290] = 10'b1111111111;
    map_test[291] = 10'b0100000000;
    map_test[292] = 10'b1111111111;
    map_test[293] = 10'b0100000000;
    map_test[294] = 10'b1111111111;
    map_test[295] = 10'b0100000000;
    map_test[296] = 10'b0100000000;
    map_test[297] = 10'b0100000000;
    map_test[298] = 10'b1111111111;
    map_test[299] = 10'b0100000000;
    map_test[300] = 10'b0100000000;
    map_test[301] = 10'b0100000000;
    map_test[302] = 10'b1111111111;
    map_test[303] = 10'b0100000000;
    map_test[304] = 10'b0100000000;
    map_test[305] = 10'b0100000000;
    map_test[306] = 10'b0100000000;
    map_test[307] = 10'b0100000000;
    map_test[308] = 10'b0100000000;
    map_test[309] = 10'b0100000000;
    map_test[310] = 10'b0100000000;
    map_test[311] = 10'b0100000000;
    map_test[312] = 10'b1111111111;
    map_test[313] = 10'b0100000000;
    map_test[314] = 10'b0100000000;
    map_test[315] = 10'b0100000000;
    map_test[316] = 10'b0100000000;
    map_test[317] = 10'b0100000000;
    map_test[318] = 10'b0100000000;
    map_test[319] = 10'b1111111111;
    map_test[320] = 10'b1111111111;
    map_test[321] = 10'b0100000000;
    map_test[322] = 10'b1111111111;
    map_test[323] = 10'b0100000000;
    map_test[324] = 10'b1111111111;
    map_test[325] = 10'b1111111111;
    map_test[326] = 10'b1111111111;
    map_test[327] = 10'b0100000000;
    map_test[328] = 10'b1111111111;
    map_test[329] = 10'b1111111111;
    map_test[330] = 10'b1111111111;
    map_test[331] = 10'b0100000000;
    map_test[332] = 10'b1111111111;
    map_test[333] = 10'b0100000000;
    map_test[334] = 10'b1111111111;
    map_test[335] = 10'b1111111111;
    map_test[336] = 10'b1111111111;
    map_test[337] = 10'b1111111111;
    map_test[338] = 10'b1111111111;
    map_test[339] = 10'b1111111111;
    map_test[340] = 10'b1111111111;
    map_test[341] = 10'b0100000000;
    map_test[342] = 10'b1111111111;
    map_test[343] = 10'b1111111111;
    map_test[344] = 10'b1111111111;
    map_test[345] = 10'b0100000000;
    map_test[346] = 10'b1111111111;
    map_test[347] = 10'b1111111111;
    map_test[348] = 10'b1111111111;
    map_test[349] = 10'b1111111111;
    map_test[350] = 10'b0100000000;
    map_test[351] = 10'b1111111111;
    map_test[352] = 10'b1111111111;
    map_test[353] = 10'b0100000000;
    map_test[354] = 10'b1111111111;
    map_test[355] = 10'b0100000000;
    map_test[356] = 10'b1111111111;
    map_test[357] = 10'b0100000000;
    map_test[358] = 10'b0100000000;
    map_test[359] = 10'b0100000000;
    map_test[360] = 10'b1111111111;
    map_test[361] = 10'b0100000000;
    map_test[362] = 10'b0100000000;
    map_test[363] = 10'b0100000000;
    map_test[364] = 10'b1111111111;
    map_test[365] = 10'b0100000000;
    map_test[366] = 10'b1111111111;
    map_test[367] = 10'b0100000000;
    map_test[368] = 10'b0100000000;
    map_test[369] = 10'b0100000000;
    map_test[370] = 10'b1111111111;
    map_test[371] = 10'b0100000000;
    map_test[372] = 10'b0100000000;
    map_test[373] = 10'b0100000000;
    map_test[374] = 10'b1111111111;
    map_test[375] = 10'b0100000000;
    map_test[376] = 10'b0100000000;
    map_test[377] = 10'b0100000000;
    map_test[378] = 10'b1111111111;
    map_test[379] = 10'b0100000000;
    map_test[380] = 10'b0100000000;
    map_test[381] = 10'b0100000000;
    map_test[382] = 10'b0100000000;
    map_test[383] = 10'b1111111111;
    map_test[384] = 10'b1111111111;
    map_test[385] = 10'b0100000000;
    map_test[386] = 10'b1111111111;
    map_test[387] = 10'b0100000000;
    map_test[388] = 10'b1111111111;
    map_test[389] = 10'b0100000000;
    map_test[390] = 10'b1111111111;
    map_test[391] = 10'b1111111111;
    map_test[392] = 10'b1111111111;
    map_test[393] = 10'b0100000000;
    map_test[394] = 10'b1111111111;
    map_test[395] = 10'b0100000000;
    map_test[396] = 10'b1111111111;
    map_test[397] = 10'b1111111111;
    map_test[398] = 10'b1111111111;
    map_test[399] = 10'b0100000000;
    map_test[400] = 10'b1111111111;
    map_test[401] = 10'b0100000000;
    map_test[402] = 10'b1111111111;
    map_test[403] = 10'b1111111111;
    map_test[404] = 10'b1111111111;
    map_test[405] = 10'b1111111111;
    map_test[406] = 10'b1111111111;
    map_test[407] = 10'b0100000000;
    map_test[408] = 10'b1111111111;
    map_test[409] = 10'b1111111111;
    map_test[410] = 10'b1111111111;
    map_test[411] = 10'b0100000000;
    map_test[412] = 10'b1111111111;
    map_test[413] = 10'b1111111111;
    map_test[414] = 10'b1111111111;
    map_test[415] = 10'b1111111111;
    map_test[416] = 10'b1111111111;
    map_test[417] = 10'b0100000000;
    map_test[418] = 10'b1111111111;
    map_test[419] = 10'b0100000000;
    map_test[420] = 10'b1111111111;
    map_test[421] = 10'b0100000000;
    map_test[422] = 10'b1111111111;
    map_test[423] = 10'b0100000000;
    map_test[424] = 10'b1111111111;
    map_test[425] = 10'b0100000000;
    map_test[426] = 10'b1111111111;
    map_test[427] = 10'b0100000000;
    map_test[428] = 10'b1111111111;
    map_test[429] = 10'b0100000000;
    map_test[430] = 10'b1111111111;
    map_test[431] = 10'b0100000000;
    map_test[432] = 10'b1111111111;
    map_test[433] = 10'b0100000000;
    map_test[434] = 10'b0100000000;
    map_test[435] = 10'b0100000000;
    map_test[436] = 10'b0100000000;
    map_test[437] = 10'b0100000000;
    map_test[438] = 10'b0100000000;
    map_test[439] = 10'b0100000000;
    map_test[440] = 10'b1111111111;
    map_test[441] = 10'b0100000000;
    map_test[442] = 10'b1111111111;
    map_test[443] = 10'b0100000000;
    map_test[444] = 10'b1111111111;
    map_test[445] = 10'b0100000000;
    map_test[446] = 10'b1111111111;
    map_test[447] = 10'b1111111111;
    map_test[448] = 10'b1111111111;
    map_test[449] = 10'b0100000000;
    map_test[450] = 10'b1111111111;
    map_test[451] = 10'b0100000000;
    map_test[452] = 10'b0100000000;
    map_test[453] = 10'b0100000000;
    map_test[454] = 10'b0100000000;
    map_test[455] = 10'b0100000000;
    map_test[456] = 10'b1111111111;
    map_test[457] = 10'b0100000000;
    map_test[458] = 10'b0100000000;
    map_test[459] = 10'b0100000000;
    map_test[460] = 10'b0100000000;
    map_test[461] = 10'b0100000000;
    map_test[462] = 10'b0100000000;
    map_test[463] = 10'b0100000000;
    map_test[464] = 10'b0100000000;
    map_test[465] = 10'b1111111111;
    map_test[466] = 10'b1111111111;
    map_test[467] = 10'b1111111111;
    map_test[468] = 10'b1111111111;
    map_test[469] = 10'b0100000000;
    map_test[470] = 10'b1111111111;
    map_test[471] = 10'b0100000000;
    map_test[472] = 10'b0100000000;
    map_test[473] = 10'b0100000000;
    map_test[474] = 10'b0100000000;
    map_test[475] = 10'b0100000000;
    map_test[476] = 10'b0100000000;
    map_test[477] = 10'b0100000000;
    map_test[478] = 10'b1111111111;
    map_test[479] = 10'b1111111111;
    map_test[480] = 10'b1111111111;
    map_test[481] = 10'b1111111111;
    map_test[482] = 10'b1111111111;
    map_test[483] = 10'b1111111111;
    map_test[484] = 10'b1111111111;
    map_test[485] = 10'b1111111111;
    map_test[486] = 10'b1111111111;
    map_test[487] = 10'b1111111111;
    map_test[488] = 10'b1111111111;
    map_test[489] = 10'b1111111111;
    map_test[490] = 10'b1111111111;
    map_test[491] = 10'b1111111111;
    map_test[492] = 10'b1111111111;
    map_test[493] = 10'b1111111111;
    map_test[494] = 10'b1111111111;
    map_test[495] = 10'b1111111111;
    map_test[496] = 10'b1111111111;
    map_test[497] = 10'b1111111111;
    map_test[498] = 10'b1111111111;
    map_test[499] = 10'b1111111111;
    map_test[500] = 10'b1111111111;
    map_test[501] = 10'b1111111111;
    map_test[502] = 10'b1111111111;
    map_test[503] = 10'b1111111111;
    map_test[504] = 10'b1111111111;
    map_test[505] = 10'b1111111111;
    map_test[506] = 10'b1111111111;
    map_test[507] = 10'b1111111111;
    map_test[508] = 10'b1111111111;
    map_test[509] = 10'b1111111111;
    map_test[510] = 10'b1111111111;
    map_test[511] = 10'b1111111111;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     out_put_flag <= 1'b0;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     first <= 4'b0000;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     second <= 4'b0000;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     third <= 4'b0000;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     count <= 32'b00000000000000000000000000000000;
end
initial begin
    encode[0] = 8'b00111111;
    encode[1] = 8'b00000110;
    encode[2] = 8'b01011011;
    encode[3] = 8'b01001111;
    encode[4] = 8'b01100110;
    encode[5] = 8'b01101101;
    encode[6] = 8'b01111101;
    encode[7] = 8'b00100111;
    encode[8] = 8'b01111111;
    encode[9] = 8'b01101111;
    encode[10] = 8'b01110111;
    encode[11] = 8'b01111100;
    encode[12] = 8'b00111001;
    encode[13] = 8'b01011110;
    encode[14] = 8'b01111001;
    encode[15] = 8'b01110001;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     end_reg <= 2'b00;
else if ((_net_1)|(_net_0)) 
      end_reg <= ((_net_1) ?(end_reg+2'b01):2'b0)|
    ((_net_0) ?2'b10:2'b0);

end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_3 <= 1'b0;
else if ((_reg_3)) 
      _reg_3 <= 1'b0;
end
endmodule

/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 19:04:52 2023
 Licensed to :EVALUATION USER*/
