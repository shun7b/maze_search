
/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Wed Dec 28 07:19:22 2022
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module subs ( p_reset , m_clock , data_in33 , data_in35 , data_in37 , data_in39 , data_in41 , data_in43 , data_in45 , data_in47 , data_in49 , data_in51 , data_in53 , data_in55 , data_in57 , data_in59 , data_in61 , data_in65 , data_in67 , data_in69 , data_in71 , data_in73 , data_in75 , data_in77 , data_in79 , data_in81 , data_in83 , data_in85 , data_in87 , data_in89 , data_in91 , data_in93 , data_in97 , data_in99 , data_in101 , data_in103 , data_in105 , data_in107 , data_in109 , data_in111 , data_in113 , data_in115 , data_in117 , data_in119 , data_in121 , data_in123 , data_in125 , data_in129 , data_in131 , data_in133 , data_in135 , data_in137 , data_in139 , data_in141 , data_in143 , data_in145 , data_in147 , data_in149 , data_in151 , data_in153 , data_in155 , data_in157 , data_in161 , data_in163 , data_in165 , data_in167 , data_in169 , data_in171 , data_in173 , data_in175 , data_in177 , data_in179 , data_in181 , data_in183 , data_in185 , data_in187 , data_in189 , data_in193 , data_in195 , data_in197 , data_in199 , data_in201 , data_in203 , data_in205 , data_in207 , data_in209 , data_in211 , data_in213 , data_in215 , data_in217 , data_in219 , data_in221 , data_in225 , data_in227 , data_in229 , data_in231 , data_in233 , data_in235 , data_in237 , data_in239 , data_in241 , data_in243 , data_in245 , data_in247 , data_in249 , data_in251 , data_in253 , data_in257 , data_in259 , data_in261 , data_in263 , data_in265 , data_in267 , data_in269 , data_in271 , data_in273 , data_in275 , data_in277 , data_in279 , data_in281 , data_in283 , data_in285 , data_in289 , data_in291 , data_in293 , data_in295 , data_in297 , data_in299 , data_in301 , data_in303 , data_in305 , data_in307 , data_in309 , data_in311 , data_in313 , data_in315 , data_in317 , data_in321 , data_in323 , data_in325 , data_in327 , data_in329 , data_in331 , data_in333 , data_in335 , data_in337 , data_in339 , data_in341 , data_in343 , data_in345 , data_in347 , data_in349 , data_in353 , data_in355 , data_in357 , data_in359 , data_in361 , data_in363 , data_in365 , data_in367 , data_in369 , data_in371 , data_in373 , data_in375 , data_in377 , data_in379 , data_in381 , data_in385 , data_in387 , data_in389 , data_in391 , data_in393 , data_in395 , data_in397 , data_in399 , data_in401 , data_in403 , data_in405 , data_in407 , data_in409 , data_in411 , data_in413 , data_in417 , data_in419 , data_in421 , data_in423 , data_in425 , data_in427 , data_in429 , data_in431 , data_in433 , data_in435 , data_in437 , data_in439 , data_in441 , data_in443 , data_in445 , data_in449 , data_in451 , data_in453 , data_in455 , data_in457 , data_in459 , data_in461 , data_in463 , data_in465 , data_in467 , data_in469 , data_in471 , data_in473 , data_in475 , data_in477 , data_in_index33 , data_in_index35 , data_in_index37 , data_in_index39 , data_in_index41 , data_in_index43 , data_in_index45 , data_in_index47 , data_in_index49 , data_in_index51 , data_in_index53 , data_in_index55 , data_in_index57 , data_in_index59 , data_in_index61 , data_in_index65 , data_in_index67 , data_in_index69 , data_in_index71 , data_in_index73 , data_in_index75 , data_in_index77 , data_in_index79 , data_in_index81 , data_in_index83 , data_in_index85 , data_in_index87 , data_in_index89 , data_in_index91 , data_in_index93 , data_in_index97 , data_in_index99 , data_in_index101 , data_in_index103 , data_in_index105 , data_in_index107 , data_in_index109 , data_in_index111 , data_in_index113 , data_in_index115 , data_in_index117 , data_in_index119 , data_in_index121 , data_in_index123 , data_in_index125 , data_in_index129 , data_in_index131 , data_in_index133 , data_in_index135 , data_in_index137 , data_in_index139 , data_in_index141 , data_in_index143 , data_in_index145 , data_in_index147 , data_in_index149 , data_in_index151 , data_in_index153 , data_in_index155 , data_in_index157 , data_in_index161 , data_in_index163 , data_in_index165 , data_in_index167 , data_in_index169 , data_in_index171 , data_in_index173 , data_in_index175 , data_in_index177 , data_in_index179 , data_in_index181 , data_in_index183 , data_in_index185 , data_in_index187 , data_in_index189 , data_in_index193 , data_in_index195 , data_in_index197 , data_in_index199 , data_in_index201 , data_in_index203 , data_in_index205 , data_in_index207 , data_in_index209 , data_in_index211 , data_in_index213 , data_in_index215 , data_in_index217 , data_in_index219 , data_in_index221 , data_in_index225 , data_in_index227 , data_in_index229 , data_in_index231 , data_in_index233 , data_in_index235 , data_in_index237 , data_in_index239 , data_in_index241 , data_in_index243 , data_in_index245 , data_in_index247 , data_in_index249 , data_in_index251 , data_in_index253 , data_in_index257 , data_in_index259 , data_in_index261 , data_in_index263 , data_in_index265 , data_in_index267 , data_in_index269 , data_in_index271 , data_in_index273 , data_in_index275 , data_in_index277 , data_in_index279 , data_in_index281 , data_in_index283 , data_in_index285 , data_in_index289 , data_in_index291 , data_in_index293 , data_in_index295 , data_in_index297 , data_in_index299 , data_in_index301 , data_in_index303 , data_in_index305 , data_in_index307 , data_in_index309 , data_in_index311 , data_in_index313 , data_in_index315 , data_in_index317 , data_in_index321 , data_in_index323 , data_in_index325 , data_in_index327 , data_in_index329 , data_in_index331 , data_in_index333 , data_in_index335 , data_in_index337 , data_in_index339 , data_in_index341 , data_in_index343 , data_in_index345 , data_in_index347 , data_in_index349 , data_in_index353 , data_in_index355 , data_in_index357 , data_in_index359 , data_in_index361 , data_in_index363 , data_in_index365 , data_in_index367 , data_in_index369 , data_in_index371 , data_in_index373 , data_in_index375 , data_in_index377 , data_in_index379 , data_in_index381 , data_in_index385 , data_in_index387 , data_in_index389 , data_in_index391 , data_in_index393 , data_in_index395 , data_in_index397 , data_in_index399 , data_in_index401 , data_in_index403 , data_in_index405 , data_in_index407 , data_in_index409 , data_in_index411 , data_in_index413 , data_in_index417 , data_in_index419 , data_in_index421 , data_in_index423 , data_in_index425 , data_in_index427 , data_in_index429 , data_in_index431 , data_in_index433 , data_in_index435 , data_in_index437 , data_in_index439 , data_in_index441 , data_in_index443 , data_in_index445 , data_in_index449 , data_in_index451 , data_in_index453 , data_in_index455 , data_in_index457 , data_in_index459 , data_in_index461 , data_in_index463 , data_in_index465 , data_in_index467 , data_in_index469 , data_in_index471 , data_in_index473 , data_in_index475 , data_in_index477 , sub_array_out , subs_exe );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input [9:0] data_in33;
  wire [9:0] data_in33;
  input [9:0] data_in35;
  wire [9:0] data_in35;
  input [9:0] data_in37;
  wire [9:0] data_in37;
  input [9:0] data_in39;
  wire [9:0] data_in39;
  input [9:0] data_in41;
  wire [9:0] data_in41;
  input [9:0] data_in43;
  wire [9:0] data_in43;
  input [9:0] data_in45;
  wire [9:0] data_in45;
  input [9:0] data_in47;
  wire [9:0] data_in47;
  input [9:0] data_in49;
  wire [9:0] data_in49;
  input [9:0] data_in51;
  wire [9:0] data_in51;
  input [9:0] data_in53;
  wire [9:0] data_in53;
  input [9:0] data_in55;
  wire [9:0] data_in55;
  input [9:0] data_in57;
  wire [9:0] data_in57;
  input [9:0] data_in59;
  wire [9:0] data_in59;
  input [9:0] data_in61;
  wire [9:0] data_in61;
  input [9:0] data_in65;
  wire [9:0] data_in65;
  input [9:0] data_in67;
  wire [9:0] data_in67;
  input [9:0] data_in69;
  wire [9:0] data_in69;
  input [9:0] data_in71;
  wire [9:0] data_in71;
  input [9:0] data_in73;
  wire [9:0] data_in73;
  input [9:0] data_in75;
  wire [9:0] data_in75;
  input [9:0] data_in77;
  wire [9:0] data_in77;
  input [9:0] data_in79;
  wire [9:0] data_in79;
  input [9:0] data_in81;
  wire [9:0] data_in81;
  input [9:0] data_in83;
  wire [9:0] data_in83;
  input [9:0] data_in85;
  wire [9:0] data_in85;
  input [9:0] data_in87;
  wire [9:0] data_in87;
  input [9:0] data_in89;
  wire [9:0] data_in89;
  input [9:0] data_in91;
  wire [9:0] data_in91;
  input [9:0] data_in93;
  wire [9:0] data_in93;
  input [9:0] data_in97;
  wire [9:0] data_in97;
  input [9:0] data_in99;
  wire [9:0] data_in99;
  input [9:0] data_in101;
  wire [9:0] data_in101;
  input [9:0] data_in103;
  wire [9:0] data_in103;
  input [9:0] data_in105;
  wire [9:0] data_in105;
  input [9:0] data_in107;
  wire [9:0] data_in107;
  input [9:0] data_in109;
  wire [9:0] data_in109;
  input [9:0] data_in111;
  wire [9:0] data_in111;
  input [9:0] data_in113;
  wire [9:0] data_in113;
  input [9:0] data_in115;
  wire [9:0] data_in115;
  input [9:0] data_in117;
  wire [9:0] data_in117;
  input [9:0] data_in119;
  wire [9:0] data_in119;
  input [9:0] data_in121;
  wire [9:0] data_in121;
  input [9:0] data_in123;
  wire [9:0] data_in123;
  input [9:0] data_in125;
  wire [9:0] data_in125;
  input [9:0] data_in129;
  wire [9:0] data_in129;
  input [9:0] data_in131;
  wire [9:0] data_in131;
  input [9:0] data_in133;
  wire [9:0] data_in133;
  input [9:0] data_in135;
  wire [9:0] data_in135;
  input [9:0] data_in137;
  wire [9:0] data_in137;
  input [9:0] data_in139;
  wire [9:0] data_in139;
  input [9:0] data_in141;
  wire [9:0] data_in141;
  input [9:0] data_in143;
  wire [9:0] data_in143;
  input [9:0] data_in145;
  wire [9:0] data_in145;
  input [9:0] data_in147;
  wire [9:0] data_in147;
  input [9:0] data_in149;
  wire [9:0] data_in149;
  input [9:0] data_in151;
  wire [9:0] data_in151;
  input [9:0] data_in153;
  wire [9:0] data_in153;
  input [9:0] data_in155;
  wire [9:0] data_in155;
  input [9:0] data_in157;
  wire [9:0] data_in157;
  input [9:0] data_in161;
  wire [9:0] data_in161;
  input [9:0] data_in163;
  wire [9:0] data_in163;
  input [9:0] data_in165;
  wire [9:0] data_in165;
  input [9:0] data_in167;
  wire [9:0] data_in167;
  input [9:0] data_in169;
  wire [9:0] data_in169;
  input [9:0] data_in171;
  wire [9:0] data_in171;
  input [9:0] data_in173;
  wire [9:0] data_in173;
  input [9:0] data_in175;
  wire [9:0] data_in175;
  input [9:0] data_in177;
  wire [9:0] data_in177;
  input [9:0] data_in179;
  wire [9:0] data_in179;
  input [9:0] data_in181;
  wire [9:0] data_in181;
  input [9:0] data_in183;
  wire [9:0] data_in183;
  input [9:0] data_in185;
  wire [9:0] data_in185;
  input [9:0] data_in187;
  wire [9:0] data_in187;
  input [9:0] data_in189;
  wire [9:0] data_in189;
  input [9:0] data_in193;
  wire [9:0] data_in193;
  input [9:0] data_in195;
  wire [9:0] data_in195;
  input [9:0] data_in197;
  wire [9:0] data_in197;
  input [9:0] data_in199;
  wire [9:0] data_in199;
  input [9:0] data_in201;
  wire [9:0] data_in201;
  input [9:0] data_in203;
  wire [9:0] data_in203;
  input [9:0] data_in205;
  wire [9:0] data_in205;
  input [9:0] data_in207;
  wire [9:0] data_in207;
  input [9:0] data_in209;
  wire [9:0] data_in209;
  input [9:0] data_in211;
  wire [9:0] data_in211;
  input [9:0] data_in213;
  wire [9:0] data_in213;
  input [9:0] data_in215;
  wire [9:0] data_in215;
  input [9:0] data_in217;
  wire [9:0] data_in217;
  input [9:0] data_in219;
  wire [9:0] data_in219;
  input [9:0] data_in221;
  wire [9:0] data_in221;
  input [9:0] data_in225;
  wire [9:0] data_in225;
  input [9:0] data_in227;
  wire [9:0] data_in227;
  input [9:0] data_in229;
  wire [9:0] data_in229;
  input [9:0] data_in231;
  wire [9:0] data_in231;
  input [9:0] data_in233;
  wire [9:0] data_in233;
  input [9:0] data_in235;
  wire [9:0] data_in235;
  input [9:0] data_in237;
  wire [9:0] data_in237;
  input [9:0] data_in239;
  wire [9:0] data_in239;
  input [9:0] data_in241;
  wire [9:0] data_in241;
  input [9:0] data_in243;
  wire [9:0] data_in243;
  input [9:0] data_in245;
  wire [9:0] data_in245;
  input [9:0] data_in247;
  wire [9:0] data_in247;
  input [9:0] data_in249;
  wire [9:0] data_in249;
  input [9:0] data_in251;
  wire [9:0] data_in251;
  input [9:0] data_in253;
  wire [9:0] data_in253;
  input [9:0] data_in257;
  wire [9:0] data_in257;
  input [9:0] data_in259;
  wire [9:0] data_in259;
  input [9:0] data_in261;
  wire [9:0] data_in261;
  input [9:0] data_in263;
  wire [9:0] data_in263;
  input [9:0] data_in265;
  wire [9:0] data_in265;
  input [9:0] data_in267;
  wire [9:0] data_in267;
  input [9:0] data_in269;
  wire [9:0] data_in269;
  input [9:0] data_in271;
  wire [9:0] data_in271;
  input [9:0] data_in273;
  wire [9:0] data_in273;
  input [9:0] data_in275;
  wire [9:0] data_in275;
  input [9:0] data_in277;
  wire [9:0] data_in277;
  input [9:0] data_in279;
  wire [9:0] data_in279;
  input [9:0] data_in281;
  wire [9:0] data_in281;
  input [9:0] data_in283;
  wire [9:0] data_in283;
  input [9:0] data_in285;
  wire [9:0] data_in285;
  input [9:0] data_in289;
  wire [9:0] data_in289;
  input [9:0] data_in291;
  wire [9:0] data_in291;
  input [9:0] data_in293;
  wire [9:0] data_in293;
  input [9:0] data_in295;
  wire [9:0] data_in295;
  input [9:0] data_in297;
  wire [9:0] data_in297;
  input [9:0] data_in299;
  wire [9:0] data_in299;
  input [9:0] data_in301;
  wire [9:0] data_in301;
  input [9:0] data_in303;
  wire [9:0] data_in303;
  input [9:0] data_in305;
  wire [9:0] data_in305;
  input [9:0] data_in307;
  wire [9:0] data_in307;
  input [9:0] data_in309;
  wire [9:0] data_in309;
  input [9:0] data_in311;
  wire [9:0] data_in311;
  input [9:0] data_in313;
  wire [9:0] data_in313;
  input [9:0] data_in315;
  wire [9:0] data_in315;
  input [9:0] data_in317;
  wire [9:0] data_in317;
  input [9:0] data_in321;
  wire [9:0] data_in321;
  input [9:0] data_in323;
  wire [9:0] data_in323;
  input [9:0] data_in325;
  wire [9:0] data_in325;
  input [9:0] data_in327;
  wire [9:0] data_in327;
  input [9:0] data_in329;
  wire [9:0] data_in329;
  input [9:0] data_in331;
  wire [9:0] data_in331;
  input [9:0] data_in333;
  wire [9:0] data_in333;
  input [9:0] data_in335;
  wire [9:0] data_in335;
  input [9:0] data_in337;
  wire [9:0] data_in337;
  input [9:0] data_in339;
  wire [9:0] data_in339;
  input [9:0] data_in341;
  wire [9:0] data_in341;
  input [9:0] data_in343;
  wire [9:0] data_in343;
  input [9:0] data_in345;
  wire [9:0] data_in345;
  input [9:0] data_in347;
  wire [9:0] data_in347;
  input [9:0] data_in349;
  wire [9:0] data_in349;
  input [9:0] data_in353;
  wire [9:0] data_in353;
  input [9:0] data_in355;
  wire [9:0] data_in355;
  input [9:0] data_in357;
  wire [9:0] data_in357;
  input [9:0] data_in359;
  wire [9:0] data_in359;
  input [9:0] data_in361;
  wire [9:0] data_in361;
  input [9:0] data_in363;
  wire [9:0] data_in363;
  input [9:0] data_in365;
  wire [9:0] data_in365;
  input [9:0] data_in367;
  wire [9:0] data_in367;
  input [9:0] data_in369;
  wire [9:0] data_in369;
  input [9:0] data_in371;
  wire [9:0] data_in371;
  input [9:0] data_in373;
  wire [9:0] data_in373;
  input [9:0] data_in375;
  wire [9:0] data_in375;
  input [9:0] data_in377;
  wire [9:0] data_in377;
  input [9:0] data_in379;
  wire [9:0] data_in379;
  input [9:0] data_in381;
  wire [9:0] data_in381;
  input [9:0] data_in385;
  wire [9:0] data_in385;
  input [9:0] data_in387;
  wire [9:0] data_in387;
  input [9:0] data_in389;
  wire [9:0] data_in389;
  input [9:0] data_in391;
  wire [9:0] data_in391;
  input [9:0] data_in393;
  wire [9:0] data_in393;
  input [9:0] data_in395;
  wire [9:0] data_in395;
  input [9:0] data_in397;
  wire [9:0] data_in397;
  input [9:0] data_in399;
  wire [9:0] data_in399;
  input [9:0] data_in401;
  wire [9:0] data_in401;
  input [9:0] data_in403;
  wire [9:0] data_in403;
  input [9:0] data_in405;
  wire [9:0] data_in405;
  input [9:0] data_in407;
  wire [9:0] data_in407;
  input [9:0] data_in409;
  wire [9:0] data_in409;
  input [9:0] data_in411;
  wire [9:0] data_in411;
  input [9:0] data_in413;
  wire [9:0] data_in413;
  input [9:0] data_in417;
  wire [9:0] data_in417;
  input [9:0] data_in419;
  wire [9:0] data_in419;
  input [9:0] data_in421;
  wire [9:0] data_in421;
  input [9:0] data_in423;
  wire [9:0] data_in423;
  input [9:0] data_in425;
  wire [9:0] data_in425;
  input [9:0] data_in427;
  wire [9:0] data_in427;
  input [9:0] data_in429;
  wire [9:0] data_in429;
  input [9:0] data_in431;
  wire [9:0] data_in431;
  input [9:0] data_in433;
  wire [9:0] data_in433;
  input [9:0] data_in435;
  wire [9:0] data_in435;
  input [9:0] data_in437;
  wire [9:0] data_in437;
  input [9:0] data_in439;
  wire [9:0] data_in439;
  input [9:0] data_in441;
  wire [9:0] data_in441;
  input [9:0] data_in443;
  wire [9:0] data_in443;
  input [9:0] data_in445;
  wire [9:0] data_in445;
  input [9:0] data_in449;
  wire [9:0] data_in449;
  input [9:0] data_in451;
  wire [9:0] data_in451;
  input [9:0] data_in453;
  wire [9:0] data_in453;
  input [9:0] data_in455;
  wire [9:0] data_in455;
  input [9:0] data_in457;
  wire [9:0] data_in457;
  input [9:0] data_in459;
  wire [9:0] data_in459;
  input [9:0] data_in461;
  wire [9:0] data_in461;
  input [9:0] data_in463;
  wire [9:0] data_in463;
  input [9:0] data_in465;
  wire [9:0] data_in465;
  input [9:0] data_in467;
  wire [9:0] data_in467;
  input [9:0] data_in469;
  wire [9:0] data_in469;
  input [9:0] data_in471;
  wire [9:0] data_in471;
  input [9:0] data_in473;
  wire [9:0] data_in473;
  input [9:0] data_in475;
  wire [9:0] data_in475;
  input [9:0] data_in477;
  wire [9:0] data_in477;
  input [9:0] data_in_index33;
  wire [9:0] data_in_index33;
  input [9:0] data_in_index35;
  wire [9:0] data_in_index35;
  input [9:0] data_in_index37;
  wire [9:0] data_in_index37;
  input [9:0] data_in_index39;
  wire [9:0] data_in_index39;
  input [9:0] data_in_index41;
  wire [9:0] data_in_index41;
  input [9:0] data_in_index43;
  wire [9:0] data_in_index43;
  input [9:0] data_in_index45;
  wire [9:0] data_in_index45;
  input [9:0] data_in_index47;
  wire [9:0] data_in_index47;
  input [9:0] data_in_index49;
  wire [9:0] data_in_index49;
  input [9:0] data_in_index51;
  wire [9:0] data_in_index51;
  input [9:0] data_in_index53;
  wire [9:0] data_in_index53;
  input [9:0] data_in_index55;
  wire [9:0] data_in_index55;
  input [9:0] data_in_index57;
  wire [9:0] data_in_index57;
  input [9:0] data_in_index59;
  wire [9:0] data_in_index59;
  input [9:0] data_in_index61;
  wire [9:0] data_in_index61;
  input [9:0] data_in_index65;
  wire [9:0] data_in_index65;
  input [9:0] data_in_index67;
  wire [9:0] data_in_index67;
  input [9:0] data_in_index69;
  wire [9:0] data_in_index69;
  input [9:0] data_in_index71;
  wire [9:0] data_in_index71;
  input [9:0] data_in_index73;
  wire [9:0] data_in_index73;
  input [9:0] data_in_index75;
  wire [9:0] data_in_index75;
  input [9:0] data_in_index77;
  wire [9:0] data_in_index77;
  input [9:0] data_in_index79;
  wire [9:0] data_in_index79;
  input [9:0] data_in_index81;
  wire [9:0] data_in_index81;
  input [9:0] data_in_index83;
  wire [9:0] data_in_index83;
  input [9:0] data_in_index85;
  wire [9:0] data_in_index85;
  input [9:0] data_in_index87;
  wire [9:0] data_in_index87;
  input [9:0] data_in_index89;
  wire [9:0] data_in_index89;
  input [9:0] data_in_index91;
  wire [9:0] data_in_index91;
  input [9:0] data_in_index93;
  wire [9:0] data_in_index93;
  input [9:0] data_in_index97;
  wire [9:0] data_in_index97;
  input [9:0] data_in_index99;
  wire [9:0] data_in_index99;
  input [9:0] data_in_index101;
  wire [9:0] data_in_index101;
  input [9:0] data_in_index103;
  wire [9:0] data_in_index103;
  input [9:0] data_in_index105;
  wire [9:0] data_in_index105;
  input [9:0] data_in_index107;
  wire [9:0] data_in_index107;
  input [9:0] data_in_index109;
  wire [9:0] data_in_index109;
  input [9:0] data_in_index111;
  wire [9:0] data_in_index111;
  input [9:0] data_in_index113;
  wire [9:0] data_in_index113;
  input [9:0] data_in_index115;
  wire [9:0] data_in_index115;
  input [9:0] data_in_index117;
  wire [9:0] data_in_index117;
  input [9:0] data_in_index119;
  wire [9:0] data_in_index119;
  input [9:0] data_in_index121;
  wire [9:0] data_in_index121;
  input [9:0] data_in_index123;
  wire [9:0] data_in_index123;
  input [9:0] data_in_index125;
  wire [9:0] data_in_index125;
  input [9:0] data_in_index129;
  wire [9:0] data_in_index129;
  input [9:0] data_in_index131;
  wire [9:0] data_in_index131;
  input [9:0] data_in_index133;
  wire [9:0] data_in_index133;
  input [9:0] data_in_index135;
  wire [9:0] data_in_index135;
  input [9:0] data_in_index137;
  wire [9:0] data_in_index137;
  input [9:0] data_in_index139;
  wire [9:0] data_in_index139;
  input [9:0] data_in_index141;
  wire [9:0] data_in_index141;
  input [9:0] data_in_index143;
  wire [9:0] data_in_index143;
  input [9:0] data_in_index145;
  wire [9:0] data_in_index145;
  input [9:0] data_in_index147;
  wire [9:0] data_in_index147;
  input [9:0] data_in_index149;
  wire [9:0] data_in_index149;
  input [9:0] data_in_index151;
  wire [9:0] data_in_index151;
  input [9:0] data_in_index153;
  wire [9:0] data_in_index153;
  input [9:0] data_in_index155;
  wire [9:0] data_in_index155;
  input [9:0] data_in_index157;
  wire [9:0] data_in_index157;
  input [9:0] data_in_index161;
  wire [9:0] data_in_index161;
  input [9:0] data_in_index163;
  wire [9:0] data_in_index163;
  input [9:0] data_in_index165;
  wire [9:0] data_in_index165;
  input [9:0] data_in_index167;
  wire [9:0] data_in_index167;
  input [9:0] data_in_index169;
  wire [9:0] data_in_index169;
  input [9:0] data_in_index171;
  wire [9:0] data_in_index171;
  input [9:0] data_in_index173;
  wire [9:0] data_in_index173;
  input [9:0] data_in_index175;
  wire [9:0] data_in_index175;
  input [9:0] data_in_index177;
  wire [9:0] data_in_index177;
  input [9:0] data_in_index179;
  wire [9:0] data_in_index179;
  input [9:0] data_in_index181;
  wire [9:0] data_in_index181;
  input [9:0] data_in_index183;
  wire [9:0] data_in_index183;
  input [9:0] data_in_index185;
  wire [9:0] data_in_index185;
  input [9:0] data_in_index187;
  wire [9:0] data_in_index187;
  input [9:0] data_in_index189;
  wire [9:0] data_in_index189;
  input [9:0] data_in_index193;
  wire [9:0] data_in_index193;
  input [9:0] data_in_index195;
  wire [9:0] data_in_index195;
  input [9:0] data_in_index197;
  wire [9:0] data_in_index197;
  input [9:0] data_in_index199;
  wire [9:0] data_in_index199;
  input [9:0] data_in_index201;
  wire [9:0] data_in_index201;
  input [9:0] data_in_index203;
  wire [9:0] data_in_index203;
  input [9:0] data_in_index205;
  wire [9:0] data_in_index205;
  input [9:0] data_in_index207;
  wire [9:0] data_in_index207;
  input [9:0] data_in_index209;
  wire [9:0] data_in_index209;
  input [9:0] data_in_index211;
  wire [9:0] data_in_index211;
  input [9:0] data_in_index213;
  wire [9:0] data_in_index213;
  input [9:0] data_in_index215;
  wire [9:0] data_in_index215;
  input [9:0] data_in_index217;
  wire [9:0] data_in_index217;
  input [9:0] data_in_index219;
  wire [9:0] data_in_index219;
  input [9:0] data_in_index221;
  wire [9:0] data_in_index221;
  input [9:0] data_in_index225;
  wire [9:0] data_in_index225;
  input [9:0] data_in_index227;
  wire [9:0] data_in_index227;
  input [9:0] data_in_index229;
  wire [9:0] data_in_index229;
  input [9:0] data_in_index231;
  wire [9:0] data_in_index231;
  input [9:0] data_in_index233;
  wire [9:0] data_in_index233;
  input [9:0] data_in_index235;
  wire [9:0] data_in_index235;
  input [9:0] data_in_index237;
  wire [9:0] data_in_index237;
  input [9:0] data_in_index239;
  wire [9:0] data_in_index239;
  input [9:0] data_in_index241;
  wire [9:0] data_in_index241;
  input [9:0] data_in_index243;
  wire [9:0] data_in_index243;
  input [9:0] data_in_index245;
  wire [9:0] data_in_index245;
  input [9:0] data_in_index247;
  wire [9:0] data_in_index247;
  input [9:0] data_in_index249;
  wire [9:0] data_in_index249;
  input [9:0] data_in_index251;
  wire [9:0] data_in_index251;
  input [9:0] data_in_index253;
  wire [9:0] data_in_index253;
  input [9:0] data_in_index257;
  wire [9:0] data_in_index257;
  input [9:0] data_in_index259;
  wire [9:0] data_in_index259;
  input [9:0] data_in_index261;
  wire [9:0] data_in_index261;
  input [9:0] data_in_index263;
  wire [9:0] data_in_index263;
  input [9:0] data_in_index265;
  wire [9:0] data_in_index265;
  input [9:0] data_in_index267;
  wire [9:0] data_in_index267;
  input [9:0] data_in_index269;
  wire [9:0] data_in_index269;
  input [9:0] data_in_index271;
  wire [9:0] data_in_index271;
  input [9:0] data_in_index273;
  wire [9:0] data_in_index273;
  input [9:0] data_in_index275;
  wire [9:0] data_in_index275;
  input [9:0] data_in_index277;
  wire [9:0] data_in_index277;
  input [9:0] data_in_index279;
  wire [9:0] data_in_index279;
  input [9:0] data_in_index281;
  wire [9:0] data_in_index281;
  input [9:0] data_in_index283;
  wire [9:0] data_in_index283;
  input [9:0] data_in_index285;
  wire [9:0] data_in_index285;
  input [9:0] data_in_index289;
  wire [9:0] data_in_index289;
  input [9:0] data_in_index291;
  wire [9:0] data_in_index291;
  input [9:0] data_in_index293;
  wire [9:0] data_in_index293;
  input [9:0] data_in_index295;
  wire [9:0] data_in_index295;
  input [9:0] data_in_index297;
  wire [9:0] data_in_index297;
  input [9:0] data_in_index299;
  wire [9:0] data_in_index299;
  input [9:0] data_in_index301;
  wire [9:0] data_in_index301;
  input [9:0] data_in_index303;
  wire [9:0] data_in_index303;
  input [9:0] data_in_index305;
  wire [9:0] data_in_index305;
  input [9:0] data_in_index307;
  wire [9:0] data_in_index307;
  input [9:0] data_in_index309;
  wire [9:0] data_in_index309;
  input [9:0] data_in_index311;
  wire [9:0] data_in_index311;
  input [9:0] data_in_index313;
  wire [9:0] data_in_index313;
  input [9:0] data_in_index315;
  wire [9:0] data_in_index315;
  input [9:0] data_in_index317;
  wire [9:0] data_in_index317;
  input [9:0] data_in_index321;
  wire [9:0] data_in_index321;
  input [9:0] data_in_index323;
  wire [9:0] data_in_index323;
  input [9:0] data_in_index325;
  wire [9:0] data_in_index325;
  input [9:0] data_in_index327;
  wire [9:0] data_in_index327;
  input [9:0] data_in_index329;
  wire [9:0] data_in_index329;
  input [9:0] data_in_index331;
  wire [9:0] data_in_index331;
  input [9:0] data_in_index333;
  wire [9:0] data_in_index333;
  input [9:0] data_in_index335;
  wire [9:0] data_in_index335;
  input [9:0] data_in_index337;
  wire [9:0] data_in_index337;
  input [9:0] data_in_index339;
  wire [9:0] data_in_index339;
  input [9:0] data_in_index341;
  wire [9:0] data_in_index341;
  input [9:0] data_in_index343;
  wire [9:0] data_in_index343;
  input [9:0] data_in_index345;
  wire [9:0] data_in_index345;
  input [9:0] data_in_index347;
  wire [9:0] data_in_index347;
  input [9:0] data_in_index349;
  wire [9:0] data_in_index349;
  input [9:0] data_in_index353;
  wire [9:0] data_in_index353;
  input [9:0] data_in_index355;
  wire [9:0] data_in_index355;
  input [9:0] data_in_index357;
  wire [9:0] data_in_index357;
  input [9:0] data_in_index359;
  wire [9:0] data_in_index359;
  input [9:0] data_in_index361;
  wire [9:0] data_in_index361;
  input [9:0] data_in_index363;
  wire [9:0] data_in_index363;
  input [9:0] data_in_index365;
  wire [9:0] data_in_index365;
  input [9:0] data_in_index367;
  wire [9:0] data_in_index367;
  input [9:0] data_in_index369;
  wire [9:0] data_in_index369;
  input [9:0] data_in_index371;
  wire [9:0] data_in_index371;
  input [9:0] data_in_index373;
  wire [9:0] data_in_index373;
  input [9:0] data_in_index375;
  wire [9:0] data_in_index375;
  input [9:0] data_in_index377;
  wire [9:0] data_in_index377;
  input [9:0] data_in_index379;
  wire [9:0] data_in_index379;
  input [9:0] data_in_index381;
  wire [9:0] data_in_index381;
  input [9:0] data_in_index385;
  wire [9:0] data_in_index385;
  input [9:0] data_in_index387;
  wire [9:0] data_in_index387;
  input [9:0] data_in_index389;
  wire [9:0] data_in_index389;
  input [9:0] data_in_index391;
  wire [9:0] data_in_index391;
  input [9:0] data_in_index393;
  wire [9:0] data_in_index393;
  input [9:0] data_in_index395;
  wire [9:0] data_in_index395;
  input [9:0] data_in_index397;
  wire [9:0] data_in_index397;
  input [9:0] data_in_index399;
  wire [9:0] data_in_index399;
  input [9:0] data_in_index401;
  wire [9:0] data_in_index401;
  input [9:0] data_in_index403;
  wire [9:0] data_in_index403;
  input [9:0] data_in_index405;
  wire [9:0] data_in_index405;
  input [9:0] data_in_index407;
  wire [9:0] data_in_index407;
  input [9:0] data_in_index409;
  wire [9:0] data_in_index409;
  input [9:0] data_in_index411;
  wire [9:0] data_in_index411;
  input [9:0] data_in_index413;
  wire [9:0] data_in_index413;
  input [9:0] data_in_index417;
  wire [9:0] data_in_index417;
  input [9:0] data_in_index419;
  wire [9:0] data_in_index419;
  input [9:0] data_in_index421;
  wire [9:0] data_in_index421;
  input [9:0] data_in_index423;
  wire [9:0] data_in_index423;
  input [9:0] data_in_index425;
  wire [9:0] data_in_index425;
  input [9:0] data_in_index427;
  wire [9:0] data_in_index427;
  input [9:0] data_in_index429;
  wire [9:0] data_in_index429;
  input [9:0] data_in_index431;
  wire [9:0] data_in_index431;
  input [9:0] data_in_index433;
  wire [9:0] data_in_index433;
  input [9:0] data_in_index435;
  wire [9:0] data_in_index435;
  input [9:0] data_in_index437;
  wire [9:0] data_in_index437;
  input [9:0] data_in_index439;
  wire [9:0] data_in_index439;
  input [9:0] data_in_index441;
  wire [9:0] data_in_index441;
  input [9:0] data_in_index443;
  wire [9:0] data_in_index443;
  input [9:0] data_in_index445;
  wire [9:0] data_in_index445;
  input [9:0] data_in_index449;
  wire [9:0] data_in_index449;
  input [9:0] data_in_index451;
  wire [9:0] data_in_index451;
  input [9:0] data_in_index453;
  wire [9:0] data_in_index453;
  input [9:0] data_in_index455;
  wire [9:0] data_in_index455;
  input [9:0] data_in_index457;
  wire [9:0] data_in_index457;
  input [9:0] data_in_index459;
  wire [9:0] data_in_index459;
  input [9:0] data_in_index461;
  wire [9:0] data_in_index461;
  input [9:0] data_in_index463;
  wire [9:0] data_in_index463;
  input [9:0] data_in_index465;
  wire [9:0] data_in_index465;
  input [9:0] data_in_index467;
  wire [9:0] data_in_index467;
  input [9:0] data_in_index469;
  wire [9:0] data_in_index469;
  input [9:0] data_in_index471;
  wire [9:0] data_in_index471;
  input [9:0] data_in_index473;
  wire [9:0] data_in_index473;
  input [9:0] data_in_index475;
  wire [9:0] data_in_index475;
  input [9:0] data_in_index477;
  wire [9:0] data_in_index477;
  output [9:0] sub_array_out;
  wire [9:0] sub_array_out;
  input subs_exe;
  wire subs_exe;
  reg [9:0] sub_reg;
  wire [9:0] _sub_plot_x_hikareru;
  wire [9:0] _sub_plot_x_moto;
  wire [9:0] _sub_plot_x_sa;
  wire _sub_plot_x_in_do;
  wire _sub_plot_x_p_reset;
  wire _sub_plot_x_m_clock;
  wire [9:0] _sub_plot_x_209_hikareru;
  wire [9:0] _sub_plot_x_209_moto;
  wire [9:0] _sub_plot_x_209_sa;
  wire _sub_plot_x_209_in_do;
  wire _sub_plot_x_209_p_reset;
  wire _sub_plot_x_209_m_clock;
  wire [9:0] _sub_plot_x_208_hikareru;
  wire [9:0] _sub_plot_x_208_moto;
  wire [9:0] _sub_plot_x_208_sa;
  wire _sub_plot_x_208_in_do;
  wire _sub_plot_x_208_p_reset;
  wire _sub_plot_x_208_m_clock;
  wire [9:0] _sub_plot_x_207_hikareru;
  wire [9:0] _sub_plot_x_207_moto;
  wire [9:0] _sub_plot_x_207_sa;
  wire _sub_plot_x_207_in_do;
  wire _sub_plot_x_207_p_reset;
  wire _sub_plot_x_207_m_clock;
  wire [9:0] _sub_plot_x_206_hikareru;
  wire [9:0] _sub_plot_x_206_moto;
  wire [9:0] _sub_plot_x_206_sa;
  wire _sub_plot_x_206_in_do;
  wire _sub_plot_x_206_p_reset;
  wire _sub_plot_x_206_m_clock;
  wire [9:0] _sub_plot_x_205_hikareru;
  wire [9:0] _sub_plot_x_205_moto;
  wire [9:0] _sub_plot_x_205_sa;
  wire _sub_plot_x_205_in_do;
  wire _sub_plot_x_205_p_reset;
  wire _sub_plot_x_205_m_clock;
  wire [9:0] _sub_plot_x_204_hikareru;
  wire [9:0] _sub_plot_x_204_moto;
  wire [9:0] _sub_plot_x_204_sa;
  wire _sub_plot_x_204_in_do;
  wire _sub_plot_x_204_p_reset;
  wire _sub_plot_x_204_m_clock;
  wire [9:0] _sub_plot_x_203_hikareru;
  wire [9:0] _sub_plot_x_203_moto;
  wire [9:0] _sub_plot_x_203_sa;
  wire _sub_plot_x_203_in_do;
  wire _sub_plot_x_203_p_reset;
  wire _sub_plot_x_203_m_clock;
  wire [9:0] _sub_plot_x_202_hikareru;
  wire [9:0] _sub_plot_x_202_moto;
  wire [9:0] _sub_plot_x_202_sa;
  wire _sub_plot_x_202_in_do;
  wire _sub_plot_x_202_p_reset;
  wire _sub_plot_x_202_m_clock;
  wire [9:0] _sub_plot_x_201_hikareru;
  wire [9:0] _sub_plot_x_201_moto;
  wire [9:0] _sub_plot_x_201_sa;
  wire _sub_plot_x_201_in_do;
  wire _sub_plot_x_201_p_reset;
  wire _sub_plot_x_201_m_clock;
  wire [9:0] _sub_plot_x_200_hikareru;
  wire [9:0] _sub_plot_x_200_moto;
  wire [9:0] _sub_plot_x_200_sa;
  wire _sub_plot_x_200_in_do;
  wire _sub_plot_x_200_p_reset;
  wire _sub_plot_x_200_m_clock;
  wire [9:0] _sub_plot_x_199_hikareru;
  wire [9:0] _sub_plot_x_199_moto;
  wire [9:0] _sub_plot_x_199_sa;
  wire _sub_plot_x_199_in_do;
  wire _sub_plot_x_199_p_reset;
  wire _sub_plot_x_199_m_clock;
  wire [9:0] _sub_plot_x_198_hikareru;
  wire [9:0] _sub_plot_x_198_moto;
  wire [9:0] _sub_plot_x_198_sa;
  wire _sub_plot_x_198_in_do;
  wire _sub_plot_x_198_p_reset;
  wire _sub_plot_x_198_m_clock;
  wire [9:0] _sub_plot_x_197_hikareru;
  wire [9:0] _sub_plot_x_197_moto;
  wire [9:0] _sub_plot_x_197_sa;
  wire _sub_plot_x_197_in_do;
  wire _sub_plot_x_197_p_reset;
  wire _sub_plot_x_197_m_clock;
  wire [9:0] _sub_plot_x_196_hikareru;
  wire [9:0] _sub_plot_x_196_moto;
  wire [9:0] _sub_plot_x_196_sa;
  wire _sub_plot_x_196_in_do;
  wire _sub_plot_x_196_p_reset;
  wire _sub_plot_x_196_m_clock;
  wire [9:0] _sub_plot_x_195_hikareru;
  wire [9:0] _sub_plot_x_195_moto;
  wire [9:0] _sub_plot_x_195_sa;
  wire _sub_plot_x_195_in_do;
  wire _sub_plot_x_195_p_reset;
  wire _sub_plot_x_195_m_clock;
  wire [9:0] _sub_plot_x_194_hikareru;
  wire [9:0] _sub_plot_x_194_moto;
  wire [9:0] _sub_plot_x_194_sa;
  wire _sub_plot_x_194_in_do;
  wire _sub_plot_x_194_p_reset;
  wire _sub_plot_x_194_m_clock;
  wire [9:0] _sub_plot_x_193_hikareru;
  wire [9:0] _sub_plot_x_193_moto;
  wire [9:0] _sub_plot_x_193_sa;
  wire _sub_plot_x_193_in_do;
  wire _sub_plot_x_193_p_reset;
  wire _sub_plot_x_193_m_clock;
  wire [9:0] _sub_plot_x_192_hikareru;
  wire [9:0] _sub_plot_x_192_moto;
  wire [9:0] _sub_plot_x_192_sa;
  wire _sub_plot_x_192_in_do;
  wire _sub_plot_x_192_p_reset;
  wire _sub_plot_x_192_m_clock;
  wire [9:0] _sub_plot_x_191_hikareru;
  wire [9:0] _sub_plot_x_191_moto;
  wire [9:0] _sub_plot_x_191_sa;
  wire _sub_plot_x_191_in_do;
  wire _sub_plot_x_191_p_reset;
  wire _sub_plot_x_191_m_clock;
  wire [9:0] _sub_plot_x_190_hikareru;
  wire [9:0] _sub_plot_x_190_moto;
  wire [9:0] _sub_plot_x_190_sa;
  wire _sub_plot_x_190_in_do;
  wire _sub_plot_x_190_p_reset;
  wire _sub_plot_x_190_m_clock;
  wire [9:0] _sub_plot_x_189_hikareru;
  wire [9:0] _sub_plot_x_189_moto;
  wire [9:0] _sub_plot_x_189_sa;
  wire _sub_plot_x_189_in_do;
  wire _sub_plot_x_189_p_reset;
  wire _sub_plot_x_189_m_clock;
  wire [9:0] _sub_plot_x_188_hikareru;
  wire [9:0] _sub_plot_x_188_moto;
  wire [9:0] _sub_plot_x_188_sa;
  wire _sub_plot_x_188_in_do;
  wire _sub_plot_x_188_p_reset;
  wire _sub_plot_x_188_m_clock;
  wire [9:0] _sub_plot_x_187_hikareru;
  wire [9:0] _sub_plot_x_187_moto;
  wire [9:0] _sub_plot_x_187_sa;
  wire _sub_plot_x_187_in_do;
  wire _sub_plot_x_187_p_reset;
  wire _sub_plot_x_187_m_clock;
  wire [9:0] _sub_plot_x_186_hikareru;
  wire [9:0] _sub_plot_x_186_moto;
  wire [9:0] _sub_plot_x_186_sa;
  wire _sub_plot_x_186_in_do;
  wire _sub_plot_x_186_p_reset;
  wire _sub_plot_x_186_m_clock;
  wire [9:0] _sub_plot_x_185_hikareru;
  wire [9:0] _sub_plot_x_185_moto;
  wire [9:0] _sub_plot_x_185_sa;
  wire _sub_plot_x_185_in_do;
  wire _sub_plot_x_185_p_reset;
  wire _sub_plot_x_185_m_clock;
  wire [9:0] _sub_plot_x_184_hikareru;
  wire [9:0] _sub_plot_x_184_moto;
  wire [9:0] _sub_plot_x_184_sa;
  wire _sub_plot_x_184_in_do;
  wire _sub_plot_x_184_p_reset;
  wire _sub_plot_x_184_m_clock;
  wire [9:0] _sub_plot_x_183_hikareru;
  wire [9:0] _sub_plot_x_183_moto;
  wire [9:0] _sub_plot_x_183_sa;
  wire _sub_plot_x_183_in_do;
  wire _sub_plot_x_183_p_reset;
  wire _sub_plot_x_183_m_clock;
  wire [9:0] _sub_plot_x_182_hikareru;
  wire [9:0] _sub_plot_x_182_moto;
  wire [9:0] _sub_plot_x_182_sa;
  wire _sub_plot_x_182_in_do;
  wire _sub_plot_x_182_p_reset;
  wire _sub_plot_x_182_m_clock;
  wire [9:0] _sub_plot_x_181_hikareru;
  wire [9:0] _sub_plot_x_181_moto;
  wire [9:0] _sub_plot_x_181_sa;
  wire _sub_plot_x_181_in_do;
  wire _sub_plot_x_181_p_reset;
  wire _sub_plot_x_181_m_clock;
  wire [9:0] _sub_plot_x_180_hikareru;
  wire [9:0] _sub_plot_x_180_moto;
  wire [9:0] _sub_plot_x_180_sa;
  wire _sub_plot_x_180_in_do;
  wire _sub_plot_x_180_p_reset;
  wire _sub_plot_x_180_m_clock;
  wire [9:0] _sub_plot_x_179_hikareru;
  wire [9:0] _sub_plot_x_179_moto;
  wire [9:0] _sub_plot_x_179_sa;
  wire _sub_plot_x_179_in_do;
  wire _sub_plot_x_179_p_reset;
  wire _sub_plot_x_179_m_clock;
  wire [9:0] _sub_plot_x_178_hikareru;
  wire [9:0] _sub_plot_x_178_moto;
  wire [9:0] _sub_plot_x_178_sa;
  wire _sub_plot_x_178_in_do;
  wire _sub_plot_x_178_p_reset;
  wire _sub_plot_x_178_m_clock;
  wire [9:0] _sub_plot_x_177_hikareru;
  wire [9:0] _sub_plot_x_177_moto;
  wire [9:0] _sub_plot_x_177_sa;
  wire _sub_plot_x_177_in_do;
  wire _sub_plot_x_177_p_reset;
  wire _sub_plot_x_177_m_clock;
  wire [9:0] _sub_plot_x_176_hikareru;
  wire [9:0] _sub_plot_x_176_moto;
  wire [9:0] _sub_plot_x_176_sa;
  wire _sub_plot_x_176_in_do;
  wire _sub_plot_x_176_p_reset;
  wire _sub_plot_x_176_m_clock;
  wire [9:0] _sub_plot_x_175_hikareru;
  wire [9:0] _sub_plot_x_175_moto;
  wire [9:0] _sub_plot_x_175_sa;
  wire _sub_plot_x_175_in_do;
  wire _sub_plot_x_175_p_reset;
  wire _sub_plot_x_175_m_clock;
  wire [9:0] _sub_plot_x_174_hikareru;
  wire [9:0] _sub_plot_x_174_moto;
  wire [9:0] _sub_plot_x_174_sa;
  wire _sub_plot_x_174_in_do;
  wire _sub_plot_x_174_p_reset;
  wire _sub_plot_x_174_m_clock;
  wire [9:0] _sub_plot_x_173_hikareru;
  wire [9:0] _sub_plot_x_173_moto;
  wire [9:0] _sub_plot_x_173_sa;
  wire _sub_plot_x_173_in_do;
  wire _sub_plot_x_173_p_reset;
  wire _sub_plot_x_173_m_clock;
  wire [9:0] _sub_plot_x_172_hikareru;
  wire [9:0] _sub_plot_x_172_moto;
  wire [9:0] _sub_plot_x_172_sa;
  wire _sub_plot_x_172_in_do;
  wire _sub_plot_x_172_p_reset;
  wire _sub_plot_x_172_m_clock;
  wire [9:0] _sub_plot_x_171_hikareru;
  wire [9:0] _sub_plot_x_171_moto;
  wire [9:0] _sub_plot_x_171_sa;
  wire _sub_plot_x_171_in_do;
  wire _sub_plot_x_171_p_reset;
  wire _sub_plot_x_171_m_clock;
  wire [9:0] _sub_plot_x_170_hikareru;
  wire [9:0] _sub_plot_x_170_moto;
  wire [9:0] _sub_plot_x_170_sa;
  wire _sub_plot_x_170_in_do;
  wire _sub_plot_x_170_p_reset;
  wire _sub_plot_x_170_m_clock;
  wire [9:0] _sub_plot_x_169_hikareru;
  wire [9:0] _sub_plot_x_169_moto;
  wire [9:0] _sub_plot_x_169_sa;
  wire _sub_plot_x_169_in_do;
  wire _sub_plot_x_169_p_reset;
  wire _sub_plot_x_169_m_clock;
  wire [9:0] _sub_plot_x_168_hikareru;
  wire [9:0] _sub_plot_x_168_moto;
  wire [9:0] _sub_plot_x_168_sa;
  wire _sub_plot_x_168_in_do;
  wire _sub_plot_x_168_p_reset;
  wire _sub_plot_x_168_m_clock;
  wire [9:0] _sub_plot_x_167_hikareru;
  wire [9:0] _sub_plot_x_167_moto;
  wire [9:0] _sub_plot_x_167_sa;
  wire _sub_plot_x_167_in_do;
  wire _sub_plot_x_167_p_reset;
  wire _sub_plot_x_167_m_clock;
  wire [9:0] _sub_plot_x_166_hikareru;
  wire [9:0] _sub_plot_x_166_moto;
  wire [9:0] _sub_plot_x_166_sa;
  wire _sub_plot_x_166_in_do;
  wire _sub_plot_x_166_p_reset;
  wire _sub_plot_x_166_m_clock;
  wire [9:0] _sub_plot_x_165_hikareru;
  wire [9:0] _sub_plot_x_165_moto;
  wire [9:0] _sub_plot_x_165_sa;
  wire _sub_plot_x_165_in_do;
  wire _sub_plot_x_165_p_reset;
  wire _sub_plot_x_165_m_clock;
  wire [9:0] _sub_plot_x_164_hikareru;
  wire [9:0] _sub_plot_x_164_moto;
  wire [9:0] _sub_plot_x_164_sa;
  wire _sub_plot_x_164_in_do;
  wire _sub_plot_x_164_p_reset;
  wire _sub_plot_x_164_m_clock;
  wire [9:0] _sub_plot_x_163_hikareru;
  wire [9:0] _sub_plot_x_163_moto;
  wire [9:0] _sub_plot_x_163_sa;
  wire _sub_plot_x_163_in_do;
  wire _sub_plot_x_163_p_reset;
  wire _sub_plot_x_163_m_clock;
  wire [9:0] _sub_plot_x_162_hikareru;
  wire [9:0] _sub_plot_x_162_moto;
  wire [9:0] _sub_plot_x_162_sa;
  wire _sub_plot_x_162_in_do;
  wire _sub_plot_x_162_p_reset;
  wire _sub_plot_x_162_m_clock;
  wire [9:0] _sub_plot_x_161_hikareru;
  wire [9:0] _sub_plot_x_161_moto;
  wire [9:0] _sub_plot_x_161_sa;
  wire _sub_plot_x_161_in_do;
  wire _sub_plot_x_161_p_reset;
  wire _sub_plot_x_161_m_clock;
  wire [9:0] _sub_plot_x_160_hikareru;
  wire [9:0] _sub_plot_x_160_moto;
  wire [9:0] _sub_plot_x_160_sa;
  wire _sub_plot_x_160_in_do;
  wire _sub_plot_x_160_p_reset;
  wire _sub_plot_x_160_m_clock;
  wire [9:0] _sub_plot_x_159_hikareru;
  wire [9:0] _sub_plot_x_159_moto;
  wire [9:0] _sub_plot_x_159_sa;
  wire _sub_plot_x_159_in_do;
  wire _sub_plot_x_159_p_reset;
  wire _sub_plot_x_159_m_clock;
  wire [9:0] _sub_plot_x_158_hikareru;
  wire [9:0] _sub_plot_x_158_moto;
  wire [9:0] _sub_plot_x_158_sa;
  wire _sub_plot_x_158_in_do;
  wire _sub_plot_x_158_p_reset;
  wire _sub_plot_x_158_m_clock;
  wire [9:0] _sub_plot_x_157_hikareru;
  wire [9:0] _sub_plot_x_157_moto;
  wire [9:0] _sub_plot_x_157_sa;
  wire _sub_plot_x_157_in_do;
  wire _sub_plot_x_157_p_reset;
  wire _sub_plot_x_157_m_clock;
  wire [9:0] _sub_plot_x_156_hikareru;
  wire [9:0] _sub_plot_x_156_moto;
  wire [9:0] _sub_plot_x_156_sa;
  wire _sub_plot_x_156_in_do;
  wire _sub_plot_x_156_p_reset;
  wire _sub_plot_x_156_m_clock;
  wire [9:0] _sub_plot_x_155_hikareru;
  wire [9:0] _sub_plot_x_155_moto;
  wire [9:0] _sub_plot_x_155_sa;
  wire _sub_plot_x_155_in_do;
  wire _sub_plot_x_155_p_reset;
  wire _sub_plot_x_155_m_clock;
  wire [9:0] _sub_plot_x_154_hikareru;
  wire [9:0] _sub_plot_x_154_moto;
  wire [9:0] _sub_plot_x_154_sa;
  wire _sub_plot_x_154_in_do;
  wire _sub_plot_x_154_p_reset;
  wire _sub_plot_x_154_m_clock;
  wire [9:0] _sub_plot_x_153_hikareru;
  wire [9:0] _sub_plot_x_153_moto;
  wire [9:0] _sub_plot_x_153_sa;
  wire _sub_plot_x_153_in_do;
  wire _sub_plot_x_153_p_reset;
  wire _sub_plot_x_153_m_clock;
  wire [9:0] _sub_plot_x_152_hikareru;
  wire [9:0] _sub_plot_x_152_moto;
  wire [9:0] _sub_plot_x_152_sa;
  wire _sub_plot_x_152_in_do;
  wire _sub_plot_x_152_p_reset;
  wire _sub_plot_x_152_m_clock;
  wire [9:0] _sub_plot_x_151_hikareru;
  wire [9:0] _sub_plot_x_151_moto;
  wire [9:0] _sub_plot_x_151_sa;
  wire _sub_plot_x_151_in_do;
  wire _sub_plot_x_151_p_reset;
  wire _sub_plot_x_151_m_clock;
  wire [9:0] _sub_plot_x_150_hikareru;
  wire [9:0] _sub_plot_x_150_moto;
  wire [9:0] _sub_plot_x_150_sa;
  wire _sub_plot_x_150_in_do;
  wire _sub_plot_x_150_p_reset;
  wire _sub_plot_x_150_m_clock;
  wire [9:0] _sub_plot_x_149_hikareru;
  wire [9:0] _sub_plot_x_149_moto;
  wire [9:0] _sub_plot_x_149_sa;
  wire _sub_plot_x_149_in_do;
  wire _sub_plot_x_149_p_reset;
  wire _sub_plot_x_149_m_clock;
  wire [9:0] _sub_plot_x_148_hikareru;
  wire [9:0] _sub_plot_x_148_moto;
  wire [9:0] _sub_plot_x_148_sa;
  wire _sub_plot_x_148_in_do;
  wire _sub_plot_x_148_p_reset;
  wire _sub_plot_x_148_m_clock;
  wire [9:0] _sub_plot_x_147_hikareru;
  wire [9:0] _sub_plot_x_147_moto;
  wire [9:0] _sub_plot_x_147_sa;
  wire _sub_plot_x_147_in_do;
  wire _sub_plot_x_147_p_reset;
  wire _sub_plot_x_147_m_clock;
  wire [9:0] _sub_plot_x_146_hikareru;
  wire [9:0] _sub_plot_x_146_moto;
  wire [9:0] _sub_plot_x_146_sa;
  wire _sub_plot_x_146_in_do;
  wire _sub_plot_x_146_p_reset;
  wire _sub_plot_x_146_m_clock;
  wire [9:0] _sub_plot_x_145_hikareru;
  wire [9:0] _sub_plot_x_145_moto;
  wire [9:0] _sub_plot_x_145_sa;
  wire _sub_plot_x_145_in_do;
  wire _sub_plot_x_145_p_reset;
  wire _sub_plot_x_145_m_clock;
  wire [9:0] _sub_plot_x_144_hikareru;
  wire [9:0] _sub_plot_x_144_moto;
  wire [9:0] _sub_plot_x_144_sa;
  wire _sub_plot_x_144_in_do;
  wire _sub_plot_x_144_p_reset;
  wire _sub_plot_x_144_m_clock;
  wire [9:0] _sub_plot_x_143_hikareru;
  wire [9:0] _sub_plot_x_143_moto;
  wire [9:0] _sub_plot_x_143_sa;
  wire _sub_plot_x_143_in_do;
  wire _sub_plot_x_143_p_reset;
  wire _sub_plot_x_143_m_clock;
  wire [9:0] _sub_plot_x_142_hikareru;
  wire [9:0] _sub_plot_x_142_moto;
  wire [9:0] _sub_plot_x_142_sa;
  wire _sub_plot_x_142_in_do;
  wire _sub_plot_x_142_p_reset;
  wire _sub_plot_x_142_m_clock;
  wire [9:0] _sub_plot_x_141_hikareru;
  wire [9:0] _sub_plot_x_141_moto;
  wire [9:0] _sub_plot_x_141_sa;
  wire _sub_plot_x_141_in_do;
  wire _sub_plot_x_141_p_reset;
  wire _sub_plot_x_141_m_clock;
  wire [9:0] _sub_plot_x_140_hikareru;
  wire [9:0] _sub_plot_x_140_moto;
  wire [9:0] _sub_plot_x_140_sa;
  wire _sub_plot_x_140_in_do;
  wire _sub_plot_x_140_p_reset;
  wire _sub_plot_x_140_m_clock;
  wire [9:0] _sub_plot_x_139_hikareru;
  wire [9:0] _sub_plot_x_139_moto;
  wire [9:0] _sub_plot_x_139_sa;
  wire _sub_plot_x_139_in_do;
  wire _sub_plot_x_139_p_reset;
  wire _sub_plot_x_139_m_clock;
  wire [9:0] _sub_plot_x_138_hikareru;
  wire [9:0] _sub_plot_x_138_moto;
  wire [9:0] _sub_plot_x_138_sa;
  wire _sub_plot_x_138_in_do;
  wire _sub_plot_x_138_p_reset;
  wire _sub_plot_x_138_m_clock;
  wire [9:0] _sub_plot_x_137_hikareru;
  wire [9:0] _sub_plot_x_137_moto;
  wire [9:0] _sub_plot_x_137_sa;
  wire _sub_plot_x_137_in_do;
  wire _sub_plot_x_137_p_reset;
  wire _sub_plot_x_137_m_clock;
  wire [9:0] _sub_plot_x_136_hikareru;
  wire [9:0] _sub_plot_x_136_moto;
  wire [9:0] _sub_plot_x_136_sa;
  wire _sub_plot_x_136_in_do;
  wire _sub_plot_x_136_p_reset;
  wire _sub_plot_x_136_m_clock;
  wire [9:0] _sub_plot_x_135_hikareru;
  wire [9:0] _sub_plot_x_135_moto;
  wire [9:0] _sub_plot_x_135_sa;
  wire _sub_plot_x_135_in_do;
  wire _sub_plot_x_135_p_reset;
  wire _sub_plot_x_135_m_clock;
  wire [9:0] _sub_plot_x_134_hikareru;
  wire [9:0] _sub_plot_x_134_moto;
  wire [9:0] _sub_plot_x_134_sa;
  wire _sub_plot_x_134_in_do;
  wire _sub_plot_x_134_p_reset;
  wire _sub_plot_x_134_m_clock;
  wire [9:0] _sub_plot_x_133_hikareru;
  wire [9:0] _sub_plot_x_133_moto;
  wire [9:0] _sub_plot_x_133_sa;
  wire _sub_plot_x_133_in_do;
  wire _sub_plot_x_133_p_reset;
  wire _sub_plot_x_133_m_clock;
  wire [9:0] _sub_plot_x_132_hikareru;
  wire [9:0] _sub_plot_x_132_moto;
  wire [9:0] _sub_plot_x_132_sa;
  wire _sub_plot_x_132_in_do;
  wire _sub_plot_x_132_p_reset;
  wire _sub_plot_x_132_m_clock;
  wire [9:0] _sub_plot_x_131_hikareru;
  wire [9:0] _sub_plot_x_131_moto;
  wire [9:0] _sub_plot_x_131_sa;
  wire _sub_plot_x_131_in_do;
  wire _sub_plot_x_131_p_reset;
  wire _sub_plot_x_131_m_clock;
  wire [9:0] _sub_plot_x_130_hikareru;
  wire [9:0] _sub_plot_x_130_moto;
  wire [9:0] _sub_plot_x_130_sa;
  wire _sub_plot_x_130_in_do;
  wire _sub_plot_x_130_p_reset;
  wire _sub_plot_x_130_m_clock;
  wire [9:0] _sub_plot_x_129_hikareru;
  wire [9:0] _sub_plot_x_129_moto;
  wire [9:0] _sub_plot_x_129_sa;
  wire _sub_plot_x_129_in_do;
  wire _sub_plot_x_129_p_reset;
  wire _sub_plot_x_129_m_clock;
  wire [9:0] _sub_plot_x_128_hikareru;
  wire [9:0] _sub_plot_x_128_moto;
  wire [9:0] _sub_plot_x_128_sa;
  wire _sub_plot_x_128_in_do;
  wire _sub_plot_x_128_p_reset;
  wire _sub_plot_x_128_m_clock;
  wire [9:0] _sub_plot_x_127_hikareru;
  wire [9:0] _sub_plot_x_127_moto;
  wire [9:0] _sub_plot_x_127_sa;
  wire _sub_plot_x_127_in_do;
  wire _sub_plot_x_127_p_reset;
  wire _sub_plot_x_127_m_clock;
  wire [9:0] _sub_plot_x_126_hikareru;
  wire [9:0] _sub_plot_x_126_moto;
  wire [9:0] _sub_plot_x_126_sa;
  wire _sub_plot_x_126_in_do;
  wire _sub_plot_x_126_p_reset;
  wire _sub_plot_x_126_m_clock;
  wire [9:0] _sub_plot_x_125_hikareru;
  wire [9:0] _sub_plot_x_125_moto;
  wire [9:0] _sub_plot_x_125_sa;
  wire _sub_plot_x_125_in_do;
  wire _sub_plot_x_125_p_reset;
  wire _sub_plot_x_125_m_clock;
  wire [9:0] _sub_plot_x_124_hikareru;
  wire [9:0] _sub_plot_x_124_moto;
  wire [9:0] _sub_plot_x_124_sa;
  wire _sub_plot_x_124_in_do;
  wire _sub_plot_x_124_p_reset;
  wire _sub_plot_x_124_m_clock;
  wire [9:0] _sub_plot_x_123_hikareru;
  wire [9:0] _sub_plot_x_123_moto;
  wire [9:0] _sub_plot_x_123_sa;
  wire _sub_plot_x_123_in_do;
  wire _sub_plot_x_123_p_reset;
  wire _sub_plot_x_123_m_clock;
  wire [9:0] _sub_plot_x_122_hikareru;
  wire [9:0] _sub_plot_x_122_moto;
  wire [9:0] _sub_plot_x_122_sa;
  wire _sub_plot_x_122_in_do;
  wire _sub_plot_x_122_p_reset;
  wire _sub_plot_x_122_m_clock;
  wire [9:0] _sub_plot_x_121_hikareru;
  wire [9:0] _sub_plot_x_121_moto;
  wire [9:0] _sub_plot_x_121_sa;
  wire _sub_plot_x_121_in_do;
  wire _sub_plot_x_121_p_reset;
  wire _sub_plot_x_121_m_clock;
  wire [9:0] _sub_plot_x_120_hikareru;
  wire [9:0] _sub_plot_x_120_moto;
  wire [9:0] _sub_plot_x_120_sa;
  wire _sub_plot_x_120_in_do;
  wire _sub_plot_x_120_p_reset;
  wire _sub_plot_x_120_m_clock;
  wire [9:0] _sub_plot_x_119_hikareru;
  wire [9:0] _sub_plot_x_119_moto;
  wire [9:0] _sub_plot_x_119_sa;
  wire _sub_plot_x_119_in_do;
  wire _sub_plot_x_119_p_reset;
  wire _sub_plot_x_119_m_clock;
  wire [9:0] _sub_plot_x_118_hikareru;
  wire [9:0] _sub_plot_x_118_moto;
  wire [9:0] _sub_plot_x_118_sa;
  wire _sub_plot_x_118_in_do;
  wire _sub_plot_x_118_p_reset;
  wire _sub_plot_x_118_m_clock;
  wire [9:0] _sub_plot_x_117_hikareru;
  wire [9:0] _sub_plot_x_117_moto;
  wire [9:0] _sub_plot_x_117_sa;
  wire _sub_plot_x_117_in_do;
  wire _sub_plot_x_117_p_reset;
  wire _sub_plot_x_117_m_clock;
  wire [9:0] _sub_plot_x_116_hikareru;
  wire [9:0] _sub_plot_x_116_moto;
  wire [9:0] _sub_plot_x_116_sa;
  wire _sub_plot_x_116_in_do;
  wire _sub_plot_x_116_p_reset;
  wire _sub_plot_x_116_m_clock;
  wire [9:0] _sub_plot_x_115_hikareru;
  wire [9:0] _sub_plot_x_115_moto;
  wire [9:0] _sub_plot_x_115_sa;
  wire _sub_plot_x_115_in_do;
  wire _sub_plot_x_115_p_reset;
  wire _sub_plot_x_115_m_clock;
  wire [9:0] _sub_plot_x_114_hikareru;
  wire [9:0] _sub_plot_x_114_moto;
  wire [9:0] _sub_plot_x_114_sa;
  wire _sub_plot_x_114_in_do;
  wire _sub_plot_x_114_p_reset;
  wire _sub_plot_x_114_m_clock;
  wire [9:0] _sub_plot_x_113_hikareru;
  wire [9:0] _sub_plot_x_113_moto;
  wire [9:0] _sub_plot_x_113_sa;
  wire _sub_plot_x_113_in_do;
  wire _sub_plot_x_113_p_reset;
  wire _sub_plot_x_113_m_clock;
  wire [9:0] _sub_plot_x_112_hikareru;
  wire [9:0] _sub_plot_x_112_moto;
  wire [9:0] _sub_plot_x_112_sa;
  wire _sub_plot_x_112_in_do;
  wire _sub_plot_x_112_p_reset;
  wire _sub_plot_x_112_m_clock;
  wire [9:0] _sub_plot_x_111_hikareru;
  wire [9:0] _sub_plot_x_111_moto;
  wire [9:0] _sub_plot_x_111_sa;
  wire _sub_plot_x_111_in_do;
  wire _sub_plot_x_111_p_reset;
  wire _sub_plot_x_111_m_clock;
  wire [9:0] _sub_plot_x_110_hikareru;
  wire [9:0] _sub_plot_x_110_moto;
  wire [9:0] _sub_plot_x_110_sa;
  wire _sub_plot_x_110_in_do;
  wire _sub_plot_x_110_p_reset;
  wire _sub_plot_x_110_m_clock;
  wire [9:0] _sub_plot_x_109_hikareru;
  wire [9:0] _sub_plot_x_109_moto;
  wire [9:0] _sub_plot_x_109_sa;
  wire _sub_plot_x_109_in_do;
  wire _sub_plot_x_109_p_reset;
  wire _sub_plot_x_109_m_clock;
  wire [9:0] _sub_plot_x_108_hikareru;
  wire [9:0] _sub_plot_x_108_moto;
  wire [9:0] _sub_plot_x_108_sa;
  wire _sub_plot_x_108_in_do;
  wire _sub_plot_x_108_p_reset;
  wire _sub_plot_x_108_m_clock;
  wire [9:0] _sub_plot_x_107_hikareru;
  wire [9:0] _sub_plot_x_107_moto;
  wire [9:0] _sub_plot_x_107_sa;
  wire _sub_plot_x_107_in_do;
  wire _sub_plot_x_107_p_reset;
  wire _sub_plot_x_107_m_clock;
  wire [9:0] _sub_plot_x_106_hikareru;
  wire [9:0] _sub_plot_x_106_moto;
  wire [9:0] _sub_plot_x_106_sa;
  wire _sub_plot_x_106_in_do;
  wire _sub_plot_x_106_p_reset;
  wire _sub_plot_x_106_m_clock;
  wire [9:0] _sub_plot_x_105_hikareru;
  wire [9:0] _sub_plot_x_105_moto;
  wire [9:0] _sub_plot_x_105_sa;
  wire _sub_plot_x_105_in_do;
  wire _sub_plot_x_105_p_reset;
  wire _sub_plot_x_105_m_clock;
  wire [9:0] _sub_plot_x_104_hikareru;
  wire [9:0] _sub_plot_x_104_moto;
  wire [9:0] _sub_plot_x_104_sa;
  wire _sub_plot_x_104_in_do;
  wire _sub_plot_x_104_p_reset;
  wire _sub_plot_x_104_m_clock;
  wire [9:0] _sub_plot_x_103_hikareru;
  wire [9:0] _sub_plot_x_103_moto;
  wire [9:0] _sub_plot_x_103_sa;
  wire _sub_plot_x_103_in_do;
  wire _sub_plot_x_103_p_reset;
  wire _sub_plot_x_103_m_clock;
  wire [9:0] _sub_plot_x_102_hikareru;
  wire [9:0] _sub_plot_x_102_moto;
  wire [9:0] _sub_plot_x_102_sa;
  wire _sub_plot_x_102_in_do;
  wire _sub_plot_x_102_p_reset;
  wire _sub_plot_x_102_m_clock;
  wire [9:0] _sub_plot_x_101_hikareru;
  wire [9:0] _sub_plot_x_101_moto;
  wire [9:0] _sub_plot_x_101_sa;
  wire _sub_plot_x_101_in_do;
  wire _sub_plot_x_101_p_reset;
  wire _sub_plot_x_101_m_clock;
  wire [9:0] _sub_plot_x_100_hikareru;
  wire [9:0] _sub_plot_x_100_moto;
  wire [9:0] _sub_plot_x_100_sa;
  wire _sub_plot_x_100_in_do;
  wire _sub_plot_x_100_p_reset;
  wire _sub_plot_x_100_m_clock;
  wire [9:0] _sub_plot_x_99_hikareru;
  wire [9:0] _sub_plot_x_99_moto;
  wire [9:0] _sub_plot_x_99_sa;
  wire _sub_plot_x_99_in_do;
  wire _sub_plot_x_99_p_reset;
  wire _sub_plot_x_99_m_clock;
  wire [9:0] _sub_plot_x_98_hikareru;
  wire [9:0] _sub_plot_x_98_moto;
  wire [9:0] _sub_plot_x_98_sa;
  wire _sub_plot_x_98_in_do;
  wire _sub_plot_x_98_p_reset;
  wire _sub_plot_x_98_m_clock;
  wire [9:0] _sub_plot_x_97_hikareru;
  wire [9:0] _sub_plot_x_97_moto;
  wire [9:0] _sub_plot_x_97_sa;
  wire _sub_plot_x_97_in_do;
  wire _sub_plot_x_97_p_reset;
  wire _sub_plot_x_97_m_clock;
  wire [9:0] _sub_plot_x_96_hikareru;
  wire [9:0] _sub_plot_x_96_moto;
  wire [9:0] _sub_plot_x_96_sa;
  wire _sub_plot_x_96_in_do;
  wire _sub_plot_x_96_p_reset;
  wire _sub_plot_x_96_m_clock;
  wire [9:0] _sub_plot_x_95_hikareru;
  wire [9:0] _sub_plot_x_95_moto;
  wire [9:0] _sub_plot_x_95_sa;
  wire _sub_plot_x_95_in_do;
  wire _sub_plot_x_95_p_reset;
  wire _sub_plot_x_95_m_clock;
  wire [9:0] _sub_plot_x_94_hikareru;
  wire [9:0] _sub_plot_x_94_moto;
  wire [9:0] _sub_plot_x_94_sa;
  wire _sub_plot_x_94_in_do;
  wire _sub_plot_x_94_p_reset;
  wire _sub_plot_x_94_m_clock;
  wire [9:0] _sub_plot_x_93_hikareru;
  wire [9:0] _sub_plot_x_93_moto;
  wire [9:0] _sub_plot_x_93_sa;
  wire _sub_plot_x_93_in_do;
  wire _sub_plot_x_93_p_reset;
  wire _sub_plot_x_93_m_clock;
  wire [9:0] _sub_plot_x_92_hikareru;
  wire [9:0] _sub_plot_x_92_moto;
  wire [9:0] _sub_plot_x_92_sa;
  wire _sub_plot_x_92_in_do;
  wire _sub_plot_x_92_p_reset;
  wire _sub_plot_x_92_m_clock;
  wire [9:0] _sub_plot_x_91_hikareru;
  wire [9:0] _sub_plot_x_91_moto;
  wire [9:0] _sub_plot_x_91_sa;
  wire _sub_plot_x_91_in_do;
  wire _sub_plot_x_91_p_reset;
  wire _sub_plot_x_91_m_clock;
  wire [9:0] _sub_plot_x_90_hikareru;
  wire [9:0] _sub_plot_x_90_moto;
  wire [9:0] _sub_plot_x_90_sa;
  wire _sub_plot_x_90_in_do;
  wire _sub_plot_x_90_p_reset;
  wire _sub_plot_x_90_m_clock;
  wire [9:0] _sub_plot_x_89_hikareru;
  wire [9:0] _sub_plot_x_89_moto;
  wire [9:0] _sub_plot_x_89_sa;
  wire _sub_plot_x_89_in_do;
  wire _sub_plot_x_89_p_reset;
  wire _sub_plot_x_89_m_clock;
  wire [9:0] _sub_plot_x_88_hikareru;
  wire [9:0] _sub_plot_x_88_moto;
  wire [9:0] _sub_plot_x_88_sa;
  wire _sub_plot_x_88_in_do;
  wire _sub_plot_x_88_p_reset;
  wire _sub_plot_x_88_m_clock;
  wire [9:0] _sub_plot_x_87_hikareru;
  wire [9:0] _sub_plot_x_87_moto;
  wire [9:0] _sub_plot_x_87_sa;
  wire _sub_plot_x_87_in_do;
  wire _sub_plot_x_87_p_reset;
  wire _sub_plot_x_87_m_clock;
  wire [9:0] _sub_plot_x_86_hikareru;
  wire [9:0] _sub_plot_x_86_moto;
  wire [9:0] _sub_plot_x_86_sa;
  wire _sub_plot_x_86_in_do;
  wire _sub_plot_x_86_p_reset;
  wire _sub_plot_x_86_m_clock;
  wire [9:0] _sub_plot_x_85_hikareru;
  wire [9:0] _sub_plot_x_85_moto;
  wire [9:0] _sub_plot_x_85_sa;
  wire _sub_plot_x_85_in_do;
  wire _sub_plot_x_85_p_reset;
  wire _sub_plot_x_85_m_clock;
  wire [9:0] _sub_plot_x_84_hikareru;
  wire [9:0] _sub_plot_x_84_moto;
  wire [9:0] _sub_plot_x_84_sa;
  wire _sub_plot_x_84_in_do;
  wire _sub_plot_x_84_p_reset;
  wire _sub_plot_x_84_m_clock;
  wire [9:0] _sub_plot_x_83_hikareru;
  wire [9:0] _sub_plot_x_83_moto;
  wire [9:0] _sub_plot_x_83_sa;
  wire _sub_plot_x_83_in_do;
  wire _sub_plot_x_83_p_reset;
  wire _sub_plot_x_83_m_clock;
  wire [9:0] _sub_plot_x_82_hikareru;
  wire [9:0] _sub_plot_x_82_moto;
  wire [9:0] _sub_plot_x_82_sa;
  wire _sub_plot_x_82_in_do;
  wire _sub_plot_x_82_p_reset;
  wire _sub_plot_x_82_m_clock;
  wire [9:0] _sub_plot_x_81_hikareru;
  wire [9:0] _sub_plot_x_81_moto;
  wire [9:0] _sub_plot_x_81_sa;
  wire _sub_plot_x_81_in_do;
  wire _sub_plot_x_81_p_reset;
  wire _sub_plot_x_81_m_clock;
  wire [9:0] _sub_plot_x_80_hikareru;
  wire [9:0] _sub_plot_x_80_moto;
  wire [9:0] _sub_plot_x_80_sa;
  wire _sub_plot_x_80_in_do;
  wire _sub_plot_x_80_p_reset;
  wire _sub_plot_x_80_m_clock;
  wire [9:0] _sub_plot_x_79_hikareru;
  wire [9:0] _sub_plot_x_79_moto;
  wire [9:0] _sub_plot_x_79_sa;
  wire _sub_plot_x_79_in_do;
  wire _sub_plot_x_79_p_reset;
  wire _sub_plot_x_79_m_clock;
  wire [9:0] _sub_plot_x_78_hikareru;
  wire [9:0] _sub_plot_x_78_moto;
  wire [9:0] _sub_plot_x_78_sa;
  wire _sub_plot_x_78_in_do;
  wire _sub_plot_x_78_p_reset;
  wire _sub_plot_x_78_m_clock;
  wire [9:0] _sub_plot_x_77_hikareru;
  wire [9:0] _sub_plot_x_77_moto;
  wire [9:0] _sub_plot_x_77_sa;
  wire _sub_plot_x_77_in_do;
  wire _sub_plot_x_77_p_reset;
  wire _sub_plot_x_77_m_clock;
  wire [9:0] _sub_plot_x_76_hikareru;
  wire [9:0] _sub_plot_x_76_moto;
  wire [9:0] _sub_plot_x_76_sa;
  wire _sub_plot_x_76_in_do;
  wire _sub_plot_x_76_p_reset;
  wire _sub_plot_x_76_m_clock;
  wire [9:0] _sub_plot_x_75_hikareru;
  wire [9:0] _sub_plot_x_75_moto;
  wire [9:0] _sub_plot_x_75_sa;
  wire _sub_plot_x_75_in_do;
  wire _sub_plot_x_75_p_reset;
  wire _sub_plot_x_75_m_clock;
  wire [9:0] _sub_plot_x_74_hikareru;
  wire [9:0] _sub_plot_x_74_moto;
  wire [9:0] _sub_plot_x_74_sa;
  wire _sub_plot_x_74_in_do;
  wire _sub_plot_x_74_p_reset;
  wire _sub_plot_x_74_m_clock;
  wire [9:0] _sub_plot_x_73_hikareru;
  wire [9:0] _sub_plot_x_73_moto;
  wire [9:0] _sub_plot_x_73_sa;
  wire _sub_plot_x_73_in_do;
  wire _sub_plot_x_73_p_reset;
  wire _sub_plot_x_73_m_clock;
  wire [9:0] _sub_plot_x_72_hikareru;
  wire [9:0] _sub_plot_x_72_moto;
  wire [9:0] _sub_plot_x_72_sa;
  wire _sub_plot_x_72_in_do;
  wire _sub_plot_x_72_p_reset;
  wire _sub_plot_x_72_m_clock;
  wire [9:0] _sub_plot_x_71_hikareru;
  wire [9:0] _sub_plot_x_71_moto;
  wire [9:0] _sub_plot_x_71_sa;
  wire _sub_plot_x_71_in_do;
  wire _sub_plot_x_71_p_reset;
  wire _sub_plot_x_71_m_clock;
  wire [9:0] _sub_plot_x_70_hikareru;
  wire [9:0] _sub_plot_x_70_moto;
  wire [9:0] _sub_plot_x_70_sa;
  wire _sub_plot_x_70_in_do;
  wire _sub_plot_x_70_p_reset;
  wire _sub_plot_x_70_m_clock;
  wire [9:0] _sub_plot_x_69_hikareru;
  wire [9:0] _sub_plot_x_69_moto;
  wire [9:0] _sub_plot_x_69_sa;
  wire _sub_plot_x_69_in_do;
  wire _sub_plot_x_69_p_reset;
  wire _sub_plot_x_69_m_clock;
  wire [9:0] _sub_plot_x_68_hikareru;
  wire [9:0] _sub_plot_x_68_moto;
  wire [9:0] _sub_plot_x_68_sa;
  wire _sub_plot_x_68_in_do;
  wire _sub_plot_x_68_p_reset;
  wire _sub_plot_x_68_m_clock;
  wire [9:0] _sub_plot_x_67_hikareru;
  wire [9:0] _sub_plot_x_67_moto;
  wire [9:0] _sub_plot_x_67_sa;
  wire _sub_plot_x_67_in_do;
  wire _sub_plot_x_67_p_reset;
  wire _sub_plot_x_67_m_clock;
  wire [9:0] _sub_plot_x_66_hikareru;
  wire [9:0] _sub_plot_x_66_moto;
  wire [9:0] _sub_plot_x_66_sa;
  wire _sub_plot_x_66_in_do;
  wire _sub_plot_x_66_p_reset;
  wire _sub_plot_x_66_m_clock;
  wire [9:0] _sub_plot_x_65_hikareru;
  wire [9:0] _sub_plot_x_65_moto;
  wire [9:0] _sub_plot_x_65_sa;
  wire _sub_plot_x_65_in_do;
  wire _sub_plot_x_65_p_reset;
  wire _sub_plot_x_65_m_clock;
  wire [9:0] _sub_plot_x_64_hikareru;
  wire [9:0] _sub_plot_x_64_moto;
  wire [9:0] _sub_plot_x_64_sa;
  wire _sub_plot_x_64_in_do;
  wire _sub_plot_x_64_p_reset;
  wire _sub_plot_x_64_m_clock;
  wire [9:0] _sub_plot_x_63_hikareru;
  wire [9:0] _sub_plot_x_63_moto;
  wire [9:0] _sub_plot_x_63_sa;
  wire _sub_plot_x_63_in_do;
  wire _sub_plot_x_63_p_reset;
  wire _sub_plot_x_63_m_clock;
  wire [9:0] _sub_plot_x_62_hikareru;
  wire [9:0] _sub_plot_x_62_moto;
  wire [9:0] _sub_plot_x_62_sa;
  wire _sub_plot_x_62_in_do;
  wire _sub_plot_x_62_p_reset;
  wire _sub_plot_x_62_m_clock;
  wire [9:0] _sub_plot_x_61_hikareru;
  wire [9:0] _sub_plot_x_61_moto;
  wire [9:0] _sub_plot_x_61_sa;
  wire _sub_plot_x_61_in_do;
  wire _sub_plot_x_61_p_reset;
  wire _sub_plot_x_61_m_clock;
  wire [9:0] _sub_plot_x_60_hikareru;
  wire [9:0] _sub_plot_x_60_moto;
  wire [9:0] _sub_plot_x_60_sa;
  wire _sub_plot_x_60_in_do;
  wire _sub_plot_x_60_p_reset;
  wire _sub_plot_x_60_m_clock;
  wire [9:0] _sub_plot_x_59_hikareru;
  wire [9:0] _sub_plot_x_59_moto;
  wire [9:0] _sub_plot_x_59_sa;
  wire _sub_plot_x_59_in_do;
  wire _sub_plot_x_59_p_reset;
  wire _sub_plot_x_59_m_clock;
  wire [9:0] _sub_plot_x_58_hikareru;
  wire [9:0] _sub_plot_x_58_moto;
  wire [9:0] _sub_plot_x_58_sa;
  wire _sub_plot_x_58_in_do;
  wire _sub_plot_x_58_p_reset;
  wire _sub_plot_x_58_m_clock;
  wire [9:0] _sub_plot_x_57_hikareru;
  wire [9:0] _sub_plot_x_57_moto;
  wire [9:0] _sub_plot_x_57_sa;
  wire _sub_plot_x_57_in_do;
  wire _sub_plot_x_57_p_reset;
  wire _sub_plot_x_57_m_clock;
  wire [9:0] _sub_plot_x_56_hikareru;
  wire [9:0] _sub_plot_x_56_moto;
  wire [9:0] _sub_plot_x_56_sa;
  wire _sub_plot_x_56_in_do;
  wire _sub_plot_x_56_p_reset;
  wire _sub_plot_x_56_m_clock;
  wire [9:0] _sub_plot_x_55_hikareru;
  wire [9:0] _sub_plot_x_55_moto;
  wire [9:0] _sub_plot_x_55_sa;
  wire _sub_plot_x_55_in_do;
  wire _sub_plot_x_55_p_reset;
  wire _sub_plot_x_55_m_clock;
  wire [9:0] _sub_plot_x_54_hikareru;
  wire [9:0] _sub_plot_x_54_moto;
  wire [9:0] _sub_plot_x_54_sa;
  wire _sub_plot_x_54_in_do;
  wire _sub_plot_x_54_p_reset;
  wire _sub_plot_x_54_m_clock;
  wire [9:0] _sub_plot_x_53_hikareru;
  wire [9:0] _sub_plot_x_53_moto;
  wire [9:0] _sub_plot_x_53_sa;
  wire _sub_plot_x_53_in_do;
  wire _sub_plot_x_53_p_reset;
  wire _sub_plot_x_53_m_clock;
  wire [9:0] _sub_plot_x_52_hikareru;
  wire [9:0] _sub_plot_x_52_moto;
  wire [9:0] _sub_plot_x_52_sa;
  wire _sub_plot_x_52_in_do;
  wire _sub_plot_x_52_p_reset;
  wire _sub_plot_x_52_m_clock;
  wire [9:0] _sub_plot_x_51_hikareru;
  wire [9:0] _sub_plot_x_51_moto;
  wire [9:0] _sub_plot_x_51_sa;
  wire _sub_plot_x_51_in_do;
  wire _sub_plot_x_51_p_reset;
  wire _sub_plot_x_51_m_clock;
  wire [9:0] _sub_plot_x_50_hikareru;
  wire [9:0] _sub_plot_x_50_moto;
  wire [9:0] _sub_plot_x_50_sa;
  wire _sub_plot_x_50_in_do;
  wire _sub_plot_x_50_p_reset;
  wire _sub_plot_x_50_m_clock;
  wire [9:0] _sub_plot_x_49_hikareru;
  wire [9:0] _sub_plot_x_49_moto;
  wire [9:0] _sub_plot_x_49_sa;
  wire _sub_plot_x_49_in_do;
  wire _sub_plot_x_49_p_reset;
  wire _sub_plot_x_49_m_clock;
  wire [9:0] _sub_plot_x_48_hikareru;
  wire [9:0] _sub_plot_x_48_moto;
  wire [9:0] _sub_plot_x_48_sa;
  wire _sub_plot_x_48_in_do;
  wire _sub_plot_x_48_p_reset;
  wire _sub_plot_x_48_m_clock;
  wire [9:0] _sub_plot_x_47_hikareru;
  wire [9:0] _sub_plot_x_47_moto;
  wire [9:0] _sub_plot_x_47_sa;
  wire _sub_plot_x_47_in_do;
  wire _sub_plot_x_47_p_reset;
  wire _sub_plot_x_47_m_clock;
  wire [9:0] _sub_plot_x_46_hikareru;
  wire [9:0] _sub_plot_x_46_moto;
  wire [9:0] _sub_plot_x_46_sa;
  wire _sub_plot_x_46_in_do;
  wire _sub_plot_x_46_p_reset;
  wire _sub_plot_x_46_m_clock;
  wire [9:0] _sub_plot_x_45_hikareru;
  wire [9:0] _sub_plot_x_45_moto;
  wire [9:0] _sub_plot_x_45_sa;
  wire _sub_plot_x_45_in_do;
  wire _sub_plot_x_45_p_reset;
  wire _sub_plot_x_45_m_clock;
  wire [9:0] _sub_plot_x_44_hikareru;
  wire [9:0] _sub_plot_x_44_moto;
  wire [9:0] _sub_plot_x_44_sa;
  wire _sub_plot_x_44_in_do;
  wire _sub_plot_x_44_p_reset;
  wire _sub_plot_x_44_m_clock;
  wire [9:0] _sub_plot_x_43_hikareru;
  wire [9:0] _sub_plot_x_43_moto;
  wire [9:0] _sub_plot_x_43_sa;
  wire _sub_plot_x_43_in_do;
  wire _sub_plot_x_43_p_reset;
  wire _sub_plot_x_43_m_clock;
  wire [9:0] _sub_plot_x_42_hikareru;
  wire [9:0] _sub_plot_x_42_moto;
  wire [9:0] _sub_plot_x_42_sa;
  wire _sub_plot_x_42_in_do;
  wire _sub_plot_x_42_p_reset;
  wire _sub_plot_x_42_m_clock;
  wire [9:0] _sub_plot_x_41_hikareru;
  wire [9:0] _sub_plot_x_41_moto;
  wire [9:0] _sub_plot_x_41_sa;
  wire _sub_plot_x_41_in_do;
  wire _sub_plot_x_41_p_reset;
  wire _sub_plot_x_41_m_clock;
  wire [9:0] _sub_plot_x_40_hikareru;
  wire [9:0] _sub_plot_x_40_moto;
  wire [9:0] _sub_plot_x_40_sa;
  wire _sub_plot_x_40_in_do;
  wire _sub_plot_x_40_p_reset;
  wire _sub_plot_x_40_m_clock;
  wire [9:0] _sub_plot_x_39_hikareru;
  wire [9:0] _sub_plot_x_39_moto;
  wire [9:0] _sub_plot_x_39_sa;
  wire _sub_plot_x_39_in_do;
  wire _sub_plot_x_39_p_reset;
  wire _sub_plot_x_39_m_clock;
  wire [9:0] _sub_plot_x_38_hikareru;
  wire [9:0] _sub_plot_x_38_moto;
  wire [9:0] _sub_plot_x_38_sa;
  wire _sub_plot_x_38_in_do;
  wire _sub_plot_x_38_p_reset;
  wire _sub_plot_x_38_m_clock;
  wire [9:0] _sub_plot_x_37_hikareru;
  wire [9:0] _sub_plot_x_37_moto;
  wire [9:0] _sub_plot_x_37_sa;
  wire _sub_plot_x_37_in_do;
  wire _sub_plot_x_37_p_reset;
  wire _sub_plot_x_37_m_clock;
  wire [9:0] _sub_plot_x_36_hikareru;
  wire [9:0] _sub_plot_x_36_moto;
  wire [9:0] _sub_plot_x_36_sa;
  wire _sub_plot_x_36_in_do;
  wire _sub_plot_x_36_p_reset;
  wire _sub_plot_x_36_m_clock;
  wire [9:0] _sub_plot_x_35_hikareru;
  wire [9:0] _sub_plot_x_35_moto;
  wire [9:0] _sub_plot_x_35_sa;
  wire _sub_plot_x_35_in_do;
  wire _sub_plot_x_35_p_reset;
  wire _sub_plot_x_35_m_clock;
  wire [9:0] _sub_plot_x_34_hikareru;
  wire [9:0] _sub_plot_x_34_moto;
  wire [9:0] _sub_plot_x_34_sa;
  wire _sub_plot_x_34_in_do;
  wire _sub_plot_x_34_p_reset;
  wire _sub_plot_x_34_m_clock;
  wire [9:0] _sub_plot_x_33_hikareru;
  wire [9:0] _sub_plot_x_33_moto;
  wire [9:0] _sub_plot_x_33_sa;
  wire _sub_plot_x_33_in_do;
  wire _sub_plot_x_33_p_reset;
  wire _sub_plot_x_33_m_clock;
  wire [9:0] _sub_plot_x_32_hikareru;
  wire [9:0] _sub_plot_x_32_moto;
  wire [9:0] _sub_plot_x_32_sa;
  wire _sub_plot_x_32_in_do;
  wire _sub_plot_x_32_p_reset;
  wire _sub_plot_x_32_m_clock;
  wire [9:0] _sub_plot_x_31_hikareru;
  wire [9:0] _sub_plot_x_31_moto;
  wire [9:0] _sub_plot_x_31_sa;
  wire _sub_plot_x_31_in_do;
  wire _sub_plot_x_31_p_reset;
  wire _sub_plot_x_31_m_clock;
  wire [9:0] _sub_plot_x_30_hikareru;
  wire [9:0] _sub_plot_x_30_moto;
  wire [9:0] _sub_plot_x_30_sa;
  wire _sub_plot_x_30_in_do;
  wire _sub_plot_x_30_p_reset;
  wire _sub_plot_x_30_m_clock;
  wire [9:0] _sub_plot_x_29_hikareru;
  wire [9:0] _sub_plot_x_29_moto;
  wire [9:0] _sub_plot_x_29_sa;
  wire _sub_plot_x_29_in_do;
  wire _sub_plot_x_29_p_reset;
  wire _sub_plot_x_29_m_clock;
  wire [9:0] _sub_plot_x_28_hikareru;
  wire [9:0] _sub_plot_x_28_moto;
  wire [9:0] _sub_plot_x_28_sa;
  wire _sub_plot_x_28_in_do;
  wire _sub_plot_x_28_p_reset;
  wire _sub_plot_x_28_m_clock;
  wire [9:0] _sub_plot_x_27_hikareru;
  wire [9:0] _sub_plot_x_27_moto;
  wire [9:0] _sub_plot_x_27_sa;
  wire _sub_plot_x_27_in_do;
  wire _sub_plot_x_27_p_reset;
  wire _sub_plot_x_27_m_clock;
  wire [9:0] _sub_plot_x_26_hikareru;
  wire [9:0] _sub_plot_x_26_moto;
  wire [9:0] _sub_plot_x_26_sa;
  wire _sub_plot_x_26_in_do;
  wire _sub_plot_x_26_p_reset;
  wire _sub_plot_x_26_m_clock;
  wire [9:0] _sub_plot_x_25_hikareru;
  wire [9:0] _sub_plot_x_25_moto;
  wire [9:0] _sub_plot_x_25_sa;
  wire _sub_plot_x_25_in_do;
  wire _sub_plot_x_25_p_reset;
  wire _sub_plot_x_25_m_clock;
  wire [9:0] _sub_plot_x_24_hikareru;
  wire [9:0] _sub_plot_x_24_moto;
  wire [9:0] _sub_plot_x_24_sa;
  wire _sub_plot_x_24_in_do;
  wire _sub_plot_x_24_p_reset;
  wire _sub_plot_x_24_m_clock;
  wire [9:0] _sub_plot_x_23_hikareru;
  wire [9:0] _sub_plot_x_23_moto;
  wire [9:0] _sub_plot_x_23_sa;
  wire _sub_plot_x_23_in_do;
  wire _sub_plot_x_23_p_reset;
  wire _sub_plot_x_23_m_clock;
  wire [9:0] _sub_plot_x_22_hikareru;
  wire [9:0] _sub_plot_x_22_moto;
  wire [9:0] _sub_plot_x_22_sa;
  wire _sub_plot_x_22_in_do;
  wire _sub_plot_x_22_p_reset;
  wire _sub_plot_x_22_m_clock;
  wire [9:0] _sub_plot_x_21_hikareru;
  wire [9:0] _sub_plot_x_21_moto;
  wire [9:0] _sub_plot_x_21_sa;
  wire _sub_plot_x_21_in_do;
  wire _sub_plot_x_21_p_reset;
  wire _sub_plot_x_21_m_clock;
  wire [9:0] _sub_plot_x_20_hikareru;
  wire [9:0] _sub_plot_x_20_moto;
  wire [9:0] _sub_plot_x_20_sa;
  wire _sub_plot_x_20_in_do;
  wire _sub_plot_x_20_p_reset;
  wire _sub_plot_x_20_m_clock;
  wire [9:0] _sub_plot_x_19_hikareru;
  wire [9:0] _sub_plot_x_19_moto;
  wire [9:0] _sub_plot_x_19_sa;
  wire _sub_plot_x_19_in_do;
  wire _sub_plot_x_19_p_reset;
  wire _sub_plot_x_19_m_clock;
  wire [9:0] _sub_plot_x_18_hikareru;
  wire [9:0] _sub_plot_x_18_moto;
  wire [9:0] _sub_plot_x_18_sa;
  wire _sub_plot_x_18_in_do;
  wire _sub_plot_x_18_p_reset;
  wire _sub_plot_x_18_m_clock;
  wire [9:0] _sub_plot_x_17_hikareru;
  wire [9:0] _sub_plot_x_17_moto;
  wire [9:0] _sub_plot_x_17_sa;
  wire _sub_plot_x_17_in_do;
  wire _sub_plot_x_17_p_reset;
  wire _sub_plot_x_17_m_clock;
  wire [9:0] _sub_plot_x_16_hikareru;
  wire [9:0] _sub_plot_x_16_moto;
  wire [9:0] _sub_plot_x_16_sa;
  wire _sub_plot_x_16_in_do;
  wire _sub_plot_x_16_p_reset;
  wire _sub_plot_x_16_m_clock;
  wire [9:0] _sub_plot_x_15_hikareru;
  wire [9:0] _sub_plot_x_15_moto;
  wire [9:0] _sub_plot_x_15_sa;
  wire _sub_plot_x_15_in_do;
  wire _sub_plot_x_15_p_reset;
  wire _sub_plot_x_15_m_clock;
  wire [9:0] _sub_plot_x_14_hikareru;
  wire [9:0] _sub_plot_x_14_moto;
  wire [9:0] _sub_plot_x_14_sa;
  wire _sub_plot_x_14_in_do;
  wire _sub_plot_x_14_p_reset;
  wire _sub_plot_x_14_m_clock;
  wire [9:0] _sub_plot_x_13_hikareru;
  wire [9:0] _sub_plot_x_13_moto;
  wire [9:0] _sub_plot_x_13_sa;
  wire _sub_plot_x_13_in_do;
  wire _sub_plot_x_13_p_reset;
  wire _sub_plot_x_13_m_clock;
  wire [9:0] _sub_plot_x_12_hikareru;
  wire [9:0] _sub_plot_x_12_moto;
  wire [9:0] _sub_plot_x_12_sa;
  wire _sub_plot_x_12_in_do;
  wire _sub_plot_x_12_p_reset;
  wire _sub_plot_x_12_m_clock;
  wire [9:0] _sub_plot_x_11_hikareru;
  wire [9:0] _sub_plot_x_11_moto;
  wire [9:0] _sub_plot_x_11_sa;
  wire _sub_plot_x_11_in_do;
  wire _sub_plot_x_11_p_reset;
  wire _sub_plot_x_11_m_clock;
  wire [9:0] _sub_plot_x_10_hikareru;
  wire [9:0] _sub_plot_x_10_moto;
  wire [9:0] _sub_plot_x_10_sa;
  wire _sub_plot_x_10_in_do;
  wire _sub_plot_x_10_p_reset;
  wire _sub_plot_x_10_m_clock;
  wire [9:0] _sub_plot_x_9_hikareru;
  wire [9:0] _sub_plot_x_9_moto;
  wire [9:0] _sub_plot_x_9_sa;
  wire _sub_plot_x_9_in_do;
  wire _sub_plot_x_9_p_reset;
  wire _sub_plot_x_9_m_clock;
  wire [9:0] _sub_plot_x_8_hikareru;
  wire [9:0] _sub_plot_x_8_moto;
  wire [9:0] _sub_plot_x_8_sa;
  wire _sub_plot_x_8_in_do;
  wire _sub_plot_x_8_p_reset;
  wire _sub_plot_x_8_m_clock;
  wire [9:0] _sub_plot_x_7_hikareru;
  wire [9:0] _sub_plot_x_7_moto;
  wire [9:0] _sub_plot_x_7_sa;
  wire _sub_plot_x_7_in_do;
  wire _sub_plot_x_7_p_reset;
  wire _sub_plot_x_7_m_clock;
  wire [9:0] _sub_plot_x_6_hikareru;
  wire [9:0] _sub_plot_x_6_moto;
  wire [9:0] _sub_plot_x_6_sa;
  wire _sub_plot_x_6_in_do;
  wire _sub_plot_x_6_p_reset;
  wire _sub_plot_x_6_m_clock;
  wire [9:0] _sub_plot_x_5_hikareru;
  wire [9:0] _sub_plot_x_5_moto;
  wire [9:0] _sub_plot_x_5_sa;
  wire _sub_plot_x_5_in_do;
  wire _sub_plot_x_5_p_reset;
  wire _sub_plot_x_5_m_clock;
  wire [9:0] _sub_plot_x_4_hikareru;
  wire [9:0] _sub_plot_x_4_moto;
  wire [9:0] _sub_plot_x_4_sa;
  wire _sub_plot_x_4_in_do;
  wire _sub_plot_x_4_p_reset;
  wire _sub_plot_x_4_m_clock;
  wire [9:0] _sub_plot_x_3_hikareru;
  wire [9:0] _sub_plot_x_3_moto;
  wire [9:0] _sub_plot_x_3_sa;
  wire _sub_plot_x_3_in_do;
  wire _sub_plot_x_3_p_reset;
  wire _sub_plot_x_3_m_clock;
  wire [9:0] _sub_plot_x_2_hikareru;
  wire [9:0] _sub_plot_x_2_moto;
  wire [9:0] _sub_plot_x_2_sa;
  wire _sub_plot_x_2_in_do;
  wire _sub_plot_x_2_p_reset;
  wire _sub_plot_x_2_m_clock;
  wire [9:0] _sub_plot_x_1_hikareru;
  wire [9:0] _sub_plot_x_1_moto;
  wire [9:0] _sub_plot_x_1_sa;
  wire _sub_plot_x_1_in_do;
  wire _sub_plot_x_1_p_reset;
  wire _sub_plot_x_1_m_clock;
sub_plot sub_plot_x (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_in_do), .sa(_sub_plot_x_sa), .hikareru(_sub_plot_x_hikareru), .moto(_sub_plot_x_moto));
sub_plot sub_plot_x_209 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_209_in_do), .sa(_sub_plot_x_209_sa), .hikareru(_sub_plot_x_209_hikareru), .moto(_sub_plot_x_209_moto));
sub_plot sub_plot_x_208 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_208_in_do), .sa(_sub_plot_x_208_sa), .hikareru(_sub_plot_x_208_hikareru), .moto(_sub_plot_x_208_moto));
sub_plot sub_plot_x_207 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_207_in_do), .sa(_sub_plot_x_207_sa), .hikareru(_sub_plot_x_207_hikareru), .moto(_sub_plot_x_207_moto));
sub_plot sub_plot_x_206 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_206_in_do), .sa(_sub_plot_x_206_sa), .hikareru(_sub_plot_x_206_hikareru), .moto(_sub_plot_x_206_moto));
sub_plot sub_plot_x_205 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_205_in_do), .sa(_sub_plot_x_205_sa), .hikareru(_sub_plot_x_205_hikareru), .moto(_sub_plot_x_205_moto));
sub_plot sub_plot_x_204 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_204_in_do), .sa(_sub_plot_x_204_sa), .hikareru(_sub_plot_x_204_hikareru), .moto(_sub_plot_x_204_moto));
sub_plot sub_plot_x_203 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_203_in_do), .sa(_sub_plot_x_203_sa), .hikareru(_sub_plot_x_203_hikareru), .moto(_sub_plot_x_203_moto));
sub_plot sub_plot_x_202 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_202_in_do), .sa(_sub_plot_x_202_sa), .hikareru(_sub_plot_x_202_hikareru), .moto(_sub_plot_x_202_moto));
sub_plot sub_plot_x_201 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_201_in_do), .sa(_sub_plot_x_201_sa), .hikareru(_sub_plot_x_201_hikareru), .moto(_sub_plot_x_201_moto));
sub_plot sub_plot_x_200 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_200_in_do), .sa(_sub_plot_x_200_sa), .hikareru(_sub_plot_x_200_hikareru), .moto(_sub_plot_x_200_moto));
sub_plot sub_plot_x_199 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_199_in_do), .sa(_sub_plot_x_199_sa), .hikareru(_sub_plot_x_199_hikareru), .moto(_sub_plot_x_199_moto));
sub_plot sub_plot_x_198 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_198_in_do), .sa(_sub_plot_x_198_sa), .hikareru(_sub_plot_x_198_hikareru), .moto(_sub_plot_x_198_moto));
sub_plot sub_plot_x_197 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_197_in_do), .sa(_sub_plot_x_197_sa), .hikareru(_sub_plot_x_197_hikareru), .moto(_sub_plot_x_197_moto));
sub_plot sub_plot_x_196 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_196_in_do), .sa(_sub_plot_x_196_sa), .hikareru(_sub_plot_x_196_hikareru), .moto(_sub_plot_x_196_moto));
sub_plot sub_plot_x_195 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_195_in_do), .sa(_sub_plot_x_195_sa), .hikareru(_sub_plot_x_195_hikareru), .moto(_sub_plot_x_195_moto));
sub_plot sub_plot_x_194 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_194_in_do), .sa(_sub_plot_x_194_sa), .hikareru(_sub_plot_x_194_hikareru), .moto(_sub_plot_x_194_moto));
sub_plot sub_plot_x_193 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_193_in_do), .sa(_sub_plot_x_193_sa), .hikareru(_sub_plot_x_193_hikareru), .moto(_sub_plot_x_193_moto));
sub_plot sub_plot_x_192 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_192_in_do), .sa(_sub_plot_x_192_sa), .hikareru(_sub_plot_x_192_hikareru), .moto(_sub_plot_x_192_moto));
sub_plot sub_plot_x_191 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_191_in_do), .sa(_sub_plot_x_191_sa), .hikareru(_sub_plot_x_191_hikareru), .moto(_sub_plot_x_191_moto));
sub_plot sub_plot_x_190 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_190_in_do), .sa(_sub_plot_x_190_sa), .hikareru(_sub_plot_x_190_hikareru), .moto(_sub_plot_x_190_moto));
sub_plot sub_plot_x_189 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_189_in_do), .sa(_sub_plot_x_189_sa), .hikareru(_sub_plot_x_189_hikareru), .moto(_sub_plot_x_189_moto));
sub_plot sub_plot_x_188 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_188_in_do), .sa(_sub_plot_x_188_sa), .hikareru(_sub_plot_x_188_hikareru), .moto(_sub_plot_x_188_moto));
sub_plot sub_plot_x_187 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_187_in_do), .sa(_sub_plot_x_187_sa), .hikareru(_sub_plot_x_187_hikareru), .moto(_sub_plot_x_187_moto));
sub_plot sub_plot_x_186 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_186_in_do), .sa(_sub_plot_x_186_sa), .hikareru(_sub_plot_x_186_hikareru), .moto(_sub_plot_x_186_moto));
sub_plot sub_plot_x_185 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_185_in_do), .sa(_sub_plot_x_185_sa), .hikareru(_sub_plot_x_185_hikareru), .moto(_sub_plot_x_185_moto));
sub_plot sub_plot_x_184 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_184_in_do), .sa(_sub_plot_x_184_sa), .hikareru(_sub_plot_x_184_hikareru), .moto(_sub_plot_x_184_moto));
sub_plot sub_plot_x_183 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_183_in_do), .sa(_sub_plot_x_183_sa), .hikareru(_sub_plot_x_183_hikareru), .moto(_sub_plot_x_183_moto));
sub_plot sub_plot_x_182 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_182_in_do), .sa(_sub_plot_x_182_sa), .hikareru(_sub_plot_x_182_hikareru), .moto(_sub_plot_x_182_moto));
sub_plot sub_plot_x_181 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_181_in_do), .sa(_sub_plot_x_181_sa), .hikareru(_sub_plot_x_181_hikareru), .moto(_sub_plot_x_181_moto));
sub_plot sub_plot_x_180 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_180_in_do), .sa(_sub_plot_x_180_sa), .hikareru(_sub_plot_x_180_hikareru), .moto(_sub_plot_x_180_moto));
sub_plot sub_plot_x_179 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_179_in_do), .sa(_sub_plot_x_179_sa), .hikareru(_sub_plot_x_179_hikareru), .moto(_sub_plot_x_179_moto));
sub_plot sub_plot_x_178 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_178_in_do), .sa(_sub_plot_x_178_sa), .hikareru(_sub_plot_x_178_hikareru), .moto(_sub_plot_x_178_moto));
sub_plot sub_plot_x_177 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_177_in_do), .sa(_sub_plot_x_177_sa), .hikareru(_sub_plot_x_177_hikareru), .moto(_sub_plot_x_177_moto));
sub_plot sub_plot_x_176 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_176_in_do), .sa(_sub_plot_x_176_sa), .hikareru(_sub_plot_x_176_hikareru), .moto(_sub_plot_x_176_moto));
sub_plot sub_plot_x_175 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_175_in_do), .sa(_sub_plot_x_175_sa), .hikareru(_sub_plot_x_175_hikareru), .moto(_sub_plot_x_175_moto));
sub_plot sub_plot_x_174 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_174_in_do), .sa(_sub_plot_x_174_sa), .hikareru(_sub_plot_x_174_hikareru), .moto(_sub_plot_x_174_moto));
sub_plot sub_plot_x_173 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_173_in_do), .sa(_sub_plot_x_173_sa), .hikareru(_sub_plot_x_173_hikareru), .moto(_sub_plot_x_173_moto));
sub_plot sub_plot_x_172 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_172_in_do), .sa(_sub_plot_x_172_sa), .hikareru(_sub_plot_x_172_hikareru), .moto(_sub_plot_x_172_moto));
sub_plot sub_plot_x_171 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_171_in_do), .sa(_sub_plot_x_171_sa), .hikareru(_sub_plot_x_171_hikareru), .moto(_sub_plot_x_171_moto));
sub_plot sub_plot_x_170 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_170_in_do), .sa(_sub_plot_x_170_sa), .hikareru(_sub_plot_x_170_hikareru), .moto(_sub_plot_x_170_moto));
sub_plot sub_plot_x_169 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_169_in_do), .sa(_sub_plot_x_169_sa), .hikareru(_sub_plot_x_169_hikareru), .moto(_sub_plot_x_169_moto));
sub_plot sub_plot_x_168 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_168_in_do), .sa(_sub_plot_x_168_sa), .hikareru(_sub_plot_x_168_hikareru), .moto(_sub_plot_x_168_moto));
sub_plot sub_plot_x_167 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_167_in_do), .sa(_sub_plot_x_167_sa), .hikareru(_sub_plot_x_167_hikareru), .moto(_sub_plot_x_167_moto));
sub_plot sub_plot_x_166 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_166_in_do), .sa(_sub_plot_x_166_sa), .hikareru(_sub_plot_x_166_hikareru), .moto(_sub_plot_x_166_moto));
sub_plot sub_plot_x_165 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_165_in_do), .sa(_sub_plot_x_165_sa), .hikareru(_sub_plot_x_165_hikareru), .moto(_sub_plot_x_165_moto));
sub_plot sub_plot_x_164 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_164_in_do), .sa(_sub_plot_x_164_sa), .hikareru(_sub_plot_x_164_hikareru), .moto(_sub_plot_x_164_moto));
sub_plot sub_plot_x_163 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_163_in_do), .sa(_sub_plot_x_163_sa), .hikareru(_sub_plot_x_163_hikareru), .moto(_sub_plot_x_163_moto));
sub_plot sub_plot_x_162 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_162_in_do), .sa(_sub_plot_x_162_sa), .hikareru(_sub_plot_x_162_hikareru), .moto(_sub_plot_x_162_moto));
sub_plot sub_plot_x_161 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_161_in_do), .sa(_sub_plot_x_161_sa), .hikareru(_sub_plot_x_161_hikareru), .moto(_sub_plot_x_161_moto));
sub_plot sub_plot_x_160 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_160_in_do), .sa(_sub_plot_x_160_sa), .hikareru(_sub_plot_x_160_hikareru), .moto(_sub_plot_x_160_moto));
sub_plot sub_plot_x_159 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_159_in_do), .sa(_sub_plot_x_159_sa), .hikareru(_sub_plot_x_159_hikareru), .moto(_sub_plot_x_159_moto));
sub_plot sub_plot_x_158 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_158_in_do), .sa(_sub_plot_x_158_sa), .hikareru(_sub_plot_x_158_hikareru), .moto(_sub_plot_x_158_moto));
sub_plot sub_plot_x_157 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_157_in_do), .sa(_sub_plot_x_157_sa), .hikareru(_sub_plot_x_157_hikareru), .moto(_sub_plot_x_157_moto));
sub_plot sub_plot_x_156 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_156_in_do), .sa(_sub_plot_x_156_sa), .hikareru(_sub_plot_x_156_hikareru), .moto(_sub_plot_x_156_moto));
sub_plot sub_plot_x_155 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_155_in_do), .sa(_sub_plot_x_155_sa), .hikareru(_sub_plot_x_155_hikareru), .moto(_sub_plot_x_155_moto));
sub_plot sub_plot_x_154 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_154_in_do), .sa(_sub_plot_x_154_sa), .hikareru(_sub_plot_x_154_hikareru), .moto(_sub_plot_x_154_moto));
sub_plot sub_plot_x_153 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_153_in_do), .sa(_sub_plot_x_153_sa), .hikareru(_sub_plot_x_153_hikareru), .moto(_sub_plot_x_153_moto));
sub_plot sub_plot_x_152 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_152_in_do), .sa(_sub_plot_x_152_sa), .hikareru(_sub_plot_x_152_hikareru), .moto(_sub_plot_x_152_moto));
sub_plot sub_plot_x_151 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_151_in_do), .sa(_sub_plot_x_151_sa), .hikareru(_sub_plot_x_151_hikareru), .moto(_sub_plot_x_151_moto));
sub_plot sub_plot_x_150 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_150_in_do), .sa(_sub_plot_x_150_sa), .hikareru(_sub_plot_x_150_hikareru), .moto(_sub_plot_x_150_moto));
sub_plot sub_plot_x_149 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_149_in_do), .sa(_sub_plot_x_149_sa), .hikareru(_sub_plot_x_149_hikareru), .moto(_sub_plot_x_149_moto));
sub_plot sub_plot_x_148 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_148_in_do), .sa(_sub_plot_x_148_sa), .hikareru(_sub_plot_x_148_hikareru), .moto(_sub_plot_x_148_moto));
sub_plot sub_plot_x_147 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_147_in_do), .sa(_sub_plot_x_147_sa), .hikareru(_sub_plot_x_147_hikareru), .moto(_sub_plot_x_147_moto));
sub_plot sub_plot_x_146 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_146_in_do), .sa(_sub_plot_x_146_sa), .hikareru(_sub_plot_x_146_hikareru), .moto(_sub_plot_x_146_moto));
sub_plot sub_plot_x_145 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_145_in_do), .sa(_sub_plot_x_145_sa), .hikareru(_sub_plot_x_145_hikareru), .moto(_sub_plot_x_145_moto));
sub_plot sub_plot_x_144 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_144_in_do), .sa(_sub_plot_x_144_sa), .hikareru(_sub_plot_x_144_hikareru), .moto(_sub_plot_x_144_moto));
sub_plot sub_plot_x_143 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_143_in_do), .sa(_sub_plot_x_143_sa), .hikareru(_sub_plot_x_143_hikareru), .moto(_sub_plot_x_143_moto));
sub_plot sub_plot_x_142 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_142_in_do), .sa(_sub_plot_x_142_sa), .hikareru(_sub_plot_x_142_hikareru), .moto(_sub_plot_x_142_moto));
sub_plot sub_plot_x_141 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_141_in_do), .sa(_sub_plot_x_141_sa), .hikareru(_sub_plot_x_141_hikareru), .moto(_sub_plot_x_141_moto));
sub_plot sub_plot_x_140 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_140_in_do), .sa(_sub_plot_x_140_sa), .hikareru(_sub_plot_x_140_hikareru), .moto(_sub_plot_x_140_moto));
sub_plot sub_plot_x_139 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_139_in_do), .sa(_sub_plot_x_139_sa), .hikareru(_sub_plot_x_139_hikareru), .moto(_sub_plot_x_139_moto));
sub_plot sub_plot_x_138 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_138_in_do), .sa(_sub_plot_x_138_sa), .hikareru(_sub_plot_x_138_hikareru), .moto(_sub_plot_x_138_moto));
sub_plot sub_plot_x_137 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_137_in_do), .sa(_sub_plot_x_137_sa), .hikareru(_sub_plot_x_137_hikareru), .moto(_sub_plot_x_137_moto));
sub_plot sub_plot_x_136 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_136_in_do), .sa(_sub_plot_x_136_sa), .hikareru(_sub_plot_x_136_hikareru), .moto(_sub_plot_x_136_moto));
sub_plot sub_plot_x_135 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_135_in_do), .sa(_sub_plot_x_135_sa), .hikareru(_sub_plot_x_135_hikareru), .moto(_sub_plot_x_135_moto));
sub_plot sub_plot_x_134 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_134_in_do), .sa(_sub_plot_x_134_sa), .hikareru(_sub_plot_x_134_hikareru), .moto(_sub_plot_x_134_moto));
sub_plot sub_plot_x_133 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_133_in_do), .sa(_sub_plot_x_133_sa), .hikareru(_sub_plot_x_133_hikareru), .moto(_sub_plot_x_133_moto));
sub_plot sub_plot_x_132 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_132_in_do), .sa(_sub_plot_x_132_sa), .hikareru(_sub_plot_x_132_hikareru), .moto(_sub_plot_x_132_moto));
sub_plot sub_plot_x_131 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_131_in_do), .sa(_sub_plot_x_131_sa), .hikareru(_sub_plot_x_131_hikareru), .moto(_sub_plot_x_131_moto));
sub_plot sub_plot_x_130 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_130_in_do), .sa(_sub_plot_x_130_sa), .hikareru(_sub_plot_x_130_hikareru), .moto(_sub_plot_x_130_moto));
sub_plot sub_plot_x_129 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_129_in_do), .sa(_sub_plot_x_129_sa), .hikareru(_sub_plot_x_129_hikareru), .moto(_sub_plot_x_129_moto));
sub_plot sub_plot_x_128 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_128_in_do), .sa(_sub_plot_x_128_sa), .hikareru(_sub_plot_x_128_hikareru), .moto(_sub_plot_x_128_moto));
sub_plot sub_plot_x_127 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_127_in_do), .sa(_sub_plot_x_127_sa), .hikareru(_sub_plot_x_127_hikareru), .moto(_sub_plot_x_127_moto));
sub_plot sub_plot_x_126 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_126_in_do), .sa(_sub_plot_x_126_sa), .hikareru(_sub_plot_x_126_hikareru), .moto(_sub_plot_x_126_moto));
sub_plot sub_plot_x_125 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_125_in_do), .sa(_sub_plot_x_125_sa), .hikareru(_sub_plot_x_125_hikareru), .moto(_sub_plot_x_125_moto));
sub_plot sub_plot_x_124 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_124_in_do), .sa(_sub_plot_x_124_sa), .hikareru(_sub_plot_x_124_hikareru), .moto(_sub_plot_x_124_moto));
sub_plot sub_plot_x_123 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_123_in_do), .sa(_sub_plot_x_123_sa), .hikareru(_sub_plot_x_123_hikareru), .moto(_sub_plot_x_123_moto));
sub_plot sub_plot_x_122 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_122_in_do), .sa(_sub_plot_x_122_sa), .hikareru(_sub_plot_x_122_hikareru), .moto(_sub_plot_x_122_moto));
sub_plot sub_plot_x_121 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_121_in_do), .sa(_sub_plot_x_121_sa), .hikareru(_sub_plot_x_121_hikareru), .moto(_sub_plot_x_121_moto));
sub_plot sub_plot_x_120 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_120_in_do), .sa(_sub_plot_x_120_sa), .hikareru(_sub_plot_x_120_hikareru), .moto(_sub_plot_x_120_moto));
sub_plot sub_plot_x_119 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_119_in_do), .sa(_sub_plot_x_119_sa), .hikareru(_sub_plot_x_119_hikareru), .moto(_sub_plot_x_119_moto));
sub_plot sub_plot_x_118 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_118_in_do), .sa(_sub_plot_x_118_sa), .hikareru(_sub_plot_x_118_hikareru), .moto(_sub_plot_x_118_moto));
sub_plot sub_plot_x_117 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_117_in_do), .sa(_sub_plot_x_117_sa), .hikareru(_sub_plot_x_117_hikareru), .moto(_sub_plot_x_117_moto));
sub_plot sub_plot_x_116 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_116_in_do), .sa(_sub_plot_x_116_sa), .hikareru(_sub_plot_x_116_hikareru), .moto(_sub_plot_x_116_moto));
sub_plot sub_plot_x_115 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_115_in_do), .sa(_sub_plot_x_115_sa), .hikareru(_sub_plot_x_115_hikareru), .moto(_sub_plot_x_115_moto));
sub_plot sub_plot_x_114 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_114_in_do), .sa(_sub_plot_x_114_sa), .hikareru(_sub_plot_x_114_hikareru), .moto(_sub_plot_x_114_moto));
sub_plot sub_plot_x_113 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_113_in_do), .sa(_sub_plot_x_113_sa), .hikareru(_sub_plot_x_113_hikareru), .moto(_sub_plot_x_113_moto));
sub_plot sub_plot_x_112 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_112_in_do), .sa(_sub_plot_x_112_sa), .hikareru(_sub_plot_x_112_hikareru), .moto(_sub_plot_x_112_moto));
sub_plot sub_plot_x_111 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_111_in_do), .sa(_sub_plot_x_111_sa), .hikareru(_sub_plot_x_111_hikareru), .moto(_sub_plot_x_111_moto));
sub_plot sub_plot_x_110 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_110_in_do), .sa(_sub_plot_x_110_sa), .hikareru(_sub_plot_x_110_hikareru), .moto(_sub_plot_x_110_moto));
sub_plot sub_plot_x_109 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_109_in_do), .sa(_sub_plot_x_109_sa), .hikareru(_sub_plot_x_109_hikareru), .moto(_sub_plot_x_109_moto));
sub_plot sub_plot_x_108 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_108_in_do), .sa(_sub_plot_x_108_sa), .hikareru(_sub_plot_x_108_hikareru), .moto(_sub_plot_x_108_moto));
sub_plot sub_plot_x_107 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_107_in_do), .sa(_sub_plot_x_107_sa), .hikareru(_sub_plot_x_107_hikareru), .moto(_sub_plot_x_107_moto));
sub_plot sub_plot_x_106 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_106_in_do), .sa(_sub_plot_x_106_sa), .hikareru(_sub_plot_x_106_hikareru), .moto(_sub_plot_x_106_moto));
sub_plot sub_plot_x_105 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_105_in_do), .sa(_sub_plot_x_105_sa), .hikareru(_sub_plot_x_105_hikareru), .moto(_sub_plot_x_105_moto));
sub_plot sub_plot_x_104 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_104_in_do), .sa(_sub_plot_x_104_sa), .hikareru(_sub_plot_x_104_hikareru), .moto(_sub_plot_x_104_moto));
sub_plot sub_plot_x_103 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_103_in_do), .sa(_sub_plot_x_103_sa), .hikareru(_sub_plot_x_103_hikareru), .moto(_sub_plot_x_103_moto));
sub_plot sub_plot_x_102 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_102_in_do), .sa(_sub_plot_x_102_sa), .hikareru(_sub_plot_x_102_hikareru), .moto(_sub_plot_x_102_moto));
sub_plot sub_plot_x_101 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_101_in_do), .sa(_sub_plot_x_101_sa), .hikareru(_sub_plot_x_101_hikareru), .moto(_sub_plot_x_101_moto));
sub_plot sub_plot_x_100 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_100_in_do), .sa(_sub_plot_x_100_sa), .hikareru(_sub_plot_x_100_hikareru), .moto(_sub_plot_x_100_moto));
sub_plot sub_plot_x_99 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_99_in_do), .sa(_sub_plot_x_99_sa), .hikareru(_sub_plot_x_99_hikareru), .moto(_sub_plot_x_99_moto));
sub_plot sub_plot_x_98 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_98_in_do), .sa(_sub_plot_x_98_sa), .hikareru(_sub_plot_x_98_hikareru), .moto(_sub_plot_x_98_moto));
sub_plot sub_plot_x_97 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_97_in_do), .sa(_sub_plot_x_97_sa), .hikareru(_sub_plot_x_97_hikareru), .moto(_sub_plot_x_97_moto));
sub_plot sub_plot_x_96 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_96_in_do), .sa(_sub_plot_x_96_sa), .hikareru(_sub_plot_x_96_hikareru), .moto(_sub_plot_x_96_moto));
sub_plot sub_plot_x_95 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_95_in_do), .sa(_sub_plot_x_95_sa), .hikareru(_sub_plot_x_95_hikareru), .moto(_sub_plot_x_95_moto));
sub_plot sub_plot_x_94 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_94_in_do), .sa(_sub_plot_x_94_sa), .hikareru(_sub_plot_x_94_hikareru), .moto(_sub_plot_x_94_moto));
sub_plot sub_plot_x_93 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_93_in_do), .sa(_sub_plot_x_93_sa), .hikareru(_sub_plot_x_93_hikareru), .moto(_sub_plot_x_93_moto));
sub_plot sub_plot_x_92 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_92_in_do), .sa(_sub_plot_x_92_sa), .hikareru(_sub_plot_x_92_hikareru), .moto(_sub_plot_x_92_moto));
sub_plot sub_plot_x_91 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_91_in_do), .sa(_sub_plot_x_91_sa), .hikareru(_sub_plot_x_91_hikareru), .moto(_sub_plot_x_91_moto));
sub_plot sub_plot_x_90 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_90_in_do), .sa(_sub_plot_x_90_sa), .hikareru(_sub_plot_x_90_hikareru), .moto(_sub_plot_x_90_moto));
sub_plot sub_plot_x_89 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_89_in_do), .sa(_sub_plot_x_89_sa), .hikareru(_sub_plot_x_89_hikareru), .moto(_sub_plot_x_89_moto));
sub_plot sub_plot_x_88 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_88_in_do), .sa(_sub_plot_x_88_sa), .hikareru(_sub_plot_x_88_hikareru), .moto(_sub_plot_x_88_moto));
sub_plot sub_plot_x_87 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_87_in_do), .sa(_sub_plot_x_87_sa), .hikareru(_sub_plot_x_87_hikareru), .moto(_sub_plot_x_87_moto));
sub_plot sub_plot_x_86 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_86_in_do), .sa(_sub_plot_x_86_sa), .hikareru(_sub_plot_x_86_hikareru), .moto(_sub_plot_x_86_moto));
sub_plot sub_plot_x_85 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_85_in_do), .sa(_sub_plot_x_85_sa), .hikareru(_sub_plot_x_85_hikareru), .moto(_sub_plot_x_85_moto));
sub_plot sub_plot_x_84 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_84_in_do), .sa(_sub_plot_x_84_sa), .hikareru(_sub_plot_x_84_hikareru), .moto(_sub_plot_x_84_moto));
sub_plot sub_plot_x_83 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_83_in_do), .sa(_sub_plot_x_83_sa), .hikareru(_sub_plot_x_83_hikareru), .moto(_sub_plot_x_83_moto));
sub_plot sub_plot_x_82 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_82_in_do), .sa(_sub_plot_x_82_sa), .hikareru(_sub_plot_x_82_hikareru), .moto(_sub_plot_x_82_moto));
sub_plot sub_plot_x_81 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_81_in_do), .sa(_sub_plot_x_81_sa), .hikareru(_sub_plot_x_81_hikareru), .moto(_sub_plot_x_81_moto));
sub_plot sub_plot_x_80 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_80_in_do), .sa(_sub_plot_x_80_sa), .hikareru(_sub_plot_x_80_hikareru), .moto(_sub_plot_x_80_moto));
sub_plot sub_plot_x_79 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_79_in_do), .sa(_sub_plot_x_79_sa), .hikareru(_sub_plot_x_79_hikareru), .moto(_sub_plot_x_79_moto));
sub_plot sub_plot_x_78 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_78_in_do), .sa(_sub_plot_x_78_sa), .hikareru(_sub_plot_x_78_hikareru), .moto(_sub_plot_x_78_moto));
sub_plot sub_plot_x_77 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_77_in_do), .sa(_sub_plot_x_77_sa), .hikareru(_sub_plot_x_77_hikareru), .moto(_sub_plot_x_77_moto));
sub_plot sub_plot_x_76 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_76_in_do), .sa(_sub_plot_x_76_sa), .hikareru(_sub_plot_x_76_hikareru), .moto(_sub_plot_x_76_moto));
sub_plot sub_plot_x_75 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_75_in_do), .sa(_sub_plot_x_75_sa), .hikareru(_sub_plot_x_75_hikareru), .moto(_sub_plot_x_75_moto));
sub_plot sub_plot_x_74 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_74_in_do), .sa(_sub_plot_x_74_sa), .hikareru(_sub_plot_x_74_hikareru), .moto(_sub_plot_x_74_moto));
sub_plot sub_plot_x_73 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_73_in_do), .sa(_sub_plot_x_73_sa), .hikareru(_sub_plot_x_73_hikareru), .moto(_sub_plot_x_73_moto));
sub_plot sub_plot_x_72 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_72_in_do), .sa(_sub_plot_x_72_sa), .hikareru(_sub_plot_x_72_hikareru), .moto(_sub_plot_x_72_moto));
sub_plot sub_plot_x_71 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_71_in_do), .sa(_sub_plot_x_71_sa), .hikareru(_sub_plot_x_71_hikareru), .moto(_sub_plot_x_71_moto));
sub_plot sub_plot_x_70 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_70_in_do), .sa(_sub_plot_x_70_sa), .hikareru(_sub_plot_x_70_hikareru), .moto(_sub_plot_x_70_moto));
sub_plot sub_plot_x_69 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_69_in_do), .sa(_sub_plot_x_69_sa), .hikareru(_sub_plot_x_69_hikareru), .moto(_sub_plot_x_69_moto));
sub_plot sub_plot_x_68 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_68_in_do), .sa(_sub_plot_x_68_sa), .hikareru(_sub_plot_x_68_hikareru), .moto(_sub_plot_x_68_moto));
sub_plot sub_plot_x_67 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_67_in_do), .sa(_sub_plot_x_67_sa), .hikareru(_sub_plot_x_67_hikareru), .moto(_sub_plot_x_67_moto));
sub_plot sub_plot_x_66 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_66_in_do), .sa(_sub_plot_x_66_sa), .hikareru(_sub_plot_x_66_hikareru), .moto(_sub_plot_x_66_moto));
sub_plot sub_plot_x_65 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_65_in_do), .sa(_sub_plot_x_65_sa), .hikareru(_sub_plot_x_65_hikareru), .moto(_sub_plot_x_65_moto));
sub_plot sub_plot_x_64 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_64_in_do), .sa(_sub_plot_x_64_sa), .hikareru(_sub_plot_x_64_hikareru), .moto(_sub_plot_x_64_moto));
sub_plot sub_plot_x_63 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_63_in_do), .sa(_sub_plot_x_63_sa), .hikareru(_sub_plot_x_63_hikareru), .moto(_sub_plot_x_63_moto));
sub_plot sub_plot_x_62 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_62_in_do), .sa(_sub_plot_x_62_sa), .hikareru(_sub_plot_x_62_hikareru), .moto(_sub_plot_x_62_moto));
sub_plot sub_plot_x_61 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_61_in_do), .sa(_sub_plot_x_61_sa), .hikareru(_sub_plot_x_61_hikareru), .moto(_sub_plot_x_61_moto));
sub_plot sub_plot_x_60 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_60_in_do), .sa(_sub_plot_x_60_sa), .hikareru(_sub_plot_x_60_hikareru), .moto(_sub_plot_x_60_moto));
sub_plot sub_plot_x_59 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_59_in_do), .sa(_sub_plot_x_59_sa), .hikareru(_sub_plot_x_59_hikareru), .moto(_sub_plot_x_59_moto));
sub_plot sub_plot_x_58 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_58_in_do), .sa(_sub_plot_x_58_sa), .hikareru(_sub_plot_x_58_hikareru), .moto(_sub_plot_x_58_moto));
sub_plot sub_plot_x_57 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_57_in_do), .sa(_sub_plot_x_57_sa), .hikareru(_sub_plot_x_57_hikareru), .moto(_sub_plot_x_57_moto));
sub_plot sub_plot_x_56 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_56_in_do), .sa(_sub_plot_x_56_sa), .hikareru(_sub_plot_x_56_hikareru), .moto(_sub_plot_x_56_moto));
sub_plot sub_plot_x_55 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_55_in_do), .sa(_sub_plot_x_55_sa), .hikareru(_sub_plot_x_55_hikareru), .moto(_sub_plot_x_55_moto));
sub_plot sub_plot_x_54 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_54_in_do), .sa(_sub_plot_x_54_sa), .hikareru(_sub_plot_x_54_hikareru), .moto(_sub_plot_x_54_moto));
sub_plot sub_plot_x_53 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_53_in_do), .sa(_sub_plot_x_53_sa), .hikareru(_sub_plot_x_53_hikareru), .moto(_sub_plot_x_53_moto));
sub_plot sub_plot_x_52 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_52_in_do), .sa(_sub_plot_x_52_sa), .hikareru(_sub_plot_x_52_hikareru), .moto(_sub_plot_x_52_moto));
sub_plot sub_plot_x_51 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_51_in_do), .sa(_sub_plot_x_51_sa), .hikareru(_sub_plot_x_51_hikareru), .moto(_sub_plot_x_51_moto));
sub_plot sub_plot_x_50 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_50_in_do), .sa(_sub_plot_x_50_sa), .hikareru(_sub_plot_x_50_hikareru), .moto(_sub_plot_x_50_moto));
sub_plot sub_plot_x_49 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_49_in_do), .sa(_sub_plot_x_49_sa), .hikareru(_sub_plot_x_49_hikareru), .moto(_sub_plot_x_49_moto));
sub_plot sub_plot_x_48 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_48_in_do), .sa(_sub_plot_x_48_sa), .hikareru(_sub_plot_x_48_hikareru), .moto(_sub_plot_x_48_moto));
sub_plot sub_plot_x_47 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_47_in_do), .sa(_sub_plot_x_47_sa), .hikareru(_sub_plot_x_47_hikareru), .moto(_sub_plot_x_47_moto));
sub_plot sub_plot_x_46 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_46_in_do), .sa(_sub_plot_x_46_sa), .hikareru(_sub_plot_x_46_hikareru), .moto(_sub_plot_x_46_moto));
sub_plot sub_plot_x_45 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_45_in_do), .sa(_sub_plot_x_45_sa), .hikareru(_sub_plot_x_45_hikareru), .moto(_sub_plot_x_45_moto));
sub_plot sub_plot_x_44 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_44_in_do), .sa(_sub_plot_x_44_sa), .hikareru(_sub_plot_x_44_hikareru), .moto(_sub_plot_x_44_moto));
sub_plot sub_plot_x_43 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_43_in_do), .sa(_sub_plot_x_43_sa), .hikareru(_sub_plot_x_43_hikareru), .moto(_sub_plot_x_43_moto));
sub_plot sub_plot_x_42 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_42_in_do), .sa(_sub_plot_x_42_sa), .hikareru(_sub_plot_x_42_hikareru), .moto(_sub_plot_x_42_moto));
sub_plot sub_plot_x_41 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_41_in_do), .sa(_sub_plot_x_41_sa), .hikareru(_sub_plot_x_41_hikareru), .moto(_sub_plot_x_41_moto));
sub_plot sub_plot_x_40 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_40_in_do), .sa(_sub_plot_x_40_sa), .hikareru(_sub_plot_x_40_hikareru), .moto(_sub_plot_x_40_moto));
sub_plot sub_plot_x_39 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_39_in_do), .sa(_sub_plot_x_39_sa), .hikareru(_sub_plot_x_39_hikareru), .moto(_sub_plot_x_39_moto));
sub_plot sub_plot_x_38 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_38_in_do), .sa(_sub_plot_x_38_sa), .hikareru(_sub_plot_x_38_hikareru), .moto(_sub_plot_x_38_moto));
sub_plot sub_plot_x_37 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_37_in_do), .sa(_sub_plot_x_37_sa), .hikareru(_sub_plot_x_37_hikareru), .moto(_sub_plot_x_37_moto));
sub_plot sub_plot_x_36 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_36_in_do), .sa(_sub_plot_x_36_sa), .hikareru(_sub_plot_x_36_hikareru), .moto(_sub_plot_x_36_moto));
sub_plot sub_plot_x_35 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_35_in_do), .sa(_sub_plot_x_35_sa), .hikareru(_sub_plot_x_35_hikareru), .moto(_sub_plot_x_35_moto));
sub_plot sub_plot_x_34 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_34_in_do), .sa(_sub_plot_x_34_sa), .hikareru(_sub_plot_x_34_hikareru), .moto(_sub_plot_x_34_moto));
sub_plot sub_plot_x_33 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_33_in_do), .sa(_sub_plot_x_33_sa), .hikareru(_sub_plot_x_33_hikareru), .moto(_sub_plot_x_33_moto));
sub_plot sub_plot_x_32 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_32_in_do), .sa(_sub_plot_x_32_sa), .hikareru(_sub_plot_x_32_hikareru), .moto(_sub_plot_x_32_moto));
sub_plot sub_plot_x_31 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_31_in_do), .sa(_sub_plot_x_31_sa), .hikareru(_sub_plot_x_31_hikareru), .moto(_sub_plot_x_31_moto));
sub_plot sub_plot_x_30 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_30_in_do), .sa(_sub_plot_x_30_sa), .hikareru(_sub_plot_x_30_hikareru), .moto(_sub_plot_x_30_moto));
sub_plot sub_plot_x_29 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_29_in_do), .sa(_sub_plot_x_29_sa), .hikareru(_sub_plot_x_29_hikareru), .moto(_sub_plot_x_29_moto));
sub_plot sub_plot_x_28 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_28_in_do), .sa(_sub_plot_x_28_sa), .hikareru(_sub_plot_x_28_hikareru), .moto(_sub_plot_x_28_moto));
sub_plot sub_plot_x_27 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_27_in_do), .sa(_sub_plot_x_27_sa), .hikareru(_sub_plot_x_27_hikareru), .moto(_sub_plot_x_27_moto));
sub_plot sub_plot_x_26 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_26_in_do), .sa(_sub_plot_x_26_sa), .hikareru(_sub_plot_x_26_hikareru), .moto(_sub_plot_x_26_moto));
sub_plot sub_plot_x_25 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_25_in_do), .sa(_sub_plot_x_25_sa), .hikareru(_sub_plot_x_25_hikareru), .moto(_sub_plot_x_25_moto));
sub_plot sub_plot_x_24 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_24_in_do), .sa(_sub_plot_x_24_sa), .hikareru(_sub_plot_x_24_hikareru), .moto(_sub_plot_x_24_moto));
sub_plot sub_plot_x_23 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_23_in_do), .sa(_sub_plot_x_23_sa), .hikareru(_sub_plot_x_23_hikareru), .moto(_sub_plot_x_23_moto));
sub_plot sub_plot_x_22 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_22_in_do), .sa(_sub_plot_x_22_sa), .hikareru(_sub_plot_x_22_hikareru), .moto(_sub_plot_x_22_moto));
sub_plot sub_plot_x_21 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_21_in_do), .sa(_sub_plot_x_21_sa), .hikareru(_sub_plot_x_21_hikareru), .moto(_sub_plot_x_21_moto));
sub_plot sub_plot_x_20 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_20_in_do), .sa(_sub_plot_x_20_sa), .hikareru(_sub_plot_x_20_hikareru), .moto(_sub_plot_x_20_moto));
sub_plot sub_plot_x_19 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_19_in_do), .sa(_sub_plot_x_19_sa), .hikareru(_sub_plot_x_19_hikareru), .moto(_sub_plot_x_19_moto));
sub_plot sub_plot_x_18 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_18_in_do), .sa(_sub_plot_x_18_sa), .hikareru(_sub_plot_x_18_hikareru), .moto(_sub_plot_x_18_moto));
sub_plot sub_plot_x_17 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_17_in_do), .sa(_sub_plot_x_17_sa), .hikareru(_sub_plot_x_17_hikareru), .moto(_sub_plot_x_17_moto));
sub_plot sub_plot_x_16 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_16_in_do), .sa(_sub_plot_x_16_sa), .hikareru(_sub_plot_x_16_hikareru), .moto(_sub_plot_x_16_moto));
sub_plot sub_plot_x_15 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_15_in_do), .sa(_sub_plot_x_15_sa), .hikareru(_sub_plot_x_15_hikareru), .moto(_sub_plot_x_15_moto));
sub_plot sub_plot_x_14 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_14_in_do), .sa(_sub_plot_x_14_sa), .hikareru(_sub_plot_x_14_hikareru), .moto(_sub_plot_x_14_moto));
sub_plot sub_plot_x_13 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_13_in_do), .sa(_sub_plot_x_13_sa), .hikareru(_sub_plot_x_13_hikareru), .moto(_sub_plot_x_13_moto));
sub_plot sub_plot_x_12 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_12_in_do), .sa(_sub_plot_x_12_sa), .hikareru(_sub_plot_x_12_hikareru), .moto(_sub_plot_x_12_moto));
sub_plot sub_plot_x_11 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_11_in_do), .sa(_sub_plot_x_11_sa), .hikareru(_sub_plot_x_11_hikareru), .moto(_sub_plot_x_11_moto));
sub_plot sub_plot_x_10 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_10_in_do), .sa(_sub_plot_x_10_sa), .hikareru(_sub_plot_x_10_hikareru), .moto(_sub_plot_x_10_moto));
sub_plot sub_plot_x_9 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_9_in_do), .sa(_sub_plot_x_9_sa), .hikareru(_sub_plot_x_9_hikareru), .moto(_sub_plot_x_9_moto));
sub_plot sub_plot_x_8 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_8_in_do), .sa(_sub_plot_x_8_sa), .hikareru(_sub_plot_x_8_hikareru), .moto(_sub_plot_x_8_moto));
sub_plot sub_plot_x_7 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_7_in_do), .sa(_sub_plot_x_7_sa), .hikareru(_sub_plot_x_7_hikareru), .moto(_sub_plot_x_7_moto));
sub_plot sub_plot_x_6 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_6_in_do), .sa(_sub_plot_x_6_sa), .hikareru(_sub_plot_x_6_hikareru), .moto(_sub_plot_x_6_moto));
sub_plot sub_plot_x_5 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_5_in_do), .sa(_sub_plot_x_5_sa), .hikareru(_sub_plot_x_5_hikareru), .moto(_sub_plot_x_5_moto));
sub_plot sub_plot_x_4 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_4_in_do), .sa(_sub_plot_x_4_sa), .hikareru(_sub_plot_x_4_hikareru), .moto(_sub_plot_x_4_moto));
sub_plot sub_plot_x_3 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_3_in_do), .sa(_sub_plot_x_3_sa), .hikareru(_sub_plot_x_3_hikareru), .moto(_sub_plot_x_3_moto));
sub_plot sub_plot_x_2 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_2_in_do), .sa(_sub_plot_x_2_sa), .hikareru(_sub_plot_x_2_hikareru), .moto(_sub_plot_x_2_moto));
sub_plot sub_plot_x_1 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_sub_plot_x_1_in_do), .sa(_sub_plot_x_1_sa), .hikareru(_sub_plot_x_1_hikareru), .moto(_sub_plot_x_1_moto));

   assign  _sub_plot_x_hikareru = data_in33;
   assign  _sub_plot_x_moto = data_in_index33;
   assign  _sub_plot_x_in_do = subs_exe;
   assign  _sub_plot_x_p_reset = p_reset;
   assign  _sub_plot_x_m_clock = m_clock;
   assign  _sub_plot_x_209_hikareru = data_in477;
   assign  _sub_plot_x_209_moto = data_in_index477;
   assign  _sub_plot_x_209_in_do = subs_exe;
   assign  _sub_plot_x_209_p_reset = p_reset;
   assign  _sub_plot_x_209_m_clock = m_clock;
   assign  _sub_plot_x_208_hikareru = data_in475;
   assign  _sub_plot_x_208_moto = data_in_index475;
   assign  _sub_plot_x_208_in_do = subs_exe;
   assign  _sub_plot_x_208_p_reset = p_reset;
   assign  _sub_plot_x_208_m_clock = m_clock;
   assign  _sub_plot_x_207_hikareru = data_in473;
   assign  _sub_plot_x_207_moto = data_in_index473;
   assign  _sub_plot_x_207_in_do = subs_exe;
   assign  _sub_plot_x_207_p_reset = p_reset;
   assign  _sub_plot_x_207_m_clock = m_clock;
   assign  _sub_plot_x_206_hikareru = data_in471;
   assign  _sub_plot_x_206_moto = data_in_index471;
   assign  _sub_plot_x_206_in_do = subs_exe;
   assign  _sub_plot_x_206_p_reset = p_reset;
   assign  _sub_plot_x_206_m_clock = m_clock;
   assign  _sub_plot_x_205_hikareru = data_in469;
   assign  _sub_plot_x_205_moto = data_in_index469;
   assign  _sub_plot_x_205_in_do = subs_exe;
   assign  _sub_plot_x_205_p_reset = p_reset;
   assign  _sub_plot_x_205_m_clock = m_clock;
   assign  _sub_plot_x_204_hikareru = data_in467;
   assign  _sub_plot_x_204_moto = data_in_index467;
   assign  _sub_plot_x_204_in_do = subs_exe;
   assign  _sub_plot_x_204_p_reset = p_reset;
   assign  _sub_plot_x_204_m_clock = m_clock;
   assign  _sub_plot_x_203_hikareru = data_in465;
   assign  _sub_plot_x_203_moto = data_in_index465;
   assign  _sub_plot_x_203_in_do = subs_exe;
   assign  _sub_plot_x_203_p_reset = p_reset;
   assign  _sub_plot_x_203_m_clock = m_clock;
   assign  _sub_plot_x_202_hikareru = data_in463;
   assign  _sub_plot_x_202_moto = data_in_index463;
   assign  _sub_plot_x_202_in_do = subs_exe;
   assign  _sub_plot_x_202_p_reset = p_reset;
   assign  _sub_plot_x_202_m_clock = m_clock;
   assign  _sub_plot_x_201_hikareru = data_in461;
   assign  _sub_plot_x_201_moto = data_in_index461;
   assign  _sub_plot_x_201_in_do = subs_exe;
   assign  _sub_plot_x_201_p_reset = p_reset;
   assign  _sub_plot_x_201_m_clock = m_clock;
   assign  _sub_plot_x_200_hikareru = data_in459;
   assign  _sub_plot_x_200_moto = data_in_index459;
   assign  _sub_plot_x_200_in_do = subs_exe;
   assign  _sub_plot_x_200_p_reset = p_reset;
   assign  _sub_plot_x_200_m_clock = m_clock;
   assign  _sub_plot_x_199_hikareru = data_in457;
   assign  _sub_plot_x_199_moto = data_in_index457;
   assign  _sub_plot_x_199_in_do = subs_exe;
   assign  _sub_plot_x_199_p_reset = p_reset;
   assign  _sub_plot_x_199_m_clock = m_clock;
   assign  _sub_plot_x_198_hikareru = data_in455;
   assign  _sub_plot_x_198_moto = data_in_index455;
   assign  _sub_plot_x_198_in_do = subs_exe;
   assign  _sub_plot_x_198_p_reset = p_reset;
   assign  _sub_plot_x_198_m_clock = m_clock;
   assign  _sub_plot_x_197_hikareru = data_in453;
   assign  _sub_plot_x_197_moto = data_in_index453;
   assign  _sub_plot_x_197_in_do = subs_exe;
   assign  _sub_plot_x_197_p_reset = p_reset;
   assign  _sub_plot_x_197_m_clock = m_clock;
   assign  _sub_plot_x_196_hikareru = data_in451;
   assign  _sub_plot_x_196_moto = data_in_index451;
   assign  _sub_plot_x_196_in_do = subs_exe;
   assign  _sub_plot_x_196_p_reset = p_reset;
   assign  _sub_plot_x_196_m_clock = m_clock;
   assign  _sub_plot_x_195_hikareru = data_in449;
   assign  _sub_plot_x_195_moto = data_in_index449;
   assign  _sub_plot_x_195_in_do = subs_exe;
   assign  _sub_plot_x_195_p_reset = p_reset;
   assign  _sub_plot_x_195_m_clock = m_clock;
   assign  _sub_plot_x_194_hikareru = data_in445;
   assign  _sub_plot_x_194_moto = data_in_index445;
   assign  _sub_plot_x_194_in_do = subs_exe;
   assign  _sub_plot_x_194_p_reset = p_reset;
   assign  _sub_plot_x_194_m_clock = m_clock;
   assign  _sub_plot_x_193_hikareru = data_in443;
   assign  _sub_plot_x_193_moto = data_in_index443;
   assign  _sub_plot_x_193_in_do = subs_exe;
   assign  _sub_plot_x_193_p_reset = p_reset;
   assign  _sub_plot_x_193_m_clock = m_clock;
   assign  _sub_plot_x_192_hikareru = data_in441;
   assign  _sub_plot_x_192_moto = data_in_index441;
   assign  _sub_plot_x_192_in_do = subs_exe;
   assign  _sub_plot_x_192_p_reset = p_reset;
   assign  _sub_plot_x_192_m_clock = m_clock;
   assign  _sub_plot_x_191_hikareru = data_in439;
   assign  _sub_plot_x_191_moto = data_in_index439;
   assign  _sub_plot_x_191_in_do = subs_exe;
   assign  _sub_plot_x_191_p_reset = p_reset;
   assign  _sub_plot_x_191_m_clock = m_clock;
   assign  _sub_plot_x_190_hikareru = data_in437;
   assign  _sub_plot_x_190_moto = data_in_index437;
   assign  _sub_plot_x_190_in_do = subs_exe;
   assign  _sub_plot_x_190_p_reset = p_reset;
   assign  _sub_plot_x_190_m_clock = m_clock;
   assign  _sub_plot_x_189_hikareru = data_in435;
   assign  _sub_plot_x_189_moto = data_in_index435;
   assign  _sub_plot_x_189_in_do = subs_exe;
   assign  _sub_plot_x_189_p_reset = p_reset;
   assign  _sub_plot_x_189_m_clock = m_clock;
   assign  _sub_plot_x_188_hikareru = data_in433;
   assign  _sub_plot_x_188_moto = data_in_index433;
   assign  _sub_plot_x_188_in_do = subs_exe;
   assign  _sub_plot_x_188_p_reset = p_reset;
   assign  _sub_plot_x_188_m_clock = m_clock;
   assign  _sub_plot_x_187_hikareru = data_in431;
   assign  _sub_plot_x_187_moto = data_in_index431;
   assign  _sub_plot_x_187_in_do = subs_exe;
   assign  _sub_plot_x_187_p_reset = p_reset;
   assign  _sub_plot_x_187_m_clock = m_clock;
   assign  _sub_plot_x_186_hikareru = data_in429;
   assign  _sub_plot_x_186_moto = data_in_index429;
   assign  _sub_plot_x_186_in_do = subs_exe;
   assign  _sub_plot_x_186_p_reset = p_reset;
   assign  _sub_plot_x_186_m_clock = m_clock;
   assign  _sub_plot_x_185_hikareru = data_in427;
   assign  _sub_plot_x_185_moto = data_in_index427;
   assign  _sub_plot_x_185_in_do = subs_exe;
   assign  _sub_plot_x_185_p_reset = p_reset;
   assign  _sub_plot_x_185_m_clock = m_clock;
   assign  _sub_plot_x_184_hikareru = data_in425;
   assign  _sub_plot_x_184_moto = data_in_index425;
   assign  _sub_plot_x_184_in_do = subs_exe;
   assign  _sub_plot_x_184_p_reset = p_reset;
   assign  _sub_plot_x_184_m_clock = m_clock;
   assign  _sub_plot_x_183_hikareru = data_in423;
   assign  _sub_plot_x_183_moto = data_in_index423;
   assign  _sub_plot_x_183_in_do = subs_exe;
   assign  _sub_plot_x_183_p_reset = p_reset;
   assign  _sub_plot_x_183_m_clock = m_clock;
   assign  _sub_plot_x_182_hikareru = data_in421;
   assign  _sub_plot_x_182_moto = data_in_index421;
   assign  _sub_plot_x_182_in_do = subs_exe;
   assign  _sub_plot_x_182_p_reset = p_reset;
   assign  _sub_plot_x_182_m_clock = m_clock;
   assign  _sub_plot_x_181_hikareru = data_in419;
   assign  _sub_plot_x_181_moto = data_in_index419;
   assign  _sub_plot_x_181_in_do = subs_exe;
   assign  _sub_plot_x_181_p_reset = p_reset;
   assign  _sub_plot_x_181_m_clock = m_clock;
   assign  _sub_plot_x_180_hikareru = data_in417;
   assign  _sub_plot_x_180_moto = data_in_index417;
   assign  _sub_plot_x_180_in_do = subs_exe;
   assign  _sub_plot_x_180_p_reset = p_reset;
   assign  _sub_plot_x_180_m_clock = m_clock;
   assign  _sub_plot_x_179_hikareru = data_in413;
   assign  _sub_plot_x_179_moto = data_in_index413;
   assign  _sub_plot_x_179_in_do = subs_exe;
   assign  _sub_plot_x_179_p_reset = p_reset;
   assign  _sub_plot_x_179_m_clock = m_clock;
   assign  _sub_plot_x_178_hikareru = data_in411;
   assign  _sub_plot_x_178_moto = data_in_index411;
   assign  _sub_plot_x_178_in_do = subs_exe;
   assign  _sub_plot_x_178_p_reset = p_reset;
   assign  _sub_plot_x_178_m_clock = m_clock;
   assign  _sub_plot_x_177_hikareru = data_in409;
   assign  _sub_plot_x_177_moto = data_in_index409;
   assign  _sub_plot_x_177_in_do = subs_exe;
   assign  _sub_plot_x_177_p_reset = p_reset;
   assign  _sub_plot_x_177_m_clock = m_clock;
   assign  _sub_plot_x_176_hikareru = data_in407;
   assign  _sub_plot_x_176_moto = data_in_index407;
   assign  _sub_plot_x_176_in_do = subs_exe;
   assign  _sub_plot_x_176_p_reset = p_reset;
   assign  _sub_plot_x_176_m_clock = m_clock;
   assign  _sub_plot_x_175_hikareru = data_in405;
   assign  _sub_plot_x_175_moto = data_in_index405;
   assign  _sub_plot_x_175_in_do = subs_exe;
   assign  _sub_plot_x_175_p_reset = p_reset;
   assign  _sub_plot_x_175_m_clock = m_clock;
   assign  _sub_plot_x_174_hikareru = data_in403;
   assign  _sub_plot_x_174_moto = data_in_index403;
   assign  _sub_plot_x_174_in_do = subs_exe;
   assign  _sub_plot_x_174_p_reset = p_reset;
   assign  _sub_plot_x_174_m_clock = m_clock;
   assign  _sub_plot_x_173_hikareru = data_in401;
   assign  _sub_plot_x_173_moto = data_in_index401;
   assign  _sub_plot_x_173_in_do = subs_exe;
   assign  _sub_plot_x_173_p_reset = p_reset;
   assign  _sub_plot_x_173_m_clock = m_clock;
   assign  _sub_plot_x_172_hikareru = data_in399;
   assign  _sub_plot_x_172_moto = data_in_index399;
   assign  _sub_plot_x_172_in_do = subs_exe;
   assign  _sub_plot_x_172_p_reset = p_reset;
   assign  _sub_plot_x_172_m_clock = m_clock;
   assign  _sub_plot_x_171_hikareru = data_in397;
   assign  _sub_plot_x_171_moto = data_in_index397;
   assign  _sub_plot_x_171_in_do = subs_exe;
   assign  _sub_plot_x_171_p_reset = p_reset;
   assign  _sub_plot_x_171_m_clock = m_clock;
   assign  _sub_plot_x_170_hikareru = data_in395;
   assign  _sub_plot_x_170_moto = data_in_index395;
   assign  _sub_plot_x_170_in_do = subs_exe;
   assign  _sub_plot_x_170_p_reset = p_reset;
   assign  _sub_plot_x_170_m_clock = m_clock;
   assign  _sub_plot_x_169_hikareru = data_in393;
   assign  _sub_plot_x_169_moto = data_in_index393;
   assign  _sub_plot_x_169_in_do = subs_exe;
   assign  _sub_plot_x_169_p_reset = p_reset;
   assign  _sub_plot_x_169_m_clock = m_clock;
   assign  _sub_plot_x_168_hikareru = data_in391;
   assign  _sub_plot_x_168_moto = data_in_index391;
   assign  _sub_plot_x_168_in_do = subs_exe;
   assign  _sub_plot_x_168_p_reset = p_reset;
   assign  _sub_plot_x_168_m_clock = m_clock;
   assign  _sub_plot_x_167_hikareru = data_in389;
   assign  _sub_plot_x_167_moto = data_in_index389;
   assign  _sub_plot_x_167_in_do = subs_exe;
   assign  _sub_plot_x_167_p_reset = p_reset;
   assign  _sub_plot_x_167_m_clock = m_clock;
   assign  _sub_plot_x_166_hikareru = data_in387;
   assign  _sub_plot_x_166_moto = data_in_index387;
   assign  _sub_plot_x_166_in_do = subs_exe;
   assign  _sub_plot_x_166_p_reset = p_reset;
   assign  _sub_plot_x_166_m_clock = m_clock;
   assign  _sub_plot_x_165_hikareru = data_in385;
   assign  _sub_plot_x_165_moto = data_in_index385;
   assign  _sub_plot_x_165_in_do = subs_exe;
   assign  _sub_plot_x_165_p_reset = p_reset;
   assign  _sub_plot_x_165_m_clock = m_clock;
   assign  _sub_plot_x_164_hikareru = data_in381;
   assign  _sub_plot_x_164_moto = data_in_index381;
   assign  _sub_plot_x_164_in_do = subs_exe;
   assign  _sub_plot_x_164_p_reset = p_reset;
   assign  _sub_plot_x_164_m_clock = m_clock;
   assign  _sub_plot_x_163_hikareru = data_in379;
   assign  _sub_plot_x_163_moto = data_in_index379;
   assign  _sub_plot_x_163_in_do = subs_exe;
   assign  _sub_plot_x_163_p_reset = p_reset;
   assign  _sub_plot_x_163_m_clock = m_clock;
   assign  _sub_plot_x_162_hikareru = data_in377;
   assign  _sub_plot_x_162_moto = data_in_index377;
   assign  _sub_plot_x_162_in_do = subs_exe;
   assign  _sub_plot_x_162_p_reset = p_reset;
   assign  _sub_plot_x_162_m_clock = m_clock;
   assign  _sub_plot_x_161_hikareru = data_in375;
   assign  _sub_plot_x_161_moto = data_in_index375;
   assign  _sub_plot_x_161_in_do = subs_exe;
   assign  _sub_plot_x_161_p_reset = p_reset;
   assign  _sub_plot_x_161_m_clock = m_clock;
   assign  _sub_plot_x_160_hikareru = data_in373;
   assign  _sub_plot_x_160_moto = data_in_index373;
   assign  _sub_plot_x_160_in_do = subs_exe;
   assign  _sub_plot_x_160_p_reset = p_reset;
   assign  _sub_plot_x_160_m_clock = m_clock;
   assign  _sub_plot_x_159_hikareru = data_in371;
   assign  _sub_plot_x_159_moto = data_in_index371;
   assign  _sub_plot_x_159_in_do = subs_exe;
   assign  _sub_plot_x_159_p_reset = p_reset;
   assign  _sub_plot_x_159_m_clock = m_clock;
   assign  _sub_plot_x_158_hikareru = data_in369;
   assign  _sub_plot_x_158_moto = data_in_index369;
   assign  _sub_plot_x_158_in_do = subs_exe;
   assign  _sub_plot_x_158_p_reset = p_reset;
   assign  _sub_plot_x_158_m_clock = m_clock;
   assign  _sub_plot_x_157_hikareru = data_in367;
   assign  _sub_plot_x_157_moto = data_in_index367;
   assign  _sub_plot_x_157_in_do = subs_exe;
   assign  _sub_plot_x_157_p_reset = p_reset;
   assign  _sub_plot_x_157_m_clock = m_clock;
   assign  _sub_plot_x_156_hikareru = data_in365;
   assign  _sub_plot_x_156_moto = data_in_index365;
   assign  _sub_plot_x_156_in_do = subs_exe;
   assign  _sub_plot_x_156_p_reset = p_reset;
   assign  _sub_plot_x_156_m_clock = m_clock;
   assign  _sub_plot_x_155_hikareru = data_in363;
   assign  _sub_plot_x_155_moto = data_in_index363;
   assign  _sub_plot_x_155_in_do = subs_exe;
   assign  _sub_plot_x_155_p_reset = p_reset;
   assign  _sub_plot_x_155_m_clock = m_clock;
   assign  _sub_plot_x_154_hikareru = data_in361;
   assign  _sub_plot_x_154_moto = data_in_index361;
   assign  _sub_plot_x_154_in_do = subs_exe;
   assign  _sub_plot_x_154_p_reset = p_reset;
   assign  _sub_plot_x_154_m_clock = m_clock;
   assign  _sub_plot_x_153_hikareru = data_in359;
   assign  _sub_plot_x_153_moto = data_in_index359;
   assign  _sub_plot_x_153_in_do = subs_exe;
   assign  _sub_plot_x_153_p_reset = p_reset;
   assign  _sub_plot_x_153_m_clock = m_clock;
   assign  _sub_plot_x_152_hikareru = data_in357;
   assign  _sub_plot_x_152_moto = data_in_index357;
   assign  _sub_plot_x_152_in_do = subs_exe;
   assign  _sub_plot_x_152_p_reset = p_reset;
   assign  _sub_plot_x_152_m_clock = m_clock;
   assign  _sub_plot_x_151_hikareru = data_in355;
   assign  _sub_plot_x_151_moto = data_in_index355;
   assign  _sub_plot_x_151_in_do = subs_exe;
   assign  _sub_plot_x_151_p_reset = p_reset;
   assign  _sub_plot_x_151_m_clock = m_clock;
   assign  _sub_plot_x_150_hikareru = data_in353;
   assign  _sub_plot_x_150_moto = data_in_index353;
   assign  _sub_plot_x_150_in_do = subs_exe;
   assign  _sub_plot_x_150_p_reset = p_reset;
   assign  _sub_plot_x_150_m_clock = m_clock;
   assign  _sub_plot_x_149_hikareru = data_in349;
   assign  _sub_plot_x_149_moto = data_in_index349;
   assign  _sub_plot_x_149_in_do = subs_exe;
   assign  _sub_plot_x_149_p_reset = p_reset;
   assign  _sub_plot_x_149_m_clock = m_clock;
   assign  _sub_plot_x_148_hikareru = data_in347;
   assign  _sub_plot_x_148_moto = data_in_index347;
   assign  _sub_plot_x_148_in_do = subs_exe;
   assign  _sub_plot_x_148_p_reset = p_reset;
   assign  _sub_plot_x_148_m_clock = m_clock;
   assign  _sub_plot_x_147_hikareru = data_in345;
   assign  _sub_plot_x_147_moto = data_in_index345;
   assign  _sub_plot_x_147_in_do = subs_exe;
   assign  _sub_plot_x_147_p_reset = p_reset;
   assign  _sub_plot_x_147_m_clock = m_clock;
   assign  _sub_plot_x_146_hikareru = data_in343;
   assign  _sub_plot_x_146_moto = data_in_index343;
   assign  _sub_plot_x_146_in_do = subs_exe;
   assign  _sub_plot_x_146_p_reset = p_reset;
   assign  _sub_plot_x_146_m_clock = m_clock;
   assign  _sub_plot_x_145_hikareru = data_in341;
   assign  _sub_plot_x_145_moto = data_in_index341;
   assign  _sub_plot_x_145_in_do = subs_exe;
   assign  _sub_plot_x_145_p_reset = p_reset;
   assign  _sub_plot_x_145_m_clock = m_clock;
   assign  _sub_plot_x_144_hikareru = data_in339;
   assign  _sub_plot_x_144_moto = data_in_index339;
   assign  _sub_plot_x_144_in_do = subs_exe;
   assign  _sub_plot_x_144_p_reset = p_reset;
   assign  _sub_plot_x_144_m_clock = m_clock;
   assign  _sub_plot_x_143_hikareru = data_in337;
   assign  _sub_plot_x_143_moto = data_in_index337;
   assign  _sub_plot_x_143_in_do = subs_exe;
   assign  _sub_plot_x_143_p_reset = p_reset;
   assign  _sub_plot_x_143_m_clock = m_clock;
   assign  _sub_plot_x_142_hikareru = data_in335;
   assign  _sub_plot_x_142_moto = data_in_index335;
   assign  _sub_plot_x_142_in_do = subs_exe;
   assign  _sub_plot_x_142_p_reset = p_reset;
   assign  _sub_plot_x_142_m_clock = m_clock;
   assign  _sub_plot_x_141_hikareru = data_in333;
   assign  _sub_plot_x_141_moto = data_in_index333;
   assign  _sub_plot_x_141_in_do = subs_exe;
   assign  _sub_plot_x_141_p_reset = p_reset;
   assign  _sub_plot_x_141_m_clock = m_clock;
   assign  _sub_plot_x_140_hikareru = data_in331;
   assign  _sub_plot_x_140_moto = data_in_index331;
   assign  _sub_plot_x_140_in_do = subs_exe;
   assign  _sub_plot_x_140_p_reset = p_reset;
   assign  _sub_plot_x_140_m_clock = m_clock;
   assign  _sub_plot_x_139_hikareru = data_in329;
   assign  _sub_plot_x_139_moto = data_in_index329;
   assign  _sub_plot_x_139_in_do = subs_exe;
   assign  _sub_plot_x_139_p_reset = p_reset;
   assign  _sub_plot_x_139_m_clock = m_clock;
   assign  _sub_plot_x_138_hikareru = data_in327;
   assign  _sub_plot_x_138_moto = data_in_index327;
   assign  _sub_plot_x_138_in_do = subs_exe;
   assign  _sub_plot_x_138_p_reset = p_reset;
   assign  _sub_plot_x_138_m_clock = m_clock;
   assign  _sub_plot_x_137_hikareru = data_in325;
   assign  _sub_plot_x_137_moto = data_in_index325;
   assign  _sub_plot_x_137_in_do = subs_exe;
   assign  _sub_plot_x_137_p_reset = p_reset;
   assign  _sub_plot_x_137_m_clock = m_clock;
   assign  _sub_plot_x_136_hikareru = data_in323;
   assign  _sub_plot_x_136_moto = data_in_index323;
   assign  _sub_plot_x_136_in_do = subs_exe;
   assign  _sub_plot_x_136_p_reset = p_reset;
   assign  _sub_plot_x_136_m_clock = m_clock;
   assign  _sub_plot_x_135_hikareru = data_in321;
   assign  _sub_plot_x_135_moto = data_in_index321;
   assign  _sub_plot_x_135_in_do = subs_exe;
   assign  _sub_plot_x_135_p_reset = p_reset;
   assign  _sub_plot_x_135_m_clock = m_clock;
   assign  _sub_plot_x_134_hikareru = data_in317;
   assign  _sub_plot_x_134_moto = data_in_index317;
   assign  _sub_plot_x_134_in_do = subs_exe;
   assign  _sub_plot_x_134_p_reset = p_reset;
   assign  _sub_plot_x_134_m_clock = m_clock;
   assign  _sub_plot_x_133_hikareru = data_in315;
   assign  _sub_plot_x_133_moto = data_in_index315;
   assign  _sub_plot_x_133_in_do = subs_exe;
   assign  _sub_plot_x_133_p_reset = p_reset;
   assign  _sub_plot_x_133_m_clock = m_clock;
   assign  _sub_plot_x_132_hikareru = data_in313;
   assign  _sub_plot_x_132_moto = data_in_index313;
   assign  _sub_plot_x_132_in_do = subs_exe;
   assign  _sub_plot_x_132_p_reset = p_reset;
   assign  _sub_plot_x_132_m_clock = m_clock;
   assign  _sub_plot_x_131_hikareru = data_in311;
   assign  _sub_plot_x_131_moto = data_in_index311;
   assign  _sub_plot_x_131_in_do = subs_exe;
   assign  _sub_plot_x_131_p_reset = p_reset;
   assign  _sub_plot_x_131_m_clock = m_clock;
   assign  _sub_plot_x_130_hikareru = data_in309;
   assign  _sub_plot_x_130_moto = data_in_index309;
   assign  _sub_plot_x_130_in_do = subs_exe;
   assign  _sub_plot_x_130_p_reset = p_reset;
   assign  _sub_plot_x_130_m_clock = m_clock;
   assign  _sub_plot_x_129_hikareru = data_in307;
   assign  _sub_plot_x_129_moto = data_in_index307;
   assign  _sub_plot_x_129_in_do = subs_exe;
   assign  _sub_plot_x_129_p_reset = p_reset;
   assign  _sub_plot_x_129_m_clock = m_clock;
   assign  _sub_plot_x_128_hikareru = data_in305;
   assign  _sub_plot_x_128_moto = data_in_index305;
   assign  _sub_plot_x_128_in_do = subs_exe;
   assign  _sub_plot_x_128_p_reset = p_reset;
   assign  _sub_plot_x_128_m_clock = m_clock;
   assign  _sub_plot_x_127_hikareru = data_in303;
   assign  _sub_plot_x_127_moto = data_in_index303;
   assign  _sub_plot_x_127_in_do = subs_exe;
   assign  _sub_plot_x_127_p_reset = p_reset;
   assign  _sub_plot_x_127_m_clock = m_clock;
   assign  _sub_plot_x_126_hikareru = data_in301;
   assign  _sub_plot_x_126_moto = data_in_index301;
   assign  _sub_plot_x_126_in_do = subs_exe;
   assign  _sub_plot_x_126_p_reset = p_reset;
   assign  _sub_plot_x_126_m_clock = m_clock;
   assign  _sub_plot_x_125_hikareru = data_in299;
   assign  _sub_plot_x_125_moto = data_in_index299;
   assign  _sub_plot_x_125_in_do = subs_exe;
   assign  _sub_plot_x_125_p_reset = p_reset;
   assign  _sub_plot_x_125_m_clock = m_clock;
   assign  _sub_plot_x_124_hikareru = data_in297;
   assign  _sub_plot_x_124_moto = data_in_index297;
   assign  _sub_plot_x_124_in_do = subs_exe;
   assign  _sub_plot_x_124_p_reset = p_reset;
   assign  _sub_plot_x_124_m_clock = m_clock;
   assign  _sub_plot_x_123_hikareru = data_in295;
   assign  _sub_plot_x_123_moto = data_in_index295;
   assign  _sub_plot_x_123_in_do = subs_exe;
   assign  _sub_plot_x_123_p_reset = p_reset;
   assign  _sub_plot_x_123_m_clock = m_clock;
   assign  _sub_plot_x_122_hikareru = data_in293;
   assign  _sub_plot_x_122_moto = data_in_index293;
   assign  _sub_plot_x_122_in_do = subs_exe;
   assign  _sub_plot_x_122_p_reset = p_reset;
   assign  _sub_plot_x_122_m_clock = m_clock;
   assign  _sub_plot_x_121_hikareru = data_in291;
   assign  _sub_plot_x_121_moto = data_in_index291;
   assign  _sub_plot_x_121_in_do = subs_exe;
   assign  _sub_plot_x_121_p_reset = p_reset;
   assign  _sub_plot_x_121_m_clock = m_clock;
   assign  _sub_plot_x_120_hikareru = data_in289;
   assign  _sub_plot_x_120_moto = data_in_index289;
   assign  _sub_plot_x_120_in_do = subs_exe;
   assign  _sub_plot_x_120_p_reset = p_reset;
   assign  _sub_plot_x_120_m_clock = m_clock;
   assign  _sub_plot_x_119_hikareru = data_in285;
   assign  _sub_plot_x_119_moto = data_in_index285;
   assign  _sub_plot_x_119_in_do = subs_exe;
   assign  _sub_plot_x_119_p_reset = p_reset;
   assign  _sub_plot_x_119_m_clock = m_clock;
   assign  _sub_plot_x_118_hikareru = data_in283;
   assign  _sub_plot_x_118_moto = data_in_index283;
   assign  _sub_plot_x_118_in_do = subs_exe;
   assign  _sub_plot_x_118_p_reset = p_reset;
   assign  _sub_plot_x_118_m_clock = m_clock;
   assign  _sub_plot_x_117_hikareru = data_in281;
   assign  _sub_plot_x_117_moto = data_in_index281;
   assign  _sub_plot_x_117_in_do = subs_exe;
   assign  _sub_plot_x_117_p_reset = p_reset;
   assign  _sub_plot_x_117_m_clock = m_clock;
   assign  _sub_plot_x_116_hikareru = data_in279;
   assign  _sub_plot_x_116_moto = data_in_index279;
   assign  _sub_plot_x_116_in_do = subs_exe;
   assign  _sub_plot_x_116_p_reset = p_reset;
   assign  _sub_plot_x_116_m_clock = m_clock;
   assign  _sub_plot_x_115_hikareru = data_in277;
   assign  _sub_plot_x_115_moto = data_in_index277;
   assign  _sub_plot_x_115_in_do = subs_exe;
   assign  _sub_plot_x_115_p_reset = p_reset;
   assign  _sub_plot_x_115_m_clock = m_clock;
   assign  _sub_plot_x_114_hikareru = data_in275;
   assign  _sub_plot_x_114_moto = data_in_index275;
   assign  _sub_plot_x_114_in_do = subs_exe;
   assign  _sub_plot_x_114_p_reset = p_reset;
   assign  _sub_plot_x_114_m_clock = m_clock;
   assign  _sub_plot_x_113_hikareru = data_in273;
   assign  _sub_plot_x_113_moto = data_in_index273;
   assign  _sub_plot_x_113_in_do = subs_exe;
   assign  _sub_plot_x_113_p_reset = p_reset;
   assign  _sub_plot_x_113_m_clock = m_clock;
   assign  _sub_plot_x_112_hikareru = data_in271;
   assign  _sub_plot_x_112_moto = data_in_index271;
   assign  _sub_plot_x_112_in_do = subs_exe;
   assign  _sub_plot_x_112_p_reset = p_reset;
   assign  _sub_plot_x_112_m_clock = m_clock;
   assign  _sub_plot_x_111_hikareru = data_in269;
   assign  _sub_plot_x_111_moto = data_in_index269;
   assign  _sub_plot_x_111_in_do = subs_exe;
   assign  _sub_plot_x_111_p_reset = p_reset;
   assign  _sub_plot_x_111_m_clock = m_clock;
   assign  _sub_plot_x_110_hikareru = data_in267;
   assign  _sub_plot_x_110_moto = data_in_index267;
   assign  _sub_plot_x_110_in_do = subs_exe;
   assign  _sub_plot_x_110_p_reset = p_reset;
   assign  _sub_plot_x_110_m_clock = m_clock;
   assign  _sub_plot_x_109_hikareru = data_in265;
   assign  _sub_plot_x_109_moto = data_in_index265;
   assign  _sub_plot_x_109_in_do = subs_exe;
   assign  _sub_plot_x_109_p_reset = p_reset;
   assign  _sub_plot_x_109_m_clock = m_clock;
   assign  _sub_plot_x_108_hikareru = data_in263;
   assign  _sub_plot_x_108_moto = data_in_index263;
   assign  _sub_plot_x_108_in_do = subs_exe;
   assign  _sub_plot_x_108_p_reset = p_reset;
   assign  _sub_plot_x_108_m_clock = m_clock;
   assign  _sub_plot_x_107_hikareru = data_in261;
   assign  _sub_plot_x_107_moto = data_in_index261;
   assign  _sub_plot_x_107_in_do = subs_exe;
   assign  _sub_plot_x_107_p_reset = p_reset;
   assign  _sub_plot_x_107_m_clock = m_clock;
   assign  _sub_plot_x_106_hikareru = data_in259;
   assign  _sub_plot_x_106_moto = data_in_index259;
   assign  _sub_plot_x_106_in_do = subs_exe;
   assign  _sub_plot_x_106_p_reset = p_reset;
   assign  _sub_plot_x_106_m_clock = m_clock;
   assign  _sub_plot_x_105_hikareru = data_in257;
   assign  _sub_plot_x_105_moto = data_in_index257;
   assign  _sub_plot_x_105_in_do = subs_exe;
   assign  _sub_plot_x_105_p_reset = p_reset;
   assign  _sub_plot_x_105_m_clock = m_clock;
   assign  _sub_plot_x_104_hikareru = data_in253;
   assign  _sub_plot_x_104_moto = data_in_index253;
   assign  _sub_plot_x_104_in_do = subs_exe;
   assign  _sub_plot_x_104_p_reset = p_reset;
   assign  _sub_plot_x_104_m_clock = m_clock;
   assign  _sub_plot_x_103_hikareru = data_in251;
   assign  _sub_plot_x_103_moto = data_in_index251;
   assign  _sub_plot_x_103_in_do = subs_exe;
   assign  _sub_plot_x_103_p_reset = p_reset;
   assign  _sub_plot_x_103_m_clock = m_clock;
   assign  _sub_plot_x_102_hikareru = data_in249;
   assign  _sub_plot_x_102_moto = data_in_index249;
   assign  _sub_plot_x_102_in_do = subs_exe;
   assign  _sub_plot_x_102_p_reset = p_reset;
   assign  _sub_plot_x_102_m_clock = m_clock;
   assign  _sub_plot_x_101_hikareru = data_in247;
   assign  _sub_plot_x_101_moto = data_in_index247;
   assign  _sub_plot_x_101_in_do = subs_exe;
   assign  _sub_plot_x_101_p_reset = p_reset;
   assign  _sub_plot_x_101_m_clock = m_clock;
   assign  _sub_plot_x_100_hikareru = data_in245;
   assign  _sub_plot_x_100_moto = data_in_index245;
   assign  _sub_plot_x_100_in_do = subs_exe;
   assign  _sub_plot_x_100_p_reset = p_reset;
   assign  _sub_plot_x_100_m_clock = m_clock;
   assign  _sub_plot_x_99_hikareru = data_in243;
   assign  _sub_plot_x_99_moto = data_in_index243;
   assign  _sub_plot_x_99_in_do = subs_exe;
   assign  _sub_plot_x_99_p_reset = p_reset;
   assign  _sub_plot_x_99_m_clock = m_clock;
   assign  _sub_plot_x_98_hikareru = data_in241;
   assign  _sub_plot_x_98_moto = data_in_index241;
   assign  _sub_plot_x_98_in_do = subs_exe;
   assign  _sub_plot_x_98_p_reset = p_reset;
   assign  _sub_plot_x_98_m_clock = m_clock;
   assign  _sub_plot_x_97_hikareru = data_in239;
   assign  _sub_plot_x_97_moto = data_in_index239;
   assign  _sub_plot_x_97_in_do = subs_exe;
   assign  _sub_plot_x_97_p_reset = p_reset;
   assign  _sub_plot_x_97_m_clock = m_clock;
   assign  _sub_plot_x_96_hikareru = data_in237;
   assign  _sub_plot_x_96_moto = data_in_index237;
   assign  _sub_plot_x_96_in_do = subs_exe;
   assign  _sub_plot_x_96_p_reset = p_reset;
   assign  _sub_plot_x_96_m_clock = m_clock;
   assign  _sub_plot_x_95_hikareru = data_in235;
   assign  _sub_plot_x_95_moto = data_in_index235;
   assign  _sub_plot_x_95_in_do = subs_exe;
   assign  _sub_plot_x_95_p_reset = p_reset;
   assign  _sub_plot_x_95_m_clock = m_clock;
   assign  _sub_plot_x_94_hikareru = data_in233;
   assign  _sub_plot_x_94_moto = data_in_index233;
   assign  _sub_plot_x_94_in_do = subs_exe;
   assign  _sub_plot_x_94_p_reset = p_reset;
   assign  _sub_plot_x_94_m_clock = m_clock;
   assign  _sub_plot_x_93_hikareru = data_in231;
   assign  _sub_plot_x_93_moto = data_in_index231;
   assign  _sub_plot_x_93_in_do = subs_exe;
   assign  _sub_plot_x_93_p_reset = p_reset;
   assign  _sub_plot_x_93_m_clock = m_clock;
   assign  _sub_plot_x_92_hikareru = data_in229;
   assign  _sub_plot_x_92_moto = data_in_index229;
   assign  _sub_plot_x_92_in_do = subs_exe;
   assign  _sub_plot_x_92_p_reset = p_reset;
   assign  _sub_plot_x_92_m_clock = m_clock;
   assign  _sub_plot_x_91_hikareru = data_in227;
   assign  _sub_plot_x_91_moto = data_in_index227;
   assign  _sub_plot_x_91_in_do = subs_exe;
   assign  _sub_plot_x_91_p_reset = p_reset;
   assign  _sub_plot_x_91_m_clock = m_clock;
   assign  _sub_plot_x_90_hikareru = data_in225;
   assign  _sub_plot_x_90_moto = data_in_index225;
   assign  _sub_plot_x_90_in_do = subs_exe;
   assign  _sub_plot_x_90_p_reset = p_reset;
   assign  _sub_plot_x_90_m_clock = m_clock;
   assign  _sub_plot_x_89_hikareru = data_in221;
   assign  _sub_plot_x_89_moto = data_in_index221;
   assign  _sub_plot_x_89_in_do = subs_exe;
   assign  _sub_plot_x_89_p_reset = p_reset;
   assign  _sub_plot_x_89_m_clock = m_clock;
   assign  _sub_plot_x_88_hikareru = data_in219;
   assign  _sub_plot_x_88_moto = data_in_index219;
   assign  _sub_plot_x_88_in_do = subs_exe;
   assign  _sub_plot_x_88_p_reset = p_reset;
   assign  _sub_plot_x_88_m_clock = m_clock;
   assign  _sub_plot_x_87_hikareru = data_in217;
   assign  _sub_plot_x_87_moto = data_in_index217;
   assign  _sub_plot_x_87_in_do = subs_exe;
   assign  _sub_plot_x_87_p_reset = p_reset;
   assign  _sub_plot_x_87_m_clock = m_clock;
   assign  _sub_plot_x_86_hikareru = data_in215;
   assign  _sub_plot_x_86_moto = data_in_index215;
   assign  _sub_plot_x_86_in_do = subs_exe;
   assign  _sub_plot_x_86_p_reset = p_reset;
   assign  _sub_plot_x_86_m_clock = m_clock;
   assign  _sub_plot_x_85_hikareru = data_in213;
   assign  _sub_plot_x_85_moto = data_in_index213;
   assign  _sub_plot_x_85_in_do = subs_exe;
   assign  _sub_plot_x_85_p_reset = p_reset;
   assign  _sub_plot_x_85_m_clock = m_clock;
   assign  _sub_plot_x_84_hikareru = data_in211;
   assign  _sub_plot_x_84_moto = data_in_index211;
   assign  _sub_plot_x_84_in_do = subs_exe;
   assign  _sub_plot_x_84_p_reset = p_reset;
   assign  _sub_plot_x_84_m_clock = m_clock;
   assign  _sub_plot_x_83_hikareru = data_in209;
   assign  _sub_plot_x_83_moto = data_in_index209;
   assign  _sub_plot_x_83_in_do = subs_exe;
   assign  _sub_plot_x_83_p_reset = p_reset;
   assign  _sub_plot_x_83_m_clock = m_clock;
   assign  _sub_plot_x_82_hikareru = data_in207;
   assign  _sub_plot_x_82_moto = data_in_index207;
   assign  _sub_plot_x_82_in_do = subs_exe;
   assign  _sub_plot_x_82_p_reset = p_reset;
   assign  _sub_plot_x_82_m_clock = m_clock;
   assign  _sub_plot_x_81_hikareru = data_in205;
   assign  _sub_plot_x_81_moto = data_in_index205;
   assign  _sub_plot_x_81_in_do = subs_exe;
   assign  _sub_plot_x_81_p_reset = p_reset;
   assign  _sub_plot_x_81_m_clock = m_clock;
   assign  _sub_plot_x_80_hikareru = data_in203;
   assign  _sub_plot_x_80_moto = data_in_index203;
   assign  _sub_plot_x_80_in_do = subs_exe;
   assign  _sub_plot_x_80_p_reset = p_reset;
   assign  _sub_plot_x_80_m_clock = m_clock;
   assign  _sub_plot_x_79_hikareru = data_in201;
   assign  _sub_plot_x_79_moto = data_in_index201;
   assign  _sub_plot_x_79_in_do = subs_exe;
   assign  _sub_plot_x_79_p_reset = p_reset;
   assign  _sub_plot_x_79_m_clock = m_clock;
   assign  _sub_plot_x_78_hikareru = data_in199;
   assign  _sub_plot_x_78_moto = data_in_index199;
   assign  _sub_plot_x_78_in_do = subs_exe;
   assign  _sub_plot_x_78_p_reset = p_reset;
   assign  _sub_plot_x_78_m_clock = m_clock;
   assign  _sub_plot_x_77_hikareru = data_in197;
   assign  _sub_plot_x_77_moto = data_in_index197;
   assign  _sub_plot_x_77_in_do = subs_exe;
   assign  _sub_plot_x_77_p_reset = p_reset;
   assign  _sub_plot_x_77_m_clock = m_clock;
   assign  _sub_plot_x_76_hikareru = data_in195;
   assign  _sub_plot_x_76_moto = data_in_index195;
   assign  _sub_plot_x_76_in_do = subs_exe;
   assign  _sub_plot_x_76_p_reset = p_reset;
   assign  _sub_plot_x_76_m_clock = m_clock;
   assign  _sub_plot_x_75_hikareru = data_in193;
   assign  _sub_plot_x_75_moto = data_in_index193;
   assign  _sub_plot_x_75_in_do = subs_exe;
   assign  _sub_plot_x_75_p_reset = p_reset;
   assign  _sub_plot_x_75_m_clock = m_clock;
   assign  _sub_plot_x_74_hikareru = data_in189;
   assign  _sub_plot_x_74_moto = data_in_index189;
   assign  _sub_plot_x_74_in_do = subs_exe;
   assign  _sub_plot_x_74_p_reset = p_reset;
   assign  _sub_plot_x_74_m_clock = m_clock;
   assign  _sub_plot_x_73_hikareru = data_in187;
   assign  _sub_plot_x_73_moto = data_in_index187;
   assign  _sub_plot_x_73_in_do = subs_exe;
   assign  _sub_plot_x_73_p_reset = p_reset;
   assign  _sub_plot_x_73_m_clock = m_clock;
   assign  _sub_plot_x_72_hikareru = data_in185;
   assign  _sub_plot_x_72_moto = data_in_index185;
   assign  _sub_plot_x_72_in_do = subs_exe;
   assign  _sub_plot_x_72_p_reset = p_reset;
   assign  _sub_plot_x_72_m_clock = m_clock;
   assign  _sub_plot_x_71_hikareru = data_in183;
   assign  _sub_plot_x_71_moto = data_in_index183;
   assign  _sub_plot_x_71_in_do = subs_exe;
   assign  _sub_plot_x_71_p_reset = p_reset;
   assign  _sub_plot_x_71_m_clock = m_clock;
   assign  _sub_plot_x_70_hikareru = data_in181;
   assign  _sub_plot_x_70_moto = data_in_index181;
   assign  _sub_plot_x_70_in_do = subs_exe;
   assign  _sub_plot_x_70_p_reset = p_reset;
   assign  _sub_plot_x_70_m_clock = m_clock;
   assign  _sub_plot_x_69_hikareru = data_in179;
   assign  _sub_plot_x_69_moto = data_in_index179;
   assign  _sub_plot_x_69_in_do = subs_exe;
   assign  _sub_plot_x_69_p_reset = p_reset;
   assign  _sub_plot_x_69_m_clock = m_clock;
   assign  _sub_plot_x_68_hikareru = data_in177;
   assign  _sub_plot_x_68_moto = data_in_index177;
   assign  _sub_plot_x_68_in_do = subs_exe;
   assign  _sub_plot_x_68_p_reset = p_reset;
   assign  _sub_plot_x_68_m_clock = m_clock;
   assign  _sub_plot_x_67_hikareru = data_in175;
   assign  _sub_plot_x_67_moto = data_in_index175;
   assign  _sub_plot_x_67_in_do = subs_exe;
   assign  _sub_plot_x_67_p_reset = p_reset;
   assign  _sub_plot_x_67_m_clock = m_clock;
   assign  _sub_plot_x_66_hikareru = data_in173;
   assign  _sub_plot_x_66_moto = data_in_index173;
   assign  _sub_plot_x_66_in_do = subs_exe;
   assign  _sub_plot_x_66_p_reset = p_reset;
   assign  _sub_plot_x_66_m_clock = m_clock;
   assign  _sub_plot_x_65_hikareru = data_in171;
   assign  _sub_plot_x_65_moto = data_in_index171;
   assign  _sub_plot_x_65_in_do = subs_exe;
   assign  _sub_plot_x_65_p_reset = p_reset;
   assign  _sub_plot_x_65_m_clock = m_clock;
   assign  _sub_plot_x_64_hikareru = data_in169;
   assign  _sub_plot_x_64_moto = data_in_index169;
   assign  _sub_plot_x_64_in_do = subs_exe;
   assign  _sub_plot_x_64_p_reset = p_reset;
   assign  _sub_plot_x_64_m_clock = m_clock;
   assign  _sub_plot_x_63_hikareru = data_in167;
   assign  _sub_plot_x_63_moto = data_in_index167;
   assign  _sub_plot_x_63_in_do = subs_exe;
   assign  _sub_plot_x_63_p_reset = p_reset;
   assign  _sub_plot_x_63_m_clock = m_clock;
   assign  _sub_plot_x_62_hikareru = data_in165;
   assign  _sub_plot_x_62_moto = data_in_index165;
   assign  _sub_plot_x_62_in_do = subs_exe;
   assign  _sub_plot_x_62_p_reset = p_reset;
   assign  _sub_plot_x_62_m_clock = m_clock;
   assign  _sub_plot_x_61_hikareru = data_in163;
   assign  _sub_plot_x_61_moto = data_in_index163;
   assign  _sub_plot_x_61_in_do = subs_exe;
   assign  _sub_plot_x_61_p_reset = p_reset;
   assign  _sub_plot_x_61_m_clock = m_clock;
   assign  _sub_plot_x_60_hikareru = data_in161;
   assign  _sub_plot_x_60_moto = data_in_index161;
   assign  _sub_plot_x_60_in_do = subs_exe;
   assign  _sub_plot_x_60_p_reset = p_reset;
   assign  _sub_plot_x_60_m_clock = m_clock;
   assign  _sub_plot_x_59_hikareru = data_in157;
   assign  _sub_plot_x_59_moto = data_in_index157;
   assign  _sub_plot_x_59_in_do = subs_exe;
   assign  _sub_plot_x_59_p_reset = p_reset;
   assign  _sub_plot_x_59_m_clock = m_clock;
   assign  _sub_plot_x_58_hikareru = data_in155;
   assign  _sub_plot_x_58_moto = data_in_index155;
   assign  _sub_plot_x_58_in_do = subs_exe;
   assign  _sub_plot_x_58_p_reset = p_reset;
   assign  _sub_plot_x_58_m_clock = m_clock;
   assign  _sub_plot_x_57_hikareru = data_in153;
   assign  _sub_plot_x_57_moto = data_in_index153;
   assign  _sub_plot_x_57_in_do = subs_exe;
   assign  _sub_plot_x_57_p_reset = p_reset;
   assign  _sub_plot_x_57_m_clock = m_clock;
   assign  _sub_plot_x_56_hikareru = data_in151;
   assign  _sub_plot_x_56_moto = data_in_index151;
   assign  _sub_plot_x_56_in_do = subs_exe;
   assign  _sub_plot_x_56_p_reset = p_reset;
   assign  _sub_plot_x_56_m_clock = m_clock;
   assign  _sub_plot_x_55_hikareru = data_in149;
   assign  _sub_plot_x_55_moto = data_in_index149;
   assign  _sub_plot_x_55_in_do = subs_exe;
   assign  _sub_plot_x_55_p_reset = p_reset;
   assign  _sub_plot_x_55_m_clock = m_clock;
   assign  _sub_plot_x_54_hikareru = data_in147;
   assign  _sub_plot_x_54_moto = data_in_index147;
   assign  _sub_plot_x_54_in_do = subs_exe;
   assign  _sub_plot_x_54_p_reset = p_reset;
   assign  _sub_plot_x_54_m_clock = m_clock;
   assign  _sub_plot_x_53_hikareru = data_in145;
   assign  _sub_plot_x_53_moto = data_in_index145;
   assign  _sub_plot_x_53_in_do = subs_exe;
   assign  _sub_plot_x_53_p_reset = p_reset;
   assign  _sub_plot_x_53_m_clock = m_clock;
   assign  _sub_plot_x_52_hikareru = data_in143;
   assign  _sub_plot_x_52_moto = data_in_index143;
   assign  _sub_plot_x_52_in_do = subs_exe;
   assign  _sub_plot_x_52_p_reset = p_reset;
   assign  _sub_plot_x_52_m_clock = m_clock;
   assign  _sub_plot_x_51_hikareru = data_in141;
   assign  _sub_plot_x_51_moto = data_in_index141;
   assign  _sub_plot_x_51_in_do = subs_exe;
   assign  _sub_plot_x_51_p_reset = p_reset;
   assign  _sub_plot_x_51_m_clock = m_clock;
   assign  _sub_plot_x_50_hikareru = data_in139;
   assign  _sub_plot_x_50_moto = data_in_index139;
   assign  _sub_plot_x_50_in_do = subs_exe;
   assign  _sub_plot_x_50_p_reset = p_reset;
   assign  _sub_plot_x_50_m_clock = m_clock;
   assign  _sub_plot_x_49_hikareru = data_in137;
   assign  _sub_plot_x_49_moto = data_in_index137;
   assign  _sub_plot_x_49_in_do = subs_exe;
   assign  _sub_plot_x_49_p_reset = p_reset;
   assign  _sub_plot_x_49_m_clock = m_clock;
   assign  _sub_plot_x_48_hikareru = data_in135;
   assign  _sub_plot_x_48_moto = data_in_index135;
   assign  _sub_plot_x_48_in_do = subs_exe;
   assign  _sub_plot_x_48_p_reset = p_reset;
   assign  _sub_plot_x_48_m_clock = m_clock;
   assign  _sub_plot_x_47_hikareru = data_in133;
   assign  _sub_plot_x_47_moto = data_in_index133;
   assign  _sub_plot_x_47_in_do = subs_exe;
   assign  _sub_plot_x_47_p_reset = p_reset;
   assign  _sub_plot_x_47_m_clock = m_clock;
   assign  _sub_plot_x_46_hikareru = data_in131;
   assign  _sub_plot_x_46_moto = data_in_index131;
   assign  _sub_plot_x_46_in_do = subs_exe;
   assign  _sub_plot_x_46_p_reset = p_reset;
   assign  _sub_plot_x_46_m_clock = m_clock;
   assign  _sub_plot_x_45_hikareru = data_in129;
   assign  _sub_plot_x_45_moto = data_in_index129;
   assign  _sub_plot_x_45_in_do = subs_exe;
   assign  _sub_plot_x_45_p_reset = p_reset;
   assign  _sub_plot_x_45_m_clock = m_clock;
   assign  _sub_plot_x_44_hikareru = data_in125;
   assign  _sub_plot_x_44_moto = data_in_index125;
   assign  _sub_plot_x_44_in_do = subs_exe;
   assign  _sub_plot_x_44_p_reset = p_reset;
   assign  _sub_plot_x_44_m_clock = m_clock;
   assign  _sub_plot_x_43_hikareru = data_in123;
   assign  _sub_plot_x_43_moto = data_in_index123;
   assign  _sub_plot_x_43_in_do = subs_exe;
   assign  _sub_plot_x_43_p_reset = p_reset;
   assign  _sub_plot_x_43_m_clock = m_clock;
   assign  _sub_plot_x_42_hikareru = data_in121;
   assign  _sub_plot_x_42_moto = data_in_index121;
   assign  _sub_plot_x_42_in_do = subs_exe;
   assign  _sub_plot_x_42_p_reset = p_reset;
   assign  _sub_plot_x_42_m_clock = m_clock;
   assign  _sub_plot_x_41_hikareru = data_in119;
   assign  _sub_plot_x_41_moto = data_in_index119;
   assign  _sub_plot_x_41_in_do = subs_exe;
   assign  _sub_plot_x_41_p_reset = p_reset;
   assign  _sub_plot_x_41_m_clock = m_clock;
   assign  _sub_plot_x_40_hikareru = data_in117;
   assign  _sub_plot_x_40_moto = data_in_index117;
   assign  _sub_plot_x_40_in_do = subs_exe;
   assign  _sub_plot_x_40_p_reset = p_reset;
   assign  _sub_plot_x_40_m_clock = m_clock;
   assign  _sub_plot_x_39_hikareru = data_in115;
   assign  _sub_plot_x_39_moto = data_in_index115;
   assign  _sub_plot_x_39_in_do = subs_exe;
   assign  _sub_plot_x_39_p_reset = p_reset;
   assign  _sub_plot_x_39_m_clock = m_clock;
   assign  _sub_plot_x_38_hikareru = data_in113;
   assign  _sub_plot_x_38_moto = data_in_index113;
   assign  _sub_plot_x_38_in_do = subs_exe;
   assign  _sub_plot_x_38_p_reset = p_reset;
   assign  _sub_plot_x_38_m_clock = m_clock;
   assign  _sub_plot_x_37_hikareru = data_in111;
   assign  _sub_plot_x_37_moto = data_in_index111;
   assign  _sub_plot_x_37_in_do = subs_exe;
   assign  _sub_plot_x_37_p_reset = p_reset;
   assign  _sub_plot_x_37_m_clock = m_clock;
   assign  _sub_plot_x_36_hikareru = data_in109;
   assign  _sub_plot_x_36_moto = data_in_index109;
   assign  _sub_plot_x_36_in_do = subs_exe;
   assign  _sub_plot_x_36_p_reset = p_reset;
   assign  _sub_plot_x_36_m_clock = m_clock;
   assign  _sub_plot_x_35_hikareru = data_in107;
   assign  _sub_plot_x_35_moto = data_in_index107;
   assign  _sub_plot_x_35_in_do = subs_exe;
   assign  _sub_plot_x_35_p_reset = p_reset;
   assign  _sub_plot_x_35_m_clock = m_clock;
   assign  _sub_plot_x_34_hikareru = data_in105;
   assign  _sub_plot_x_34_moto = data_in_index105;
   assign  _sub_plot_x_34_in_do = subs_exe;
   assign  _sub_plot_x_34_p_reset = p_reset;
   assign  _sub_plot_x_34_m_clock = m_clock;
   assign  _sub_plot_x_33_hikareru = data_in103;
   assign  _sub_plot_x_33_moto = data_in_index103;
   assign  _sub_plot_x_33_in_do = subs_exe;
   assign  _sub_plot_x_33_p_reset = p_reset;
   assign  _sub_plot_x_33_m_clock = m_clock;
   assign  _sub_plot_x_32_hikareru = data_in101;
   assign  _sub_plot_x_32_moto = data_in_index101;
   assign  _sub_plot_x_32_in_do = subs_exe;
   assign  _sub_plot_x_32_p_reset = p_reset;
   assign  _sub_plot_x_32_m_clock = m_clock;
   assign  _sub_plot_x_31_hikareru = data_in99;
   assign  _sub_plot_x_31_moto = data_in_index99;
   assign  _sub_plot_x_31_in_do = subs_exe;
   assign  _sub_plot_x_31_p_reset = p_reset;
   assign  _sub_plot_x_31_m_clock = m_clock;
   assign  _sub_plot_x_30_hikareru = data_in97;
   assign  _sub_plot_x_30_moto = data_in_index97;
   assign  _sub_plot_x_30_in_do = subs_exe;
   assign  _sub_plot_x_30_p_reset = p_reset;
   assign  _sub_plot_x_30_m_clock = m_clock;
   assign  _sub_plot_x_29_hikareru = data_in93;
   assign  _sub_plot_x_29_moto = data_in_index93;
   assign  _sub_plot_x_29_in_do = subs_exe;
   assign  _sub_plot_x_29_p_reset = p_reset;
   assign  _sub_plot_x_29_m_clock = m_clock;
   assign  _sub_plot_x_28_hikareru = data_in91;
   assign  _sub_plot_x_28_moto = data_in_index91;
   assign  _sub_plot_x_28_in_do = subs_exe;
   assign  _sub_plot_x_28_p_reset = p_reset;
   assign  _sub_plot_x_28_m_clock = m_clock;
   assign  _sub_plot_x_27_hikareru = data_in89;
   assign  _sub_plot_x_27_moto = data_in_index89;
   assign  _sub_plot_x_27_in_do = subs_exe;
   assign  _sub_plot_x_27_p_reset = p_reset;
   assign  _sub_plot_x_27_m_clock = m_clock;
   assign  _sub_plot_x_26_hikareru = data_in87;
   assign  _sub_plot_x_26_moto = data_in_index87;
   assign  _sub_plot_x_26_in_do = subs_exe;
   assign  _sub_plot_x_26_p_reset = p_reset;
   assign  _sub_plot_x_26_m_clock = m_clock;
   assign  _sub_plot_x_25_hikareru = data_in85;
   assign  _sub_plot_x_25_moto = data_in_index85;
   assign  _sub_plot_x_25_in_do = subs_exe;
   assign  _sub_plot_x_25_p_reset = p_reset;
   assign  _sub_plot_x_25_m_clock = m_clock;
   assign  _sub_plot_x_24_hikareru = data_in83;
   assign  _sub_plot_x_24_moto = data_in_index83;
   assign  _sub_plot_x_24_in_do = subs_exe;
   assign  _sub_plot_x_24_p_reset = p_reset;
   assign  _sub_plot_x_24_m_clock = m_clock;
   assign  _sub_plot_x_23_hikareru = data_in81;
   assign  _sub_plot_x_23_moto = data_in_index81;
   assign  _sub_plot_x_23_in_do = subs_exe;
   assign  _sub_plot_x_23_p_reset = p_reset;
   assign  _sub_plot_x_23_m_clock = m_clock;
   assign  _sub_plot_x_22_hikareru = data_in79;
   assign  _sub_plot_x_22_moto = data_in_index79;
   assign  _sub_plot_x_22_in_do = subs_exe;
   assign  _sub_plot_x_22_p_reset = p_reset;
   assign  _sub_plot_x_22_m_clock = m_clock;
   assign  _sub_plot_x_21_hikareru = data_in77;
   assign  _sub_plot_x_21_moto = data_in_index77;
   assign  _sub_plot_x_21_in_do = subs_exe;
   assign  _sub_plot_x_21_p_reset = p_reset;
   assign  _sub_plot_x_21_m_clock = m_clock;
   assign  _sub_plot_x_20_hikareru = data_in75;
   assign  _sub_plot_x_20_moto = data_in_index75;
   assign  _sub_plot_x_20_in_do = subs_exe;
   assign  _sub_plot_x_20_p_reset = p_reset;
   assign  _sub_plot_x_20_m_clock = m_clock;
   assign  _sub_plot_x_19_hikareru = data_in73;
   assign  _sub_plot_x_19_moto = data_in_index73;
   assign  _sub_plot_x_19_in_do = subs_exe;
   assign  _sub_plot_x_19_p_reset = p_reset;
   assign  _sub_plot_x_19_m_clock = m_clock;
   assign  _sub_plot_x_18_hikareru = data_in71;
   assign  _sub_plot_x_18_moto = data_in_index71;
   assign  _sub_plot_x_18_in_do = subs_exe;
   assign  _sub_plot_x_18_p_reset = p_reset;
   assign  _sub_plot_x_18_m_clock = m_clock;
   assign  _sub_plot_x_17_hikareru = data_in69;
   assign  _sub_plot_x_17_moto = data_in_index69;
   assign  _sub_plot_x_17_in_do = subs_exe;
   assign  _sub_plot_x_17_p_reset = p_reset;
   assign  _sub_plot_x_17_m_clock = m_clock;
   assign  _sub_plot_x_16_hikareru = data_in67;
   assign  _sub_plot_x_16_moto = data_in_index67;
   assign  _sub_plot_x_16_in_do = subs_exe;
   assign  _sub_plot_x_16_p_reset = p_reset;
   assign  _sub_plot_x_16_m_clock = m_clock;
   assign  _sub_plot_x_15_hikareru = data_in65;
   assign  _sub_plot_x_15_moto = data_in_index65;
   assign  _sub_plot_x_15_in_do = subs_exe;
   assign  _sub_plot_x_15_p_reset = p_reset;
   assign  _sub_plot_x_15_m_clock = m_clock;
   assign  _sub_plot_x_14_hikareru = data_in61;
   assign  _sub_plot_x_14_moto = data_in_index61;
   assign  _sub_plot_x_14_in_do = subs_exe;
   assign  _sub_plot_x_14_p_reset = p_reset;
   assign  _sub_plot_x_14_m_clock = m_clock;
   assign  _sub_plot_x_13_hikareru = data_in59;
   assign  _sub_plot_x_13_moto = data_in_index59;
   assign  _sub_plot_x_13_in_do = subs_exe;
   assign  _sub_plot_x_13_p_reset = p_reset;
   assign  _sub_plot_x_13_m_clock = m_clock;
   assign  _sub_plot_x_12_hikareru = data_in57;
   assign  _sub_plot_x_12_moto = data_in_index57;
   assign  _sub_plot_x_12_in_do = subs_exe;
   assign  _sub_plot_x_12_p_reset = p_reset;
   assign  _sub_plot_x_12_m_clock = m_clock;
   assign  _sub_plot_x_11_hikareru = data_in55;
   assign  _sub_plot_x_11_moto = data_in_index55;
   assign  _sub_plot_x_11_in_do = subs_exe;
   assign  _sub_plot_x_11_p_reset = p_reset;
   assign  _sub_plot_x_11_m_clock = m_clock;
   assign  _sub_plot_x_10_hikareru = data_in53;
   assign  _sub_plot_x_10_moto = data_in_index53;
   assign  _sub_plot_x_10_in_do = subs_exe;
   assign  _sub_plot_x_10_p_reset = p_reset;
   assign  _sub_plot_x_10_m_clock = m_clock;
   assign  _sub_plot_x_9_hikareru = data_in51;
   assign  _sub_plot_x_9_moto = data_in_index51;
   assign  _sub_plot_x_9_in_do = subs_exe;
   assign  _sub_plot_x_9_p_reset = p_reset;
   assign  _sub_plot_x_9_m_clock = m_clock;
   assign  _sub_plot_x_8_hikareru = data_in49;
   assign  _sub_plot_x_8_moto = data_in_index49;
   assign  _sub_plot_x_8_in_do = subs_exe;
   assign  _sub_plot_x_8_p_reset = p_reset;
   assign  _sub_plot_x_8_m_clock = m_clock;
   assign  _sub_plot_x_7_hikareru = data_in47;
   assign  _sub_plot_x_7_moto = data_in_index47;
   assign  _sub_plot_x_7_in_do = subs_exe;
   assign  _sub_plot_x_7_p_reset = p_reset;
   assign  _sub_plot_x_7_m_clock = m_clock;
   assign  _sub_plot_x_6_hikareru = data_in45;
   assign  _sub_plot_x_6_moto = data_in_index45;
   assign  _sub_plot_x_6_in_do = subs_exe;
   assign  _sub_plot_x_6_p_reset = p_reset;
   assign  _sub_plot_x_6_m_clock = m_clock;
   assign  _sub_plot_x_5_hikareru = data_in43;
   assign  _sub_plot_x_5_moto = data_in_index43;
   assign  _sub_plot_x_5_in_do = subs_exe;
   assign  _sub_plot_x_5_p_reset = p_reset;
   assign  _sub_plot_x_5_m_clock = m_clock;
   assign  _sub_plot_x_4_hikareru = data_in41;
   assign  _sub_plot_x_4_moto = data_in_index41;
   assign  _sub_plot_x_4_in_do = subs_exe;
   assign  _sub_plot_x_4_p_reset = p_reset;
   assign  _sub_plot_x_4_m_clock = m_clock;
   assign  _sub_plot_x_3_hikareru = data_in39;
   assign  _sub_plot_x_3_moto = data_in_index39;
   assign  _sub_plot_x_3_in_do = subs_exe;
   assign  _sub_plot_x_3_p_reset = p_reset;
   assign  _sub_plot_x_3_m_clock = m_clock;
   assign  _sub_plot_x_2_hikareru = data_in37;
   assign  _sub_plot_x_2_moto = data_in_index37;
   assign  _sub_plot_x_2_in_do = subs_exe;
   assign  _sub_plot_x_2_p_reset = p_reset;
   assign  _sub_plot_x_2_m_clock = m_clock;
   assign  _sub_plot_x_1_hikareru = data_in35;
   assign  _sub_plot_x_1_moto = data_in_index35;
   assign  _sub_plot_x_1_in_do = subs_exe;
   assign  _sub_plot_x_1_p_reset = p_reset;
   assign  _sub_plot_x_1_m_clock = m_clock;
   assign  sub_array_out = sub_reg;
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     sub_reg <= 10'b0000000000;
else if ((subs_exe)) 
      sub_reg <= (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_sub_plot_x_sa|_sub_plot_x_1_sa)|_sub_plot_x_2_sa)|_sub_plot_x_3_sa)|_sub_plot_x_4_sa)|_sub_plot_x_5_sa)|_sub_plot_x_6_sa)|_sub_plot_x_7_sa)|_sub_plot_x_8_sa)|_sub_plot_x_9_sa)|_sub_plot_x_10_sa)|_sub_plot_x_11_sa)|_sub_plot_x_12_sa)|_sub_plot_x_13_sa)|_sub_plot_x_14_sa)|_sub_plot_x_15_sa)|_sub_plot_x_16_sa)|_sub_plot_x_17_sa)|_sub_plot_x_18_sa)|_sub_plot_x_19_sa)|_sub_plot_x_20_sa)|_sub_plot_x_21_sa)|_sub_plot_x_22_sa)|_sub_plot_x_23_sa)|_sub_plot_x_24_sa)|_sub_plot_x_25_sa)|_sub_plot_x_26_sa)|_sub_plot_x_27_sa)|_sub_plot_x_28_sa)|_sub_plot_x_29_sa)|_sub_plot_x_30_sa)|_sub_plot_x_31_sa)|_sub_plot_x_32_sa)|_sub_plot_x_33_sa)|_sub_plot_x_34_sa)|_sub_plot_x_35_sa)|_sub_plot_x_36_sa)|_sub_plot_x_37_sa)|_sub_plot_x_38_sa)|_sub_plot_x_39_sa)|_sub_plot_x_40_sa)|_sub_plot_x_41_sa)|_sub_plot_x_42_sa)|_sub_plot_x_43_sa)|_sub_plot_x_44_sa)|_sub_plot_x_45_sa)|_sub_plot_x_46_sa)|_sub_plot_x_47_sa)|_sub_plot_x_48_sa)|_sub_plot_x_49_sa)|_sub_plot_x_50_sa)|_sub_plot_x_51_sa)|_sub_plot_x_52_sa)|_sub_plot_x_53_sa)|_sub_plot_x_54_sa)|_sub_plot_x_55_sa)|_sub_plot_x_56_sa)|_sub_plot_x_57_sa)|_sub_plot_x_58_sa)|_sub_plot_x_59_sa)|_sub_plot_x_60_sa)|_sub_plot_x_61_sa)|_sub_plot_x_62_sa)|_sub_plot_x_63_sa)|_sub_plot_x_64_sa)|_sub_plot_x_65_sa)|_sub_plot_x_66_sa)|_sub_plot_x_67_sa)|_sub_plot_x_68_sa)|_sub_plot_x_69_sa)|_sub_plot_x_70_sa)|_sub_plot_x_71_sa)|_sub_plot_x_72_sa)|_sub_plot_x_73_sa)|_sub_plot_x_74_sa)|_sub_plot_x_75_sa)|_sub_plot_x_76_sa)|_sub_plot_x_77_sa)|_sub_plot_x_78_sa)|_sub_plot_x_79_sa)|_sub_plot_x_80_sa)|_sub_plot_x_81_sa)|_sub_plot_x_82_sa)|_sub_plot_x_83_sa)|_sub_plot_x_84_sa)|_sub_plot_x_85_sa)|_sub_plot_x_86_sa)|_sub_plot_x_87_sa)|_sub_plot_x_88_sa)|_sub_plot_x_89_sa)|_sub_plot_x_90_sa)|_sub_plot_x_91_sa)|_sub_plot_x_92_sa)|_sub_plot_x_93_sa)|_sub_plot_x_94_sa)|_sub_plot_x_95_sa)|_sub_plot_x_96_sa)|_sub_plot_x_97_sa)|_sub_plot_x_98_sa)|_sub_plot_x_99_sa)|_sub_plot_x_100_sa)|_sub_plot_x_101_sa)|_sub_plot_x_102_sa)|_sub_plot_x_103_sa)|_sub_plot_x_104_sa)|_sub_plot_x_105_sa)|_sub_plot_x_106_sa)|_sub_plot_x_107_sa)|_sub_plot_x_108_sa)|_sub_plot_x_109_sa)|_sub_plot_x_110_sa)|_sub_plot_x_111_sa)|_sub_plot_x_112_sa)|_sub_plot_x_113_sa)|_sub_plot_x_114_sa)|_sub_plot_x_115_sa)|_sub_plot_x_116_sa)|_sub_plot_x_117_sa)|_sub_plot_x_118_sa)|_sub_plot_x_119_sa)|_sub_plot_x_120_sa)|_sub_plot_x_121_sa)|_sub_plot_x_122_sa)|_sub_plot_x_123_sa)|_sub_plot_x_124_sa)|_sub_plot_x_125_sa)|_sub_plot_x_126_sa)|_sub_plot_x_127_sa)|_sub_plot_x_128_sa)|_sub_plot_x_129_sa)|_sub_plot_x_130_sa)|_sub_plot_x_131_sa)|_sub_plot_x_132_sa)|_sub_plot_x_133_sa)|_sub_plot_x_134_sa)|_sub_plot_x_135_sa)|_sub_plot_x_136_sa)|_sub_plot_x_137_sa)|_sub_plot_x_138_sa)|_sub_plot_x_139_sa)|_sub_plot_x_140_sa)|_sub_plot_x_141_sa)|_sub_plot_x_142_sa)|_sub_plot_x_143_sa)|_sub_plot_x_144_sa)|_sub_plot_x_145_sa)|_sub_plot_x_146_sa)|_sub_plot_x_147_sa)|_sub_plot_x_148_sa)|_sub_plot_x_149_sa)|_sub_plot_x_150_sa)|_sub_plot_x_151_sa)|_sub_plot_x_152_sa)|_sub_plot_x_153_sa)|_sub_plot_x_154_sa)|_sub_plot_x_155_sa)|_sub_plot_x_156_sa)|_sub_plot_x_157_sa)|_sub_plot_x_158_sa)|_sub_plot_x_159_sa)|_sub_plot_x_160_sa)|_sub_plot_x_161_sa)|_sub_plot_x_162_sa)|_sub_plot_x_163_sa)|_sub_plot_x_164_sa)|_sub_plot_x_165_sa)|_sub_plot_x_166_sa)|_sub_plot_x_167_sa)|_sub_plot_x_168_sa)|_sub_plot_x_169_sa)|_sub_plot_x_170_sa)|_sub_plot_x_171_sa)|_sub_plot_x_172_sa)|_sub_plot_x_173_sa)|_sub_plot_x_174_sa)|_sub_plot_x_175_sa)|_sub_plot_x_176_sa)|_sub_plot_x_177_sa)|_sub_plot_x_178_sa)|_sub_plot_x_179_sa)|_sub_plot_x_180_sa)|_sub_plot_x_181_sa)|_sub_plot_x_182_sa)|_sub_plot_x_183_sa)|_sub_plot_x_184_sa)|_sub_plot_x_185_sa)|_sub_plot_x_186_sa)|_sub_plot_x_187_sa)|_sub_plot_x_188_sa)|_sub_plot_x_189_sa)|_sub_plot_x_190_sa)|_sub_plot_x_191_sa)|_sub_plot_x_192_sa)|_sub_plot_x_193_sa)|_sub_plot_x_194_sa)|_sub_plot_x_195_sa)|_sub_plot_x_196_sa)|_sub_plot_x_197_sa)|_sub_plot_x_198_sa)|_sub_plot_x_199_sa)|_sub_plot_x_200_sa)|_sub_plot_x_201_sa)|_sub_plot_x_202_sa)|_sub_plot_x_203_sa)|_sub_plot_x_204_sa)|_sub_plot_x_205_sa)|_sub_plot_x_206_sa)|_sub_plot_x_207_sa)|_sub_plot_x_208_sa)|_sub_plot_x_209_sa);
end
endmodule

/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Wed Dec 28 07:19:22 2022
 Licensed to :EVALUATION USER*/
