
/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 14:47:40 2023
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module meiro ( p_reset , m_clock , map_value_arg0 , map_value_arg1 , map_value_arg2 , map_value_arg3 , map_value_arg4 , map_value_arg5 , map_value_arg6 , map_value_arg7 , map_value_arg8 , map_value_arg9 , map_value_arg10 , map_value_arg11 , map_value_arg12 , map_value_arg13 , map_value_arg14 , map_value_arg15 , map_value_arg16 , map_value_arg17 , map_value_arg18 , map_value_arg19 , map_value_arg20 , map_value_arg21 , map_value_arg22 , map_value_arg23 , map_value_arg24 , map_value_arg25 , map_value_arg26 , map_value_arg27 , map_value_arg28 , map_value_arg29 , map_value_arg30 , map_value_arg31 , map_value_arg32 , map_value_arg33 , map_value_arg34 , map_value_arg35 , map_value_arg36 , map_value_arg37 , map_value_arg38 , map_value_arg39 , map_value_arg40 , map_value_arg41 , map_value_arg42 , map_value_arg43 , map_value_arg44 , map_value_arg45 , map_value_arg46 , map_value_arg47 , map_value_arg48 , map_value_arg49 , map_value_arg50 , map_value_arg51 , map_value_arg52 , map_value_arg53 , map_value_arg54 , map_value_arg55 , map_value_arg56 , map_value_arg57 , map_value_arg58 , map_value_arg59 , map_value_arg60 , map_value_arg61 , map_value_arg62 , map_value_arg63 , map_value_arg64 , map_value_arg65 , map_value_arg66 , map_value_arg67 , map_value_arg68 , map_value_arg69 , map_value_arg70 , map_value_arg71 , map_value_arg72 , map_value_arg73 , map_value_arg74 , map_value_arg75 , map_value_arg76 , map_value_arg77 , map_value_arg78 , map_value_arg79 , map_value_arg80 , map_value_arg81 , map_value_arg82 , map_value_arg83 , map_value_arg84 , map_value_arg85 , map_value_arg86 , map_value_arg87 , map_value_arg88 , map_value_arg89 , map_value_arg90 , map_value_arg91 , map_value_arg92 , map_value_arg93 , map_value_arg94 , map_value_arg95 , map_value_arg96 , map_value_arg97 , map_value_arg98 , map_value_arg99 , map_value_arg100 , map_value_arg101 , map_value_arg102 , map_value_arg103 , map_value_arg104 , map_value_arg105 , map_value_arg106 , map_value_arg107 , map_value_arg108 , map_value_arg109 , map_value_arg110 , map_value_arg111 , map_value_arg112 , map_value_arg113 , map_value_arg114 , map_value_arg115 , map_value_arg116 , map_value_arg117 , map_value_arg118 , map_value_arg119 , map_value_arg120 , map_value_arg121 , map_value_arg122 , map_value_arg123 , map_value_arg124 , map_value_arg125 , map_value_arg126 , map_value_arg127 , map_value_arg128 , map_value_arg129 , map_value_arg130 , map_value_arg131 , map_value_arg132 , map_value_arg133 , map_value_arg134 , map_value_arg135 , map_value_arg136 , map_value_arg137 , map_value_arg138 , map_value_arg139 , map_value_arg140 , map_value_arg141 , map_value_arg142 , map_value_arg143 , map_value_arg144 , map_value_arg145 , map_value_arg146 , map_value_arg147 , map_value_arg148 , map_value_arg149 , map_value_arg150 , map_value_arg151 , map_value_arg152 , map_value_arg153 , map_value_arg154 , map_value_arg155 , map_value_arg156 , map_value_arg157 , map_value_arg158 , map_value_arg159 , map_value_arg160 , map_value_arg161 , map_value_arg162 , map_value_arg163 , map_value_arg164 , map_value_arg165 , map_value_arg166 , map_value_arg167 , map_value_arg168 , map_value_arg169 , map_value_arg170 , map_value_arg171 , map_value_arg172 , map_value_arg173 , map_value_arg174 , map_value_arg175 , map_value_arg176 , map_value_arg177 , map_value_arg178 , map_value_arg179 , map_value_arg180 , map_value_arg181 , map_value_arg182 , map_value_arg183 , map_value_arg184 , map_value_arg185 , map_value_arg186 , map_value_arg187 , map_value_arg188 , map_value_arg189 , map_value_arg190 , map_value_arg191 , map_value_arg192 , map_value_arg193 , map_value_arg194 , map_value_arg195 , map_value_arg196 , map_value_arg197 , map_value_arg198 , map_value_arg199 , map_value_arg200 , map_value_arg201 , map_value_arg202 , map_value_arg203 , map_value_arg204 , map_value_arg205 , map_value_arg206 , map_value_arg207 , map_value_arg208 , map_value_arg209 , map_value_arg210 , map_value_arg211 , map_value_arg212 , map_value_arg213 , map_value_arg214 , map_value_arg215 , map_value_arg216 , map_value_arg217 , map_value_arg218 , map_value_arg219 , map_value_arg220 , map_value_arg221 , map_value_arg222 , map_value_arg223 , map_value_arg224 , map_value_arg225 , map_value_arg226 , map_value_arg227 , map_value_arg228 , map_value_arg229 , map_value_arg230 , map_value_arg231 , map_value_arg232 , map_value_arg233 , map_value_arg234 , map_value_arg235 , map_value_arg236 , map_value_arg237 , map_value_arg238 , map_value_arg239 , map_value_arg240 , map_value_arg241 , map_value_arg242 , map_value_arg243 , map_value_arg244 , map_value_arg245 , map_value_arg246 , map_value_arg247 , map_value_arg248 , map_value_arg249 , map_value_arg250 , map_value_arg251 , map_value_arg252 , map_value_arg253 , map_value_arg254 , map_value_arg255 , map_value_arg256 , map_value_arg257 , map_value_arg258 , map_value_arg259 , map_value_arg260 , map_value_arg261 , map_value_arg262 , map_value_arg263 , map_value_arg264 , map_value_arg265 , map_value_arg266 , map_value_arg267 , map_value_arg268 , map_value_arg269 , map_value_arg270 , map_value_arg271 , map_value_arg272 , map_value_arg273 , map_value_arg274 , map_value_arg275 , map_value_arg276 , map_value_arg277 , map_value_arg278 , map_value_arg279 , map_value_arg280 , map_value_arg281 , map_value_arg282 , map_value_arg283 , map_value_arg284 , map_value_arg285 , map_value_arg286 , map_value_arg287 , map_value_arg288 , map_value_arg289 , map_value_arg290 , map_value_arg291 , map_value_arg292 , map_value_arg293 , map_value_arg294 , map_value_arg295 , map_value_arg296 , map_value_arg297 , map_value_arg298 , map_value_arg299 , map_value_arg300 , map_value_arg301 , map_value_arg302 , map_value_arg303 , map_value_arg304 , map_value_arg305 , map_value_arg306 , map_value_arg307 , map_value_arg308 , map_value_arg309 , map_value_arg310 , map_value_arg311 , map_value_arg312 , map_value_arg313 , map_value_arg314 , map_value_arg315 , map_value_arg316 , map_value_arg317 , map_value_arg318 , map_value_arg319 , map_value_arg320 , map_value_arg321 , map_value_arg322 , map_value_arg323 , map_value_arg324 , map_value_arg325 , map_value_arg326 , map_value_arg327 , map_value_arg328 , map_value_arg329 , map_value_arg330 , map_value_arg331 , map_value_arg332 , map_value_arg333 , map_value_arg334 , map_value_arg335 , map_value_arg336 , map_value_arg337 , map_value_arg338 , map_value_arg339 , map_value_arg340 , map_value_arg341 , map_value_arg342 , map_value_arg343 , map_value_arg344 , map_value_arg345 , map_value_arg346 , map_value_arg347 , map_value_arg348 , map_value_arg349 , map_value_arg350 , map_value_arg351 , map_value_arg352 , map_value_arg353 , map_value_arg354 , map_value_arg355 , map_value_arg356 , map_value_arg357 , map_value_arg358 , map_value_arg359 , map_value_arg360 , map_value_arg361 , map_value_arg362 , map_value_arg363 , map_value_arg364 , map_value_arg365 , map_value_arg366 , map_value_arg367 , map_value_arg368 , map_value_arg369 , map_value_arg370 , map_value_arg371 , map_value_arg372 , map_value_arg373 , map_value_arg374 , map_value_arg375 , map_value_arg376 , map_value_arg377 , map_value_arg378 , map_value_arg379 , map_value_arg380 , map_value_arg381 , map_value_arg382 , map_value_arg383 , map_value_arg384 , map_value_arg385 , map_value_arg386 , map_value_arg387 , map_value_arg388 , map_value_arg389 , map_value_arg390 , map_value_arg391 , map_value_arg392 , map_value_arg393 , map_value_arg394 , map_value_arg395 , map_value_arg396 , map_value_arg397 , map_value_arg398 , map_value_arg399 , map_value_arg400 , map_value_arg401 , map_value_arg402 , map_value_arg403 , map_value_arg404 , map_value_arg405 , map_value_arg406 , map_value_arg407 , map_value_arg408 , map_value_arg409 , map_value_arg410 , map_value_arg411 , map_value_arg412 , map_value_arg413 , map_value_arg414 , map_value_arg415 , map_value_arg416 , map_value_arg417 , map_value_arg418 , map_value_arg419 , map_value_arg420 , map_value_arg421 , map_value_arg422 , map_value_arg423 , map_value_arg424 , map_value_arg425 , map_value_arg426 , map_value_arg427 , map_value_arg428 , map_value_arg429 , map_value_arg430 , map_value_arg431 , map_value_arg432 , map_value_arg433 , map_value_arg434 , map_value_arg435 , map_value_arg436 , map_value_arg437 , map_value_arg438 , map_value_arg439 , map_value_arg440 , map_value_arg441 , map_value_arg442 , map_value_arg443 , map_value_arg444 , map_value_arg445 , map_value_arg446 , map_value_arg447 , map_value_arg448 , map_value_arg449 , map_value_arg450 , map_value_arg451 , map_value_arg452 , map_value_arg453 , map_value_arg454 , map_value_arg455 , map_value_arg456 , map_value_arg457 , map_value_arg458 , map_value_arg459 , map_value_arg460 , map_value_arg461 , map_value_arg462 , map_value_arg463 , map_value_arg464 , map_value_arg465 , map_value_arg466 , map_value_arg467 , map_value_arg468 , map_value_arg469 , map_value_arg470 , map_value_arg471 , map_value_arg472 , map_value_arg473 , map_value_arg474 , map_value_arg475 , map_value_arg476 , map_value_arg477 , map_value_arg478 , map_value_arg479 , map_value_arg480 , map_value_arg481 , map_value_arg482 , map_value_arg483 , map_value_arg484 , map_value_arg485 , map_value_arg486 , map_value_arg487 , map_value_arg488 , map_value_arg489 , map_value_arg490 , map_value_arg491 , map_value_arg492 , map_value_arg493 , map_value_arg494 , map_value_arg495 , map_value_arg496 , map_value_arg497 , map_value_arg498 , map_value_arg499 , map_value_arg500 , map_value_arg501 , map_value_arg502 , map_value_arg503 , map_value_arg504 , map_value_arg505 , map_value_arg506 , map_value_arg507 , map_value_arg508 , map_value_arg509 , map_value_arg510 , map_value_arg511 , kekka_out0 , kekka_out1 , kekka_out2 , kekka_out3 , kekka_out4 , kekka_out5 , kekka_out6 , kekka_out7 , kekka_out8 , kekka_out9 , kekka_out10 , kekka_out11 , kekka_out12 , kekka_out13 , kekka_out14 , kekka_out15 , kekka_out16 , kekka_out17 , kekka_out18 , kekka_out19 , kekka_out20 , kekka_out21 , kekka_out22 , kekka_out23 , kekka_out24 , kekka_out25 , kekka_out26 , kekka_out27 , kekka_out28 , kekka_out29 , kekka_out30 , kekka_out31 , kekka_out32 , kekka_out33 , kekka_out34 , kekka_out35 , kekka_out36 , kekka_out37 , kekka_out38 , kekka_out39 , kekka_out40 , kekka_out41 , kekka_out42 , kekka_out43 , kekka_out44 , kekka_out45 , kekka_out46 , kekka_out47 , kekka_out48 , kekka_out49 , kekka_out50 , kekka_out51 , kekka_out52 , kekka_out53 , kekka_out54 , kekka_out55 , kekka_out56 , kekka_out57 , kekka_out58 , kekka_out59 , kekka_out60 , kekka_out61 , kekka_out62 , kekka_out63 , kekka_out64 , kekka_out65 , kekka_out66 , kekka_out67 , kekka_out68 , kekka_out69 , kekka_out70 , kekka_out71 , kekka_out72 , kekka_out73 , kekka_out74 , kekka_out75 , kekka_out76 , kekka_out77 , kekka_out78 , kekka_out79 , kekka_out80 , kekka_out81 , kekka_out82 , kekka_out83 , kekka_out84 , kekka_out85 , kekka_out86 , kekka_out87 , kekka_out88 , kekka_out89 , kekka_out90 , kekka_out91 , kekka_out92 , kekka_out93 , kekka_out94 , kekka_out95 , kekka_out96 , kekka_out97 , kekka_out98 , kekka_out99 , kekka_out100 , kekka_out101 , kekka_out102 , kekka_out103 , kekka_out104 , kekka_out105 , kekka_out106 , kekka_out107 , kekka_out108 , kekka_out109 , kekka_out110 , kekka_out111 , kekka_out112 , kekka_out113 , kekka_out114 , kekka_out115 , kekka_out116 , kekka_out117 , kekka_out118 , kekka_out119 , kekka_out120 , kekka_out121 , kekka_out122 , kekka_out123 , kekka_out124 , kekka_out125 , kekka_out126 , kekka_out127 , kekka_out128 , kekka_out129 , kekka_out130 , kekka_out131 , kekka_out132 , kekka_out133 , kekka_out134 , kekka_out135 , kekka_out136 , kekka_out137 , kekka_out138 , kekka_out139 , kekka_out140 , kekka_out141 , kekka_out142 , kekka_out143 , kekka_out144 , kekka_out145 , kekka_out146 , kekka_out147 , kekka_out148 , kekka_out149 , kekka_out150 , kekka_out151 , kekka_out152 , kekka_out153 , kekka_out154 , kekka_out155 , kekka_out156 , kekka_out157 , kekka_out158 , kekka_out159 , kekka_out160 , kekka_out161 , kekka_out162 , kekka_out163 , kekka_out164 , kekka_out165 , kekka_out166 , kekka_out167 , kekka_out168 , kekka_out169 , kekka_out170 , kekka_out171 , kekka_out172 , kekka_out173 , kekka_out174 , kekka_out175 , kekka_out176 , kekka_out177 , kekka_out178 , kekka_out179 , kekka_out180 , kekka_out181 , kekka_out182 , kekka_out183 , kekka_out184 , kekka_out185 , kekka_out186 , kekka_out187 , kekka_out188 , kekka_out189 , kekka_out190 , kekka_out191 , kekka_out192 , kekka_out193 , kekka_out194 , kekka_out195 , kekka_out196 , kekka_out197 , kekka_out198 , kekka_out199 , kekka_out200 , kekka_out201 , kekka_out202 , kekka_out203 , kekka_out204 , kekka_out205 , kekka_out206 , kekka_out207 , kekka_out208 , kekka_out209 , kekka_out210 , kekka_out211 , kekka_out212 , kekka_out213 , kekka_out214 , kekka_out215 , kekka_out216 , kekka_out217 , kekka_out218 , kekka_out219 , kekka_out220 , kekka_out221 , kekka_out222 , in_do , end_meiro );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input [9:0] map_value_arg0;
  wire [9:0] map_value_arg0;
  input [9:0] map_value_arg1;
  wire [9:0] map_value_arg1;
  input [9:0] map_value_arg2;
  wire [9:0] map_value_arg2;
  input [9:0] map_value_arg3;
  wire [9:0] map_value_arg3;
  input [9:0] map_value_arg4;
  wire [9:0] map_value_arg4;
  input [9:0] map_value_arg5;
  wire [9:0] map_value_arg5;
  input [9:0] map_value_arg6;
  wire [9:0] map_value_arg6;
  input [9:0] map_value_arg7;
  wire [9:0] map_value_arg7;
  input [9:0] map_value_arg8;
  wire [9:0] map_value_arg8;
  input [9:0] map_value_arg9;
  wire [9:0] map_value_arg9;
  input [9:0] map_value_arg10;
  wire [9:0] map_value_arg10;
  input [9:0] map_value_arg11;
  wire [9:0] map_value_arg11;
  input [9:0] map_value_arg12;
  wire [9:0] map_value_arg12;
  input [9:0] map_value_arg13;
  wire [9:0] map_value_arg13;
  input [9:0] map_value_arg14;
  wire [9:0] map_value_arg14;
  input [9:0] map_value_arg15;
  wire [9:0] map_value_arg15;
  input [9:0] map_value_arg16;
  wire [9:0] map_value_arg16;
  input [9:0] map_value_arg17;
  wire [9:0] map_value_arg17;
  input [9:0] map_value_arg18;
  wire [9:0] map_value_arg18;
  input [9:0] map_value_arg19;
  wire [9:0] map_value_arg19;
  input [9:0] map_value_arg20;
  wire [9:0] map_value_arg20;
  input [9:0] map_value_arg21;
  wire [9:0] map_value_arg21;
  input [9:0] map_value_arg22;
  wire [9:0] map_value_arg22;
  input [9:0] map_value_arg23;
  wire [9:0] map_value_arg23;
  input [9:0] map_value_arg24;
  wire [9:0] map_value_arg24;
  input [9:0] map_value_arg25;
  wire [9:0] map_value_arg25;
  input [9:0] map_value_arg26;
  wire [9:0] map_value_arg26;
  input [9:0] map_value_arg27;
  wire [9:0] map_value_arg27;
  input [9:0] map_value_arg28;
  wire [9:0] map_value_arg28;
  input [9:0] map_value_arg29;
  wire [9:0] map_value_arg29;
  input [9:0] map_value_arg30;
  wire [9:0] map_value_arg30;
  input [9:0] map_value_arg31;
  wire [9:0] map_value_arg31;
  input [9:0] map_value_arg32;
  wire [9:0] map_value_arg32;
  input [9:0] map_value_arg33;
  wire [9:0] map_value_arg33;
  input [9:0] map_value_arg34;
  wire [9:0] map_value_arg34;
  input [9:0] map_value_arg35;
  wire [9:0] map_value_arg35;
  input [9:0] map_value_arg36;
  wire [9:0] map_value_arg36;
  input [9:0] map_value_arg37;
  wire [9:0] map_value_arg37;
  input [9:0] map_value_arg38;
  wire [9:0] map_value_arg38;
  input [9:0] map_value_arg39;
  wire [9:0] map_value_arg39;
  input [9:0] map_value_arg40;
  wire [9:0] map_value_arg40;
  input [9:0] map_value_arg41;
  wire [9:0] map_value_arg41;
  input [9:0] map_value_arg42;
  wire [9:0] map_value_arg42;
  input [9:0] map_value_arg43;
  wire [9:0] map_value_arg43;
  input [9:0] map_value_arg44;
  wire [9:0] map_value_arg44;
  input [9:0] map_value_arg45;
  wire [9:0] map_value_arg45;
  input [9:0] map_value_arg46;
  wire [9:0] map_value_arg46;
  input [9:0] map_value_arg47;
  wire [9:0] map_value_arg47;
  input [9:0] map_value_arg48;
  wire [9:0] map_value_arg48;
  input [9:0] map_value_arg49;
  wire [9:0] map_value_arg49;
  input [9:0] map_value_arg50;
  wire [9:0] map_value_arg50;
  input [9:0] map_value_arg51;
  wire [9:0] map_value_arg51;
  input [9:0] map_value_arg52;
  wire [9:0] map_value_arg52;
  input [9:0] map_value_arg53;
  wire [9:0] map_value_arg53;
  input [9:0] map_value_arg54;
  wire [9:0] map_value_arg54;
  input [9:0] map_value_arg55;
  wire [9:0] map_value_arg55;
  input [9:0] map_value_arg56;
  wire [9:0] map_value_arg56;
  input [9:0] map_value_arg57;
  wire [9:0] map_value_arg57;
  input [9:0] map_value_arg58;
  wire [9:0] map_value_arg58;
  input [9:0] map_value_arg59;
  wire [9:0] map_value_arg59;
  input [9:0] map_value_arg60;
  wire [9:0] map_value_arg60;
  input [9:0] map_value_arg61;
  wire [9:0] map_value_arg61;
  input [9:0] map_value_arg62;
  wire [9:0] map_value_arg62;
  input [9:0] map_value_arg63;
  wire [9:0] map_value_arg63;
  input [9:0] map_value_arg64;
  wire [9:0] map_value_arg64;
  input [9:0] map_value_arg65;
  wire [9:0] map_value_arg65;
  input [9:0] map_value_arg66;
  wire [9:0] map_value_arg66;
  input [9:0] map_value_arg67;
  wire [9:0] map_value_arg67;
  input [9:0] map_value_arg68;
  wire [9:0] map_value_arg68;
  input [9:0] map_value_arg69;
  wire [9:0] map_value_arg69;
  input [9:0] map_value_arg70;
  wire [9:0] map_value_arg70;
  input [9:0] map_value_arg71;
  wire [9:0] map_value_arg71;
  input [9:0] map_value_arg72;
  wire [9:0] map_value_arg72;
  input [9:0] map_value_arg73;
  wire [9:0] map_value_arg73;
  input [9:0] map_value_arg74;
  wire [9:0] map_value_arg74;
  input [9:0] map_value_arg75;
  wire [9:0] map_value_arg75;
  input [9:0] map_value_arg76;
  wire [9:0] map_value_arg76;
  input [9:0] map_value_arg77;
  wire [9:0] map_value_arg77;
  input [9:0] map_value_arg78;
  wire [9:0] map_value_arg78;
  input [9:0] map_value_arg79;
  wire [9:0] map_value_arg79;
  input [9:0] map_value_arg80;
  wire [9:0] map_value_arg80;
  input [9:0] map_value_arg81;
  wire [9:0] map_value_arg81;
  input [9:0] map_value_arg82;
  wire [9:0] map_value_arg82;
  input [9:0] map_value_arg83;
  wire [9:0] map_value_arg83;
  input [9:0] map_value_arg84;
  wire [9:0] map_value_arg84;
  input [9:0] map_value_arg85;
  wire [9:0] map_value_arg85;
  input [9:0] map_value_arg86;
  wire [9:0] map_value_arg86;
  input [9:0] map_value_arg87;
  wire [9:0] map_value_arg87;
  input [9:0] map_value_arg88;
  wire [9:0] map_value_arg88;
  input [9:0] map_value_arg89;
  wire [9:0] map_value_arg89;
  input [9:0] map_value_arg90;
  wire [9:0] map_value_arg90;
  input [9:0] map_value_arg91;
  wire [9:0] map_value_arg91;
  input [9:0] map_value_arg92;
  wire [9:0] map_value_arg92;
  input [9:0] map_value_arg93;
  wire [9:0] map_value_arg93;
  input [9:0] map_value_arg94;
  wire [9:0] map_value_arg94;
  input [9:0] map_value_arg95;
  wire [9:0] map_value_arg95;
  input [9:0] map_value_arg96;
  wire [9:0] map_value_arg96;
  input [9:0] map_value_arg97;
  wire [9:0] map_value_arg97;
  input [9:0] map_value_arg98;
  wire [9:0] map_value_arg98;
  input [9:0] map_value_arg99;
  wire [9:0] map_value_arg99;
  input [9:0] map_value_arg100;
  wire [9:0] map_value_arg100;
  input [9:0] map_value_arg101;
  wire [9:0] map_value_arg101;
  input [9:0] map_value_arg102;
  wire [9:0] map_value_arg102;
  input [9:0] map_value_arg103;
  wire [9:0] map_value_arg103;
  input [9:0] map_value_arg104;
  wire [9:0] map_value_arg104;
  input [9:0] map_value_arg105;
  wire [9:0] map_value_arg105;
  input [9:0] map_value_arg106;
  wire [9:0] map_value_arg106;
  input [9:0] map_value_arg107;
  wire [9:0] map_value_arg107;
  input [9:0] map_value_arg108;
  wire [9:0] map_value_arg108;
  input [9:0] map_value_arg109;
  wire [9:0] map_value_arg109;
  input [9:0] map_value_arg110;
  wire [9:0] map_value_arg110;
  input [9:0] map_value_arg111;
  wire [9:0] map_value_arg111;
  input [9:0] map_value_arg112;
  wire [9:0] map_value_arg112;
  input [9:0] map_value_arg113;
  wire [9:0] map_value_arg113;
  input [9:0] map_value_arg114;
  wire [9:0] map_value_arg114;
  input [9:0] map_value_arg115;
  wire [9:0] map_value_arg115;
  input [9:0] map_value_arg116;
  wire [9:0] map_value_arg116;
  input [9:0] map_value_arg117;
  wire [9:0] map_value_arg117;
  input [9:0] map_value_arg118;
  wire [9:0] map_value_arg118;
  input [9:0] map_value_arg119;
  wire [9:0] map_value_arg119;
  input [9:0] map_value_arg120;
  wire [9:0] map_value_arg120;
  input [9:0] map_value_arg121;
  wire [9:0] map_value_arg121;
  input [9:0] map_value_arg122;
  wire [9:0] map_value_arg122;
  input [9:0] map_value_arg123;
  wire [9:0] map_value_arg123;
  input [9:0] map_value_arg124;
  wire [9:0] map_value_arg124;
  input [9:0] map_value_arg125;
  wire [9:0] map_value_arg125;
  input [9:0] map_value_arg126;
  wire [9:0] map_value_arg126;
  input [9:0] map_value_arg127;
  wire [9:0] map_value_arg127;
  input [9:0] map_value_arg128;
  wire [9:0] map_value_arg128;
  input [9:0] map_value_arg129;
  wire [9:0] map_value_arg129;
  input [9:0] map_value_arg130;
  wire [9:0] map_value_arg130;
  input [9:0] map_value_arg131;
  wire [9:0] map_value_arg131;
  input [9:0] map_value_arg132;
  wire [9:0] map_value_arg132;
  input [9:0] map_value_arg133;
  wire [9:0] map_value_arg133;
  input [9:0] map_value_arg134;
  wire [9:0] map_value_arg134;
  input [9:0] map_value_arg135;
  wire [9:0] map_value_arg135;
  input [9:0] map_value_arg136;
  wire [9:0] map_value_arg136;
  input [9:0] map_value_arg137;
  wire [9:0] map_value_arg137;
  input [9:0] map_value_arg138;
  wire [9:0] map_value_arg138;
  input [9:0] map_value_arg139;
  wire [9:0] map_value_arg139;
  input [9:0] map_value_arg140;
  wire [9:0] map_value_arg140;
  input [9:0] map_value_arg141;
  wire [9:0] map_value_arg141;
  input [9:0] map_value_arg142;
  wire [9:0] map_value_arg142;
  input [9:0] map_value_arg143;
  wire [9:0] map_value_arg143;
  input [9:0] map_value_arg144;
  wire [9:0] map_value_arg144;
  input [9:0] map_value_arg145;
  wire [9:0] map_value_arg145;
  input [9:0] map_value_arg146;
  wire [9:0] map_value_arg146;
  input [9:0] map_value_arg147;
  wire [9:0] map_value_arg147;
  input [9:0] map_value_arg148;
  wire [9:0] map_value_arg148;
  input [9:0] map_value_arg149;
  wire [9:0] map_value_arg149;
  input [9:0] map_value_arg150;
  wire [9:0] map_value_arg150;
  input [9:0] map_value_arg151;
  wire [9:0] map_value_arg151;
  input [9:0] map_value_arg152;
  wire [9:0] map_value_arg152;
  input [9:0] map_value_arg153;
  wire [9:0] map_value_arg153;
  input [9:0] map_value_arg154;
  wire [9:0] map_value_arg154;
  input [9:0] map_value_arg155;
  wire [9:0] map_value_arg155;
  input [9:0] map_value_arg156;
  wire [9:0] map_value_arg156;
  input [9:0] map_value_arg157;
  wire [9:0] map_value_arg157;
  input [9:0] map_value_arg158;
  wire [9:0] map_value_arg158;
  input [9:0] map_value_arg159;
  wire [9:0] map_value_arg159;
  input [9:0] map_value_arg160;
  wire [9:0] map_value_arg160;
  input [9:0] map_value_arg161;
  wire [9:0] map_value_arg161;
  input [9:0] map_value_arg162;
  wire [9:0] map_value_arg162;
  input [9:0] map_value_arg163;
  wire [9:0] map_value_arg163;
  input [9:0] map_value_arg164;
  wire [9:0] map_value_arg164;
  input [9:0] map_value_arg165;
  wire [9:0] map_value_arg165;
  input [9:0] map_value_arg166;
  wire [9:0] map_value_arg166;
  input [9:0] map_value_arg167;
  wire [9:0] map_value_arg167;
  input [9:0] map_value_arg168;
  wire [9:0] map_value_arg168;
  input [9:0] map_value_arg169;
  wire [9:0] map_value_arg169;
  input [9:0] map_value_arg170;
  wire [9:0] map_value_arg170;
  input [9:0] map_value_arg171;
  wire [9:0] map_value_arg171;
  input [9:0] map_value_arg172;
  wire [9:0] map_value_arg172;
  input [9:0] map_value_arg173;
  wire [9:0] map_value_arg173;
  input [9:0] map_value_arg174;
  wire [9:0] map_value_arg174;
  input [9:0] map_value_arg175;
  wire [9:0] map_value_arg175;
  input [9:0] map_value_arg176;
  wire [9:0] map_value_arg176;
  input [9:0] map_value_arg177;
  wire [9:0] map_value_arg177;
  input [9:0] map_value_arg178;
  wire [9:0] map_value_arg178;
  input [9:0] map_value_arg179;
  wire [9:0] map_value_arg179;
  input [9:0] map_value_arg180;
  wire [9:0] map_value_arg180;
  input [9:0] map_value_arg181;
  wire [9:0] map_value_arg181;
  input [9:0] map_value_arg182;
  wire [9:0] map_value_arg182;
  input [9:0] map_value_arg183;
  wire [9:0] map_value_arg183;
  input [9:0] map_value_arg184;
  wire [9:0] map_value_arg184;
  input [9:0] map_value_arg185;
  wire [9:0] map_value_arg185;
  input [9:0] map_value_arg186;
  wire [9:0] map_value_arg186;
  input [9:0] map_value_arg187;
  wire [9:0] map_value_arg187;
  input [9:0] map_value_arg188;
  wire [9:0] map_value_arg188;
  input [9:0] map_value_arg189;
  wire [9:0] map_value_arg189;
  input [9:0] map_value_arg190;
  wire [9:0] map_value_arg190;
  input [9:0] map_value_arg191;
  wire [9:0] map_value_arg191;
  input [9:0] map_value_arg192;
  wire [9:0] map_value_arg192;
  input [9:0] map_value_arg193;
  wire [9:0] map_value_arg193;
  input [9:0] map_value_arg194;
  wire [9:0] map_value_arg194;
  input [9:0] map_value_arg195;
  wire [9:0] map_value_arg195;
  input [9:0] map_value_arg196;
  wire [9:0] map_value_arg196;
  input [9:0] map_value_arg197;
  wire [9:0] map_value_arg197;
  input [9:0] map_value_arg198;
  wire [9:0] map_value_arg198;
  input [9:0] map_value_arg199;
  wire [9:0] map_value_arg199;
  input [9:0] map_value_arg200;
  wire [9:0] map_value_arg200;
  input [9:0] map_value_arg201;
  wire [9:0] map_value_arg201;
  input [9:0] map_value_arg202;
  wire [9:0] map_value_arg202;
  input [9:0] map_value_arg203;
  wire [9:0] map_value_arg203;
  input [9:0] map_value_arg204;
  wire [9:0] map_value_arg204;
  input [9:0] map_value_arg205;
  wire [9:0] map_value_arg205;
  input [9:0] map_value_arg206;
  wire [9:0] map_value_arg206;
  input [9:0] map_value_arg207;
  wire [9:0] map_value_arg207;
  input [9:0] map_value_arg208;
  wire [9:0] map_value_arg208;
  input [9:0] map_value_arg209;
  wire [9:0] map_value_arg209;
  input [9:0] map_value_arg210;
  wire [9:0] map_value_arg210;
  input [9:0] map_value_arg211;
  wire [9:0] map_value_arg211;
  input [9:0] map_value_arg212;
  wire [9:0] map_value_arg212;
  input [9:0] map_value_arg213;
  wire [9:0] map_value_arg213;
  input [9:0] map_value_arg214;
  wire [9:0] map_value_arg214;
  input [9:0] map_value_arg215;
  wire [9:0] map_value_arg215;
  input [9:0] map_value_arg216;
  wire [9:0] map_value_arg216;
  input [9:0] map_value_arg217;
  wire [9:0] map_value_arg217;
  input [9:0] map_value_arg218;
  wire [9:0] map_value_arg218;
  input [9:0] map_value_arg219;
  wire [9:0] map_value_arg219;
  input [9:0] map_value_arg220;
  wire [9:0] map_value_arg220;
  input [9:0] map_value_arg221;
  wire [9:0] map_value_arg221;
  input [9:0] map_value_arg222;
  wire [9:0] map_value_arg222;
  input [9:0] map_value_arg223;
  wire [9:0] map_value_arg223;
  input [9:0] map_value_arg224;
  wire [9:0] map_value_arg224;
  input [9:0] map_value_arg225;
  wire [9:0] map_value_arg225;
  input [9:0] map_value_arg226;
  wire [9:0] map_value_arg226;
  input [9:0] map_value_arg227;
  wire [9:0] map_value_arg227;
  input [9:0] map_value_arg228;
  wire [9:0] map_value_arg228;
  input [9:0] map_value_arg229;
  wire [9:0] map_value_arg229;
  input [9:0] map_value_arg230;
  wire [9:0] map_value_arg230;
  input [9:0] map_value_arg231;
  wire [9:0] map_value_arg231;
  input [9:0] map_value_arg232;
  wire [9:0] map_value_arg232;
  input [9:0] map_value_arg233;
  wire [9:0] map_value_arg233;
  input [9:0] map_value_arg234;
  wire [9:0] map_value_arg234;
  input [9:0] map_value_arg235;
  wire [9:0] map_value_arg235;
  input [9:0] map_value_arg236;
  wire [9:0] map_value_arg236;
  input [9:0] map_value_arg237;
  wire [9:0] map_value_arg237;
  input [9:0] map_value_arg238;
  wire [9:0] map_value_arg238;
  input [9:0] map_value_arg239;
  wire [9:0] map_value_arg239;
  input [9:0] map_value_arg240;
  wire [9:0] map_value_arg240;
  input [9:0] map_value_arg241;
  wire [9:0] map_value_arg241;
  input [9:0] map_value_arg242;
  wire [9:0] map_value_arg242;
  input [9:0] map_value_arg243;
  wire [9:0] map_value_arg243;
  input [9:0] map_value_arg244;
  wire [9:0] map_value_arg244;
  input [9:0] map_value_arg245;
  wire [9:0] map_value_arg245;
  input [9:0] map_value_arg246;
  wire [9:0] map_value_arg246;
  input [9:0] map_value_arg247;
  wire [9:0] map_value_arg247;
  input [9:0] map_value_arg248;
  wire [9:0] map_value_arg248;
  input [9:0] map_value_arg249;
  wire [9:0] map_value_arg249;
  input [9:0] map_value_arg250;
  wire [9:0] map_value_arg250;
  input [9:0] map_value_arg251;
  wire [9:0] map_value_arg251;
  input [9:0] map_value_arg252;
  wire [9:0] map_value_arg252;
  input [9:0] map_value_arg253;
  wire [9:0] map_value_arg253;
  input [9:0] map_value_arg254;
  wire [9:0] map_value_arg254;
  input [9:0] map_value_arg255;
  wire [9:0] map_value_arg255;
  input [9:0] map_value_arg256;
  wire [9:0] map_value_arg256;
  input [9:0] map_value_arg257;
  wire [9:0] map_value_arg257;
  input [9:0] map_value_arg258;
  wire [9:0] map_value_arg258;
  input [9:0] map_value_arg259;
  wire [9:0] map_value_arg259;
  input [9:0] map_value_arg260;
  wire [9:0] map_value_arg260;
  input [9:0] map_value_arg261;
  wire [9:0] map_value_arg261;
  input [9:0] map_value_arg262;
  wire [9:0] map_value_arg262;
  input [9:0] map_value_arg263;
  wire [9:0] map_value_arg263;
  input [9:0] map_value_arg264;
  wire [9:0] map_value_arg264;
  input [9:0] map_value_arg265;
  wire [9:0] map_value_arg265;
  input [9:0] map_value_arg266;
  wire [9:0] map_value_arg266;
  input [9:0] map_value_arg267;
  wire [9:0] map_value_arg267;
  input [9:0] map_value_arg268;
  wire [9:0] map_value_arg268;
  input [9:0] map_value_arg269;
  wire [9:0] map_value_arg269;
  input [9:0] map_value_arg270;
  wire [9:0] map_value_arg270;
  input [9:0] map_value_arg271;
  wire [9:0] map_value_arg271;
  input [9:0] map_value_arg272;
  wire [9:0] map_value_arg272;
  input [9:0] map_value_arg273;
  wire [9:0] map_value_arg273;
  input [9:0] map_value_arg274;
  wire [9:0] map_value_arg274;
  input [9:0] map_value_arg275;
  wire [9:0] map_value_arg275;
  input [9:0] map_value_arg276;
  wire [9:0] map_value_arg276;
  input [9:0] map_value_arg277;
  wire [9:0] map_value_arg277;
  input [9:0] map_value_arg278;
  wire [9:0] map_value_arg278;
  input [9:0] map_value_arg279;
  wire [9:0] map_value_arg279;
  input [9:0] map_value_arg280;
  wire [9:0] map_value_arg280;
  input [9:0] map_value_arg281;
  wire [9:0] map_value_arg281;
  input [9:0] map_value_arg282;
  wire [9:0] map_value_arg282;
  input [9:0] map_value_arg283;
  wire [9:0] map_value_arg283;
  input [9:0] map_value_arg284;
  wire [9:0] map_value_arg284;
  input [9:0] map_value_arg285;
  wire [9:0] map_value_arg285;
  input [9:0] map_value_arg286;
  wire [9:0] map_value_arg286;
  input [9:0] map_value_arg287;
  wire [9:0] map_value_arg287;
  input [9:0] map_value_arg288;
  wire [9:0] map_value_arg288;
  input [9:0] map_value_arg289;
  wire [9:0] map_value_arg289;
  input [9:0] map_value_arg290;
  wire [9:0] map_value_arg290;
  input [9:0] map_value_arg291;
  wire [9:0] map_value_arg291;
  input [9:0] map_value_arg292;
  wire [9:0] map_value_arg292;
  input [9:0] map_value_arg293;
  wire [9:0] map_value_arg293;
  input [9:0] map_value_arg294;
  wire [9:0] map_value_arg294;
  input [9:0] map_value_arg295;
  wire [9:0] map_value_arg295;
  input [9:0] map_value_arg296;
  wire [9:0] map_value_arg296;
  input [9:0] map_value_arg297;
  wire [9:0] map_value_arg297;
  input [9:0] map_value_arg298;
  wire [9:0] map_value_arg298;
  input [9:0] map_value_arg299;
  wire [9:0] map_value_arg299;
  input [9:0] map_value_arg300;
  wire [9:0] map_value_arg300;
  input [9:0] map_value_arg301;
  wire [9:0] map_value_arg301;
  input [9:0] map_value_arg302;
  wire [9:0] map_value_arg302;
  input [9:0] map_value_arg303;
  wire [9:0] map_value_arg303;
  input [9:0] map_value_arg304;
  wire [9:0] map_value_arg304;
  input [9:0] map_value_arg305;
  wire [9:0] map_value_arg305;
  input [9:0] map_value_arg306;
  wire [9:0] map_value_arg306;
  input [9:0] map_value_arg307;
  wire [9:0] map_value_arg307;
  input [9:0] map_value_arg308;
  wire [9:0] map_value_arg308;
  input [9:0] map_value_arg309;
  wire [9:0] map_value_arg309;
  input [9:0] map_value_arg310;
  wire [9:0] map_value_arg310;
  input [9:0] map_value_arg311;
  wire [9:0] map_value_arg311;
  input [9:0] map_value_arg312;
  wire [9:0] map_value_arg312;
  input [9:0] map_value_arg313;
  wire [9:0] map_value_arg313;
  input [9:0] map_value_arg314;
  wire [9:0] map_value_arg314;
  input [9:0] map_value_arg315;
  wire [9:0] map_value_arg315;
  input [9:0] map_value_arg316;
  wire [9:0] map_value_arg316;
  input [9:0] map_value_arg317;
  wire [9:0] map_value_arg317;
  input [9:0] map_value_arg318;
  wire [9:0] map_value_arg318;
  input [9:0] map_value_arg319;
  wire [9:0] map_value_arg319;
  input [9:0] map_value_arg320;
  wire [9:0] map_value_arg320;
  input [9:0] map_value_arg321;
  wire [9:0] map_value_arg321;
  input [9:0] map_value_arg322;
  wire [9:0] map_value_arg322;
  input [9:0] map_value_arg323;
  wire [9:0] map_value_arg323;
  input [9:0] map_value_arg324;
  wire [9:0] map_value_arg324;
  input [9:0] map_value_arg325;
  wire [9:0] map_value_arg325;
  input [9:0] map_value_arg326;
  wire [9:0] map_value_arg326;
  input [9:0] map_value_arg327;
  wire [9:0] map_value_arg327;
  input [9:0] map_value_arg328;
  wire [9:0] map_value_arg328;
  input [9:0] map_value_arg329;
  wire [9:0] map_value_arg329;
  input [9:0] map_value_arg330;
  wire [9:0] map_value_arg330;
  input [9:0] map_value_arg331;
  wire [9:0] map_value_arg331;
  input [9:0] map_value_arg332;
  wire [9:0] map_value_arg332;
  input [9:0] map_value_arg333;
  wire [9:0] map_value_arg333;
  input [9:0] map_value_arg334;
  wire [9:0] map_value_arg334;
  input [9:0] map_value_arg335;
  wire [9:0] map_value_arg335;
  input [9:0] map_value_arg336;
  wire [9:0] map_value_arg336;
  input [9:0] map_value_arg337;
  wire [9:0] map_value_arg337;
  input [9:0] map_value_arg338;
  wire [9:0] map_value_arg338;
  input [9:0] map_value_arg339;
  wire [9:0] map_value_arg339;
  input [9:0] map_value_arg340;
  wire [9:0] map_value_arg340;
  input [9:0] map_value_arg341;
  wire [9:0] map_value_arg341;
  input [9:0] map_value_arg342;
  wire [9:0] map_value_arg342;
  input [9:0] map_value_arg343;
  wire [9:0] map_value_arg343;
  input [9:0] map_value_arg344;
  wire [9:0] map_value_arg344;
  input [9:0] map_value_arg345;
  wire [9:0] map_value_arg345;
  input [9:0] map_value_arg346;
  wire [9:0] map_value_arg346;
  input [9:0] map_value_arg347;
  wire [9:0] map_value_arg347;
  input [9:0] map_value_arg348;
  wire [9:0] map_value_arg348;
  input [9:0] map_value_arg349;
  wire [9:0] map_value_arg349;
  input [9:0] map_value_arg350;
  wire [9:0] map_value_arg350;
  input [9:0] map_value_arg351;
  wire [9:0] map_value_arg351;
  input [9:0] map_value_arg352;
  wire [9:0] map_value_arg352;
  input [9:0] map_value_arg353;
  wire [9:0] map_value_arg353;
  input [9:0] map_value_arg354;
  wire [9:0] map_value_arg354;
  input [9:0] map_value_arg355;
  wire [9:0] map_value_arg355;
  input [9:0] map_value_arg356;
  wire [9:0] map_value_arg356;
  input [9:0] map_value_arg357;
  wire [9:0] map_value_arg357;
  input [9:0] map_value_arg358;
  wire [9:0] map_value_arg358;
  input [9:0] map_value_arg359;
  wire [9:0] map_value_arg359;
  input [9:0] map_value_arg360;
  wire [9:0] map_value_arg360;
  input [9:0] map_value_arg361;
  wire [9:0] map_value_arg361;
  input [9:0] map_value_arg362;
  wire [9:0] map_value_arg362;
  input [9:0] map_value_arg363;
  wire [9:0] map_value_arg363;
  input [9:0] map_value_arg364;
  wire [9:0] map_value_arg364;
  input [9:0] map_value_arg365;
  wire [9:0] map_value_arg365;
  input [9:0] map_value_arg366;
  wire [9:0] map_value_arg366;
  input [9:0] map_value_arg367;
  wire [9:0] map_value_arg367;
  input [9:0] map_value_arg368;
  wire [9:0] map_value_arg368;
  input [9:0] map_value_arg369;
  wire [9:0] map_value_arg369;
  input [9:0] map_value_arg370;
  wire [9:0] map_value_arg370;
  input [9:0] map_value_arg371;
  wire [9:0] map_value_arg371;
  input [9:0] map_value_arg372;
  wire [9:0] map_value_arg372;
  input [9:0] map_value_arg373;
  wire [9:0] map_value_arg373;
  input [9:0] map_value_arg374;
  wire [9:0] map_value_arg374;
  input [9:0] map_value_arg375;
  wire [9:0] map_value_arg375;
  input [9:0] map_value_arg376;
  wire [9:0] map_value_arg376;
  input [9:0] map_value_arg377;
  wire [9:0] map_value_arg377;
  input [9:0] map_value_arg378;
  wire [9:0] map_value_arg378;
  input [9:0] map_value_arg379;
  wire [9:0] map_value_arg379;
  input [9:0] map_value_arg380;
  wire [9:0] map_value_arg380;
  input [9:0] map_value_arg381;
  wire [9:0] map_value_arg381;
  input [9:0] map_value_arg382;
  wire [9:0] map_value_arg382;
  input [9:0] map_value_arg383;
  wire [9:0] map_value_arg383;
  input [9:0] map_value_arg384;
  wire [9:0] map_value_arg384;
  input [9:0] map_value_arg385;
  wire [9:0] map_value_arg385;
  input [9:0] map_value_arg386;
  wire [9:0] map_value_arg386;
  input [9:0] map_value_arg387;
  wire [9:0] map_value_arg387;
  input [9:0] map_value_arg388;
  wire [9:0] map_value_arg388;
  input [9:0] map_value_arg389;
  wire [9:0] map_value_arg389;
  input [9:0] map_value_arg390;
  wire [9:0] map_value_arg390;
  input [9:0] map_value_arg391;
  wire [9:0] map_value_arg391;
  input [9:0] map_value_arg392;
  wire [9:0] map_value_arg392;
  input [9:0] map_value_arg393;
  wire [9:0] map_value_arg393;
  input [9:0] map_value_arg394;
  wire [9:0] map_value_arg394;
  input [9:0] map_value_arg395;
  wire [9:0] map_value_arg395;
  input [9:0] map_value_arg396;
  wire [9:0] map_value_arg396;
  input [9:0] map_value_arg397;
  wire [9:0] map_value_arg397;
  input [9:0] map_value_arg398;
  wire [9:0] map_value_arg398;
  input [9:0] map_value_arg399;
  wire [9:0] map_value_arg399;
  input [9:0] map_value_arg400;
  wire [9:0] map_value_arg400;
  input [9:0] map_value_arg401;
  wire [9:0] map_value_arg401;
  input [9:0] map_value_arg402;
  wire [9:0] map_value_arg402;
  input [9:0] map_value_arg403;
  wire [9:0] map_value_arg403;
  input [9:0] map_value_arg404;
  wire [9:0] map_value_arg404;
  input [9:0] map_value_arg405;
  wire [9:0] map_value_arg405;
  input [9:0] map_value_arg406;
  wire [9:0] map_value_arg406;
  input [9:0] map_value_arg407;
  wire [9:0] map_value_arg407;
  input [9:0] map_value_arg408;
  wire [9:0] map_value_arg408;
  input [9:0] map_value_arg409;
  wire [9:0] map_value_arg409;
  input [9:0] map_value_arg410;
  wire [9:0] map_value_arg410;
  input [9:0] map_value_arg411;
  wire [9:0] map_value_arg411;
  input [9:0] map_value_arg412;
  wire [9:0] map_value_arg412;
  input [9:0] map_value_arg413;
  wire [9:0] map_value_arg413;
  input [9:0] map_value_arg414;
  wire [9:0] map_value_arg414;
  input [9:0] map_value_arg415;
  wire [9:0] map_value_arg415;
  input [9:0] map_value_arg416;
  wire [9:0] map_value_arg416;
  input [9:0] map_value_arg417;
  wire [9:0] map_value_arg417;
  input [9:0] map_value_arg418;
  wire [9:0] map_value_arg418;
  input [9:0] map_value_arg419;
  wire [9:0] map_value_arg419;
  input [9:0] map_value_arg420;
  wire [9:0] map_value_arg420;
  input [9:0] map_value_arg421;
  wire [9:0] map_value_arg421;
  input [9:0] map_value_arg422;
  wire [9:0] map_value_arg422;
  input [9:0] map_value_arg423;
  wire [9:0] map_value_arg423;
  input [9:0] map_value_arg424;
  wire [9:0] map_value_arg424;
  input [9:0] map_value_arg425;
  wire [9:0] map_value_arg425;
  input [9:0] map_value_arg426;
  wire [9:0] map_value_arg426;
  input [9:0] map_value_arg427;
  wire [9:0] map_value_arg427;
  input [9:0] map_value_arg428;
  wire [9:0] map_value_arg428;
  input [9:0] map_value_arg429;
  wire [9:0] map_value_arg429;
  input [9:0] map_value_arg430;
  wire [9:0] map_value_arg430;
  input [9:0] map_value_arg431;
  wire [9:0] map_value_arg431;
  input [9:0] map_value_arg432;
  wire [9:0] map_value_arg432;
  input [9:0] map_value_arg433;
  wire [9:0] map_value_arg433;
  input [9:0] map_value_arg434;
  wire [9:0] map_value_arg434;
  input [9:0] map_value_arg435;
  wire [9:0] map_value_arg435;
  input [9:0] map_value_arg436;
  wire [9:0] map_value_arg436;
  input [9:0] map_value_arg437;
  wire [9:0] map_value_arg437;
  input [9:0] map_value_arg438;
  wire [9:0] map_value_arg438;
  input [9:0] map_value_arg439;
  wire [9:0] map_value_arg439;
  input [9:0] map_value_arg440;
  wire [9:0] map_value_arg440;
  input [9:0] map_value_arg441;
  wire [9:0] map_value_arg441;
  input [9:0] map_value_arg442;
  wire [9:0] map_value_arg442;
  input [9:0] map_value_arg443;
  wire [9:0] map_value_arg443;
  input [9:0] map_value_arg444;
  wire [9:0] map_value_arg444;
  input [9:0] map_value_arg445;
  wire [9:0] map_value_arg445;
  input [9:0] map_value_arg446;
  wire [9:0] map_value_arg446;
  input [9:0] map_value_arg447;
  wire [9:0] map_value_arg447;
  input [9:0] map_value_arg448;
  wire [9:0] map_value_arg448;
  input [9:0] map_value_arg449;
  wire [9:0] map_value_arg449;
  input [9:0] map_value_arg450;
  wire [9:0] map_value_arg450;
  input [9:0] map_value_arg451;
  wire [9:0] map_value_arg451;
  input [9:0] map_value_arg452;
  wire [9:0] map_value_arg452;
  input [9:0] map_value_arg453;
  wire [9:0] map_value_arg453;
  input [9:0] map_value_arg454;
  wire [9:0] map_value_arg454;
  input [9:0] map_value_arg455;
  wire [9:0] map_value_arg455;
  input [9:0] map_value_arg456;
  wire [9:0] map_value_arg456;
  input [9:0] map_value_arg457;
  wire [9:0] map_value_arg457;
  input [9:0] map_value_arg458;
  wire [9:0] map_value_arg458;
  input [9:0] map_value_arg459;
  wire [9:0] map_value_arg459;
  input [9:0] map_value_arg460;
  wire [9:0] map_value_arg460;
  input [9:0] map_value_arg461;
  wire [9:0] map_value_arg461;
  input [9:0] map_value_arg462;
  wire [9:0] map_value_arg462;
  input [9:0] map_value_arg463;
  wire [9:0] map_value_arg463;
  input [9:0] map_value_arg464;
  wire [9:0] map_value_arg464;
  input [9:0] map_value_arg465;
  wire [9:0] map_value_arg465;
  input [9:0] map_value_arg466;
  wire [9:0] map_value_arg466;
  input [9:0] map_value_arg467;
  wire [9:0] map_value_arg467;
  input [9:0] map_value_arg468;
  wire [9:0] map_value_arg468;
  input [9:0] map_value_arg469;
  wire [9:0] map_value_arg469;
  input [9:0] map_value_arg470;
  wire [9:0] map_value_arg470;
  input [9:0] map_value_arg471;
  wire [9:0] map_value_arg471;
  input [9:0] map_value_arg472;
  wire [9:0] map_value_arg472;
  input [9:0] map_value_arg473;
  wire [9:0] map_value_arg473;
  input [9:0] map_value_arg474;
  wire [9:0] map_value_arg474;
  input [9:0] map_value_arg475;
  wire [9:0] map_value_arg475;
  input [9:0] map_value_arg476;
  wire [9:0] map_value_arg476;
  input [9:0] map_value_arg477;
  wire [9:0] map_value_arg477;
  input [9:0] map_value_arg478;
  wire [9:0] map_value_arg478;
  input [9:0] map_value_arg479;
  wire [9:0] map_value_arg479;
  input [9:0] map_value_arg480;
  wire [9:0] map_value_arg480;
  input [9:0] map_value_arg481;
  wire [9:0] map_value_arg481;
  input [9:0] map_value_arg482;
  wire [9:0] map_value_arg482;
  input [9:0] map_value_arg483;
  wire [9:0] map_value_arg483;
  input [9:0] map_value_arg484;
  wire [9:0] map_value_arg484;
  input [9:0] map_value_arg485;
  wire [9:0] map_value_arg485;
  input [9:0] map_value_arg486;
  wire [9:0] map_value_arg486;
  input [9:0] map_value_arg487;
  wire [9:0] map_value_arg487;
  input [9:0] map_value_arg488;
  wire [9:0] map_value_arg488;
  input [9:0] map_value_arg489;
  wire [9:0] map_value_arg489;
  input [9:0] map_value_arg490;
  wire [9:0] map_value_arg490;
  input [9:0] map_value_arg491;
  wire [9:0] map_value_arg491;
  input [9:0] map_value_arg492;
  wire [9:0] map_value_arg492;
  input [9:0] map_value_arg493;
  wire [9:0] map_value_arg493;
  input [9:0] map_value_arg494;
  wire [9:0] map_value_arg494;
  input [9:0] map_value_arg495;
  wire [9:0] map_value_arg495;
  input [9:0] map_value_arg496;
  wire [9:0] map_value_arg496;
  input [9:0] map_value_arg497;
  wire [9:0] map_value_arg497;
  input [9:0] map_value_arg498;
  wire [9:0] map_value_arg498;
  input [9:0] map_value_arg499;
  wire [9:0] map_value_arg499;
  input [9:0] map_value_arg500;
  wire [9:0] map_value_arg500;
  input [9:0] map_value_arg501;
  wire [9:0] map_value_arg501;
  input [9:0] map_value_arg502;
  wire [9:0] map_value_arg502;
  input [9:0] map_value_arg503;
  wire [9:0] map_value_arg503;
  input [9:0] map_value_arg504;
  wire [9:0] map_value_arg504;
  input [9:0] map_value_arg505;
  wire [9:0] map_value_arg505;
  input [9:0] map_value_arg506;
  wire [9:0] map_value_arg506;
  input [9:0] map_value_arg507;
  wire [9:0] map_value_arg507;
  input [9:0] map_value_arg508;
  wire [9:0] map_value_arg508;
  input [9:0] map_value_arg509;
  wire [9:0] map_value_arg509;
  input [9:0] map_value_arg510;
  wire [9:0] map_value_arg510;
  input [9:0] map_value_arg511;
  wire [9:0] map_value_arg511;
  output [9:0] kekka_out0;
  wire [9:0] kekka_out0;
  output [9:0] kekka_out1;
  wire [9:0] kekka_out1;
  output [9:0] kekka_out2;
  wire [9:0] kekka_out2;
  output [9:0] kekka_out3;
  wire [9:0] kekka_out3;
  output [9:0] kekka_out4;
  wire [9:0] kekka_out4;
  output [9:0] kekka_out5;
  wire [9:0] kekka_out5;
  output [9:0] kekka_out6;
  wire [9:0] kekka_out6;
  output [9:0] kekka_out7;
  wire [9:0] kekka_out7;
  output [9:0] kekka_out8;
  wire [9:0] kekka_out8;
  output [9:0] kekka_out9;
  wire [9:0] kekka_out9;
  output [9:0] kekka_out10;
  wire [9:0] kekka_out10;
  output [9:0] kekka_out11;
  wire [9:0] kekka_out11;
  output [9:0] kekka_out12;
  wire [9:0] kekka_out12;
  output [9:0] kekka_out13;
  wire [9:0] kekka_out13;
  output [9:0] kekka_out14;
  wire [9:0] kekka_out14;
  output [9:0] kekka_out15;
  wire [9:0] kekka_out15;
  output [9:0] kekka_out16;
  wire [9:0] kekka_out16;
  output [9:0] kekka_out17;
  wire [9:0] kekka_out17;
  output [9:0] kekka_out18;
  wire [9:0] kekka_out18;
  output [9:0] kekka_out19;
  wire [9:0] kekka_out19;
  output [9:0] kekka_out20;
  wire [9:0] kekka_out20;
  output [9:0] kekka_out21;
  wire [9:0] kekka_out21;
  output [9:0] kekka_out22;
  wire [9:0] kekka_out22;
  output [9:0] kekka_out23;
  wire [9:0] kekka_out23;
  output [9:0] kekka_out24;
  wire [9:0] kekka_out24;
  output [9:0] kekka_out25;
  wire [9:0] kekka_out25;
  output [9:0] kekka_out26;
  wire [9:0] kekka_out26;
  output [9:0] kekka_out27;
  wire [9:0] kekka_out27;
  output [9:0] kekka_out28;
  wire [9:0] kekka_out28;
  output [9:0] kekka_out29;
  wire [9:0] kekka_out29;
  output [9:0] kekka_out30;
  wire [9:0] kekka_out30;
  output [9:0] kekka_out31;
  wire [9:0] kekka_out31;
  output [9:0] kekka_out32;
  wire [9:0] kekka_out32;
  output [9:0] kekka_out33;
  wire [9:0] kekka_out33;
  output [9:0] kekka_out34;
  wire [9:0] kekka_out34;
  output [9:0] kekka_out35;
  wire [9:0] kekka_out35;
  output [9:0] kekka_out36;
  wire [9:0] kekka_out36;
  output [9:0] kekka_out37;
  wire [9:0] kekka_out37;
  output [9:0] kekka_out38;
  wire [9:0] kekka_out38;
  output [9:0] kekka_out39;
  wire [9:0] kekka_out39;
  output [9:0] kekka_out40;
  wire [9:0] kekka_out40;
  output [9:0] kekka_out41;
  wire [9:0] kekka_out41;
  output [9:0] kekka_out42;
  wire [9:0] kekka_out42;
  output [9:0] kekka_out43;
  wire [9:0] kekka_out43;
  output [9:0] kekka_out44;
  wire [9:0] kekka_out44;
  output [9:0] kekka_out45;
  wire [9:0] kekka_out45;
  output [9:0] kekka_out46;
  wire [9:0] kekka_out46;
  output [9:0] kekka_out47;
  wire [9:0] kekka_out47;
  output [9:0] kekka_out48;
  wire [9:0] kekka_out48;
  output [9:0] kekka_out49;
  wire [9:0] kekka_out49;
  output [9:0] kekka_out50;
  wire [9:0] kekka_out50;
  output [9:0] kekka_out51;
  wire [9:0] kekka_out51;
  output [9:0] kekka_out52;
  wire [9:0] kekka_out52;
  output [9:0] kekka_out53;
  wire [9:0] kekka_out53;
  output [9:0] kekka_out54;
  wire [9:0] kekka_out54;
  output [9:0] kekka_out55;
  wire [9:0] kekka_out55;
  output [9:0] kekka_out56;
  wire [9:0] kekka_out56;
  output [9:0] kekka_out57;
  wire [9:0] kekka_out57;
  output [9:0] kekka_out58;
  wire [9:0] kekka_out58;
  output [9:0] kekka_out59;
  wire [9:0] kekka_out59;
  output [9:0] kekka_out60;
  wire [9:0] kekka_out60;
  output [9:0] kekka_out61;
  wire [9:0] kekka_out61;
  output [9:0] kekka_out62;
  wire [9:0] kekka_out62;
  output [9:0] kekka_out63;
  wire [9:0] kekka_out63;
  output [9:0] kekka_out64;
  wire [9:0] kekka_out64;
  output [9:0] kekka_out65;
  wire [9:0] kekka_out65;
  output [9:0] kekka_out66;
  wire [9:0] kekka_out66;
  output [9:0] kekka_out67;
  wire [9:0] kekka_out67;
  output [9:0] kekka_out68;
  wire [9:0] kekka_out68;
  output [9:0] kekka_out69;
  wire [9:0] kekka_out69;
  output [9:0] kekka_out70;
  wire [9:0] kekka_out70;
  output [9:0] kekka_out71;
  wire [9:0] kekka_out71;
  output [9:0] kekka_out72;
  wire [9:0] kekka_out72;
  output [9:0] kekka_out73;
  wire [9:0] kekka_out73;
  output [9:0] kekka_out74;
  wire [9:0] kekka_out74;
  output [9:0] kekka_out75;
  wire [9:0] kekka_out75;
  output [9:0] kekka_out76;
  wire [9:0] kekka_out76;
  output [9:0] kekka_out77;
  wire [9:0] kekka_out77;
  output [9:0] kekka_out78;
  wire [9:0] kekka_out78;
  output [9:0] kekka_out79;
  wire [9:0] kekka_out79;
  output [9:0] kekka_out80;
  wire [9:0] kekka_out80;
  output [9:0] kekka_out81;
  wire [9:0] kekka_out81;
  output [9:0] kekka_out82;
  wire [9:0] kekka_out82;
  output [9:0] kekka_out83;
  wire [9:0] kekka_out83;
  output [9:0] kekka_out84;
  wire [9:0] kekka_out84;
  output [9:0] kekka_out85;
  wire [9:0] kekka_out85;
  output [9:0] kekka_out86;
  wire [9:0] kekka_out86;
  output [9:0] kekka_out87;
  wire [9:0] kekka_out87;
  output [9:0] kekka_out88;
  wire [9:0] kekka_out88;
  output [9:0] kekka_out89;
  wire [9:0] kekka_out89;
  output [9:0] kekka_out90;
  wire [9:0] kekka_out90;
  output [9:0] kekka_out91;
  wire [9:0] kekka_out91;
  output [9:0] kekka_out92;
  wire [9:0] kekka_out92;
  output [9:0] kekka_out93;
  wire [9:0] kekka_out93;
  output [9:0] kekka_out94;
  wire [9:0] kekka_out94;
  output [9:0] kekka_out95;
  wire [9:0] kekka_out95;
  output [9:0] kekka_out96;
  wire [9:0] kekka_out96;
  output [9:0] kekka_out97;
  wire [9:0] kekka_out97;
  output [9:0] kekka_out98;
  wire [9:0] kekka_out98;
  output [9:0] kekka_out99;
  wire [9:0] kekka_out99;
  output [9:0] kekka_out100;
  wire [9:0] kekka_out100;
  output [9:0] kekka_out101;
  wire [9:0] kekka_out101;
  output [9:0] kekka_out102;
  wire [9:0] kekka_out102;
  output [9:0] kekka_out103;
  wire [9:0] kekka_out103;
  output [9:0] kekka_out104;
  wire [9:0] kekka_out104;
  output [9:0] kekka_out105;
  wire [9:0] kekka_out105;
  output [9:0] kekka_out106;
  wire [9:0] kekka_out106;
  output [9:0] kekka_out107;
  wire [9:0] kekka_out107;
  output [9:0] kekka_out108;
  wire [9:0] kekka_out108;
  output [9:0] kekka_out109;
  wire [9:0] kekka_out109;
  output [9:0] kekka_out110;
  wire [9:0] kekka_out110;
  output [9:0] kekka_out111;
  wire [9:0] kekka_out111;
  output [9:0] kekka_out112;
  wire [9:0] kekka_out112;
  output [9:0] kekka_out113;
  wire [9:0] kekka_out113;
  output [9:0] kekka_out114;
  wire [9:0] kekka_out114;
  output [9:0] kekka_out115;
  wire [9:0] kekka_out115;
  output [9:0] kekka_out116;
  wire [9:0] kekka_out116;
  output [9:0] kekka_out117;
  wire [9:0] kekka_out117;
  output [9:0] kekka_out118;
  wire [9:0] kekka_out118;
  output [9:0] kekka_out119;
  wire [9:0] kekka_out119;
  output [9:0] kekka_out120;
  wire [9:0] kekka_out120;
  output [9:0] kekka_out121;
  wire [9:0] kekka_out121;
  output [9:0] kekka_out122;
  wire [9:0] kekka_out122;
  output [9:0] kekka_out123;
  wire [9:0] kekka_out123;
  output [9:0] kekka_out124;
  wire [9:0] kekka_out124;
  output [9:0] kekka_out125;
  wire [9:0] kekka_out125;
  output [9:0] kekka_out126;
  wire [9:0] kekka_out126;
  output [9:0] kekka_out127;
  wire [9:0] kekka_out127;
  output [9:0] kekka_out128;
  wire [9:0] kekka_out128;
  output [9:0] kekka_out129;
  wire [9:0] kekka_out129;
  output [9:0] kekka_out130;
  wire [9:0] kekka_out130;
  output [9:0] kekka_out131;
  wire [9:0] kekka_out131;
  output [9:0] kekka_out132;
  wire [9:0] kekka_out132;
  output [9:0] kekka_out133;
  wire [9:0] kekka_out133;
  output [9:0] kekka_out134;
  wire [9:0] kekka_out134;
  output [9:0] kekka_out135;
  wire [9:0] kekka_out135;
  output [9:0] kekka_out136;
  wire [9:0] kekka_out136;
  output [9:0] kekka_out137;
  wire [9:0] kekka_out137;
  output [9:0] kekka_out138;
  wire [9:0] kekka_out138;
  output [9:0] kekka_out139;
  wire [9:0] kekka_out139;
  output [9:0] kekka_out140;
  wire [9:0] kekka_out140;
  output [9:0] kekka_out141;
  wire [9:0] kekka_out141;
  output [9:0] kekka_out142;
  wire [9:0] kekka_out142;
  output [9:0] kekka_out143;
  wire [9:0] kekka_out143;
  output [9:0] kekka_out144;
  wire [9:0] kekka_out144;
  output [9:0] kekka_out145;
  wire [9:0] kekka_out145;
  output [9:0] kekka_out146;
  wire [9:0] kekka_out146;
  output [9:0] kekka_out147;
  wire [9:0] kekka_out147;
  output [9:0] kekka_out148;
  wire [9:0] kekka_out148;
  output [9:0] kekka_out149;
  wire [9:0] kekka_out149;
  output [9:0] kekka_out150;
  wire [9:0] kekka_out150;
  output [9:0] kekka_out151;
  wire [9:0] kekka_out151;
  output [9:0] kekka_out152;
  wire [9:0] kekka_out152;
  output [9:0] kekka_out153;
  wire [9:0] kekka_out153;
  output [9:0] kekka_out154;
  wire [9:0] kekka_out154;
  output [9:0] kekka_out155;
  wire [9:0] kekka_out155;
  output [9:0] kekka_out156;
  wire [9:0] kekka_out156;
  output [9:0] kekka_out157;
  wire [9:0] kekka_out157;
  output [9:0] kekka_out158;
  wire [9:0] kekka_out158;
  output [9:0] kekka_out159;
  wire [9:0] kekka_out159;
  output [9:0] kekka_out160;
  wire [9:0] kekka_out160;
  output [9:0] kekka_out161;
  wire [9:0] kekka_out161;
  output [9:0] kekka_out162;
  wire [9:0] kekka_out162;
  output [9:0] kekka_out163;
  wire [9:0] kekka_out163;
  output [9:0] kekka_out164;
  wire [9:0] kekka_out164;
  output [9:0] kekka_out165;
  wire [9:0] kekka_out165;
  output [9:0] kekka_out166;
  wire [9:0] kekka_out166;
  output [9:0] kekka_out167;
  wire [9:0] kekka_out167;
  output [9:0] kekka_out168;
  wire [9:0] kekka_out168;
  output [9:0] kekka_out169;
  wire [9:0] kekka_out169;
  output [9:0] kekka_out170;
  wire [9:0] kekka_out170;
  output [9:0] kekka_out171;
  wire [9:0] kekka_out171;
  output [9:0] kekka_out172;
  wire [9:0] kekka_out172;
  output [9:0] kekka_out173;
  wire [9:0] kekka_out173;
  output [9:0] kekka_out174;
  wire [9:0] kekka_out174;
  output [9:0] kekka_out175;
  wire [9:0] kekka_out175;
  output [9:0] kekka_out176;
  wire [9:0] kekka_out176;
  output [9:0] kekka_out177;
  wire [9:0] kekka_out177;
  output [9:0] kekka_out178;
  wire [9:0] kekka_out178;
  output [9:0] kekka_out179;
  wire [9:0] kekka_out179;
  output [9:0] kekka_out180;
  wire [9:0] kekka_out180;
  output [9:0] kekka_out181;
  wire [9:0] kekka_out181;
  output [9:0] kekka_out182;
  wire [9:0] kekka_out182;
  output [9:0] kekka_out183;
  wire [9:0] kekka_out183;
  output [9:0] kekka_out184;
  wire [9:0] kekka_out184;
  output [9:0] kekka_out185;
  wire [9:0] kekka_out185;
  output [9:0] kekka_out186;
  wire [9:0] kekka_out186;
  output [9:0] kekka_out187;
  wire [9:0] kekka_out187;
  output [9:0] kekka_out188;
  wire [9:0] kekka_out188;
  output [9:0] kekka_out189;
  wire [9:0] kekka_out189;
  output [9:0] kekka_out190;
  wire [9:0] kekka_out190;
  output [9:0] kekka_out191;
  wire [9:0] kekka_out191;
  output [9:0] kekka_out192;
  wire [9:0] kekka_out192;
  output [9:0] kekka_out193;
  wire [9:0] kekka_out193;
  output [9:0] kekka_out194;
  wire [9:0] kekka_out194;
  output [9:0] kekka_out195;
  wire [9:0] kekka_out195;
  output [9:0] kekka_out196;
  wire [9:0] kekka_out196;
  output [9:0] kekka_out197;
  wire [9:0] kekka_out197;
  output [9:0] kekka_out198;
  wire [9:0] kekka_out198;
  output [9:0] kekka_out199;
  wire [9:0] kekka_out199;
  output [9:0] kekka_out200;
  wire [9:0] kekka_out200;
  output [9:0] kekka_out201;
  wire [9:0] kekka_out201;
  output [9:0] kekka_out202;
  wire [9:0] kekka_out202;
  output [9:0] kekka_out203;
  wire [9:0] kekka_out203;
  output [9:0] kekka_out204;
  wire [9:0] kekka_out204;
  output [9:0] kekka_out205;
  wire [9:0] kekka_out205;
  output [9:0] kekka_out206;
  wire [9:0] kekka_out206;
  output [9:0] kekka_out207;
  wire [9:0] kekka_out207;
  output [9:0] kekka_out208;
  wire [9:0] kekka_out208;
  output [9:0] kekka_out209;
  wire [9:0] kekka_out209;
  output [9:0] kekka_out210;
  wire [9:0] kekka_out210;
  output [9:0] kekka_out211;
  wire [9:0] kekka_out211;
  output [9:0] kekka_out212;
  wire [9:0] kekka_out212;
  output [9:0] kekka_out213;
  wire [9:0] kekka_out213;
  output [9:0] kekka_out214;
  wire [9:0] kekka_out214;
  output [9:0] kekka_out215;
  wire [9:0] kekka_out215;
  output [9:0] kekka_out216;
  wire [9:0] kekka_out216;
  output [9:0] kekka_out217;
  wire [9:0] kekka_out217;
  output [9:0] kekka_out218;
  wire [9:0] kekka_out218;
  output [9:0] kekka_out219;
  wire [9:0] kekka_out219;
  output [9:0] kekka_out220;
  wire [9:0] kekka_out220;
  output [9:0] kekka_out221;
  wire [9:0] kekka_out221;
  output [9:0] kekka_out222;
  wire [9:0] kekka_out222;
  input in_do;
  wire in_do;
  output end_meiro;
  wire end_meiro;
  reg [9:0] count;
  wire [9:0] move_out;
  wire [9:0] _seachx_data_in33;
  wire [9:0] _seachx_data_in34;
  wire [9:0] _seachx_data_in35;
  wire [9:0] _seachx_data_in36;
  wire [9:0] _seachx_data_in37;
  wire [9:0] _seachx_data_in38;
  wire [9:0] _seachx_data_in39;
  wire [9:0] _seachx_data_in40;
  wire [9:0] _seachx_data_in41;
  wire [9:0] _seachx_data_in42;
  wire [9:0] _seachx_data_in43;
  wire [9:0] _seachx_data_in44;
  wire [9:0] _seachx_data_in45;
  wire [9:0] _seachx_data_in46;
  wire [9:0] _seachx_data_in47;
  wire [9:0] _seachx_data_in48;
  wire [9:0] _seachx_data_in49;
  wire [9:0] _seachx_data_in50;
  wire [9:0] _seachx_data_in51;
  wire [9:0] _seachx_data_in52;
  wire [9:0] _seachx_data_in53;
  wire [9:0] _seachx_data_in54;
  wire [9:0] _seachx_data_in55;
  wire [9:0] _seachx_data_in56;
  wire [9:0] _seachx_data_in57;
  wire [9:0] _seachx_data_in58;
  wire [9:0] _seachx_data_in59;
  wire [9:0] _seachx_data_in60;
  wire [9:0] _seachx_data_in61;
  wire [9:0] _seachx_data_in62;
  wire [9:0] _seachx_data_in65;
  wire [9:0] _seachx_data_in66;
  wire [9:0] _seachx_data_in67;
  wire [9:0] _seachx_data_in68;
  wire [9:0] _seachx_data_in69;
  wire [9:0] _seachx_data_in70;
  wire [9:0] _seachx_data_in71;
  wire [9:0] _seachx_data_in72;
  wire [9:0] _seachx_data_in73;
  wire [9:0] _seachx_data_in74;
  wire [9:0] _seachx_data_in75;
  wire [9:0] _seachx_data_in76;
  wire [9:0] _seachx_data_in77;
  wire [9:0] _seachx_data_in78;
  wire [9:0] _seachx_data_in79;
  wire [9:0] _seachx_data_in80;
  wire [9:0] _seachx_data_in81;
  wire [9:0] _seachx_data_in82;
  wire [9:0] _seachx_data_in83;
  wire [9:0] _seachx_data_in84;
  wire [9:0] _seachx_data_in85;
  wire [9:0] _seachx_data_in86;
  wire [9:0] _seachx_data_in87;
  wire [9:0] _seachx_data_in88;
  wire [9:0] _seachx_data_in89;
  wire [9:0] _seachx_data_in90;
  wire [9:0] _seachx_data_in91;
  wire [9:0] _seachx_data_in92;
  wire [9:0] _seachx_data_in93;
  wire [9:0] _seachx_data_in94;
  wire [9:0] _seachx_data_in97;
  wire [9:0] _seachx_data_in98;
  wire [9:0] _seachx_data_in99;
  wire [9:0] _seachx_data_in100;
  wire [9:0] _seachx_data_in101;
  wire [9:0] _seachx_data_in102;
  wire [9:0] _seachx_data_in103;
  wire [9:0] _seachx_data_in104;
  wire [9:0] _seachx_data_in105;
  wire [9:0] _seachx_data_in106;
  wire [9:0] _seachx_data_in107;
  wire [9:0] _seachx_data_in108;
  wire [9:0] _seachx_data_in109;
  wire [9:0] _seachx_data_in110;
  wire [9:0] _seachx_data_in111;
  wire [9:0] _seachx_data_in112;
  wire [9:0] _seachx_data_in113;
  wire [9:0] _seachx_data_in114;
  wire [9:0] _seachx_data_in115;
  wire [9:0] _seachx_data_in116;
  wire [9:0] _seachx_data_in117;
  wire [9:0] _seachx_data_in118;
  wire [9:0] _seachx_data_in119;
  wire [9:0] _seachx_data_in120;
  wire [9:0] _seachx_data_in121;
  wire [9:0] _seachx_data_in122;
  wire [9:0] _seachx_data_in123;
  wire [9:0] _seachx_data_in124;
  wire [9:0] _seachx_data_in125;
  wire [9:0] _seachx_data_in126;
  wire [9:0] _seachx_data_in129;
  wire [9:0] _seachx_data_in130;
  wire [9:0] _seachx_data_in131;
  wire [9:0] _seachx_data_in132;
  wire [9:0] _seachx_data_in133;
  wire [9:0] _seachx_data_in134;
  wire [9:0] _seachx_data_in135;
  wire [9:0] _seachx_data_in136;
  wire [9:0] _seachx_data_in137;
  wire [9:0] _seachx_data_in138;
  wire [9:0] _seachx_data_in139;
  wire [9:0] _seachx_data_in140;
  wire [9:0] _seachx_data_in141;
  wire [9:0] _seachx_data_in142;
  wire [9:0] _seachx_data_in143;
  wire [9:0] _seachx_data_in144;
  wire [9:0] _seachx_data_in145;
  wire [9:0] _seachx_data_in146;
  wire [9:0] _seachx_data_in147;
  wire [9:0] _seachx_data_in148;
  wire [9:0] _seachx_data_in149;
  wire [9:0] _seachx_data_in150;
  wire [9:0] _seachx_data_in151;
  wire [9:0] _seachx_data_in152;
  wire [9:0] _seachx_data_in153;
  wire [9:0] _seachx_data_in154;
  wire [9:0] _seachx_data_in155;
  wire [9:0] _seachx_data_in156;
  wire [9:0] _seachx_data_in157;
  wire [9:0] _seachx_data_in158;
  wire [9:0] _seachx_data_in161;
  wire [9:0] _seachx_data_in162;
  wire [9:0] _seachx_data_in163;
  wire [9:0] _seachx_data_in164;
  wire [9:0] _seachx_data_in165;
  wire [9:0] _seachx_data_in166;
  wire [9:0] _seachx_data_in167;
  wire [9:0] _seachx_data_in168;
  wire [9:0] _seachx_data_in169;
  wire [9:0] _seachx_data_in170;
  wire [9:0] _seachx_data_in171;
  wire [9:0] _seachx_data_in172;
  wire [9:0] _seachx_data_in173;
  wire [9:0] _seachx_data_in174;
  wire [9:0] _seachx_data_in175;
  wire [9:0] _seachx_data_in176;
  wire [9:0] _seachx_data_in177;
  wire [9:0] _seachx_data_in178;
  wire [9:0] _seachx_data_in179;
  wire [9:0] _seachx_data_in180;
  wire [9:0] _seachx_data_in181;
  wire [9:0] _seachx_data_in182;
  wire [9:0] _seachx_data_in183;
  wire [9:0] _seachx_data_in184;
  wire [9:0] _seachx_data_in185;
  wire [9:0] _seachx_data_in186;
  wire [9:0] _seachx_data_in187;
  wire [9:0] _seachx_data_in188;
  wire [9:0] _seachx_data_in189;
  wire [9:0] _seachx_data_in190;
  wire [9:0] _seachx_data_in193;
  wire [9:0] _seachx_data_in194;
  wire [9:0] _seachx_data_in195;
  wire [9:0] _seachx_data_in196;
  wire [9:0] _seachx_data_in197;
  wire [9:0] _seachx_data_in198;
  wire [9:0] _seachx_data_in199;
  wire [9:0] _seachx_data_in200;
  wire [9:0] _seachx_data_in201;
  wire [9:0] _seachx_data_in202;
  wire [9:0] _seachx_data_in203;
  wire [9:0] _seachx_data_in204;
  wire [9:0] _seachx_data_in205;
  wire [9:0] _seachx_data_in206;
  wire [9:0] _seachx_data_in207;
  wire [9:0] _seachx_data_in208;
  wire [9:0] _seachx_data_in209;
  wire [9:0] _seachx_data_in210;
  wire [9:0] _seachx_data_in211;
  wire [9:0] _seachx_data_in212;
  wire [9:0] _seachx_data_in213;
  wire [9:0] _seachx_data_in214;
  wire [9:0] _seachx_data_in215;
  wire [9:0] _seachx_data_in216;
  wire [9:0] _seachx_data_in217;
  wire [9:0] _seachx_data_in218;
  wire [9:0] _seachx_data_in219;
  wire [9:0] _seachx_data_in220;
  wire [9:0] _seachx_data_in221;
  wire [9:0] _seachx_data_in222;
  wire [9:0] _seachx_data_in225;
  wire [9:0] _seachx_data_in226;
  wire [9:0] _seachx_data_in227;
  wire [9:0] _seachx_data_in228;
  wire [9:0] _seachx_data_in229;
  wire [9:0] _seachx_data_in230;
  wire [9:0] _seachx_data_in231;
  wire [9:0] _seachx_data_in232;
  wire [9:0] _seachx_data_in233;
  wire [9:0] _seachx_data_in234;
  wire [9:0] _seachx_data_in235;
  wire [9:0] _seachx_data_in236;
  wire [9:0] _seachx_data_in237;
  wire [9:0] _seachx_data_in238;
  wire [9:0] _seachx_data_in239;
  wire [9:0] _seachx_data_in240;
  wire [9:0] _seachx_data_in241;
  wire [9:0] _seachx_data_in242;
  wire [9:0] _seachx_data_in243;
  wire [9:0] _seachx_data_in244;
  wire [9:0] _seachx_data_in245;
  wire [9:0] _seachx_data_in246;
  wire [9:0] _seachx_data_in247;
  wire [9:0] _seachx_data_in248;
  wire [9:0] _seachx_data_in249;
  wire [9:0] _seachx_data_in250;
  wire [9:0] _seachx_data_in251;
  wire [9:0] _seachx_data_in252;
  wire [9:0] _seachx_data_in253;
  wire [9:0] _seachx_data_in254;
  wire [9:0] _seachx_data_in257;
  wire [9:0] _seachx_data_in258;
  wire [9:0] _seachx_data_in259;
  wire [9:0] _seachx_data_in260;
  wire [9:0] _seachx_data_in261;
  wire [9:0] _seachx_data_in262;
  wire [9:0] _seachx_data_in263;
  wire [9:0] _seachx_data_in264;
  wire [9:0] _seachx_data_in265;
  wire [9:0] _seachx_data_in266;
  wire [9:0] _seachx_data_in267;
  wire [9:0] _seachx_data_in268;
  wire [9:0] _seachx_data_in269;
  wire [9:0] _seachx_data_in270;
  wire [9:0] _seachx_data_in271;
  wire [9:0] _seachx_data_in272;
  wire [9:0] _seachx_data_in273;
  wire [9:0] _seachx_data_in274;
  wire [9:0] _seachx_data_in275;
  wire [9:0] _seachx_data_in276;
  wire [9:0] _seachx_data_in277;
  wire [9:0] _seachx_data_in278;
  wire [9:0] _seachx_data_in279;
  wire [9:0] _seachx_data_in280;
  wire [9:0] _seachx_data_in281;
  wire [9:0] _seachx_data_in282;
  wire [9:0] _seachx_data_in283;
  wire [9:0] _seachx_data_in284;
  wire [9:0] _seachx_data_in285;
  wire [9:0] _seachx_data_in286;
  wire [9:0] _seachx_data_in289;
  wire [9:0] _seachx_data_in290;
  wire [9:0] _seachx_data_in291;
  wire [9:0] _seachx_data_in292;
  wire [9:0] _seachx_data_in293;
  wire [9:0] _seachx_data_in294;
  wire [9:0] _seachx_data_in295;
  wire [9:0] _seachx_data_in296;
  wire [9:0] _seachx_data_in297;
  wire [9:0] _seachx_data_in298;
  wire [9:0] _seachx_data_in299;
  wire [9:0] _seachx_data_in300;
  wire [9:0] _seachx_data_in301;
  wire [9:0] _seachx_data_in302;
  wire [9:0] _seachx_data_in303;
  wire [9:0] _seachx_data_in304;
  wire [9:0] _seachx_data_in305;
  wire [9:0] _seachx_data_in306;
  wire [9:0] _seachx_data_in307;
  wire [9:0] _seachx_data_in308;
  wire [9:0] _seachx_data_in309;
  wire [9:0] _seachx_data_in310;
  wire [9:0] _seachx_data_in311;
  wire [9:0] _seachx_data_in312;
  wire [9:0] _seachx_data_in313;
  wire [9:0] _seachx_data_in314;
  wire [9:0] _seachx_data_in315;
  wire [9:0] _seachx_data_in316;
  wire [9:0] _seachx_data_in317;
  wire [9:0] _seachx_data_in318;
  wire [9:0] _seachx_data_in321;
  wire [9:0] _seachx_data_in322;
  wire [9:0] _seachx_data_in323;
  wire [9:0] _seachx_data_in324;
  wire [9:0] _seachx_data_in325;
  wire [9:0] _seachx_data_in326;
  wire [9:0] _seachx_data_in327;
  wire [9:0] _seachx_data_in328;
  wire [9:0] _seachx_data_in329;
  wire [9:0] _seachx_data_in330;
  wire [9:0] _seachx_data_in331;
  wire [9:0] _seachx_data_in332;
  wire [9:0] _seachx_data_in333;
  wire [9:0] _seachx_data_in334;
  wire [9:0] _seachx_data_in335;
  wire [9:0] _seachx_data_in336;
  wire [9:0] _seachx_data_in337;
  wire [9:0] _seachx_data_in338;
  wire [9:0] _seachx_data_in339;
  wire [9:0] _seachx_data_in340;
  wire [9:0] _seachx_data_in341;
  wire [9:0] _seachx_data_in342;
  wire [9:0] _seachx_data_in343;
  wire [9:0] _seachx_data_in344;
  wire [9:0] _seachx_data_in345;
  wire [9:0] _seachx_data_in346;
  wire [9:0] _seachx_data_in347;
  wire [9:0] _seachx_data_in348;
  wire [9:0] _seachx_data_in349;
  wire [9:0] _seachx_data_in350;
  wire [9:0] _seachx_data_in353;
  wire [9:0] _seachx_data_in354;
  wire [9:0] _seachx_data_in355;
  wire [9:0] _seachx_data_in356;
  wire [9:0] _seachx_data_in357;
  wire [9:0] _seachx_data_in358;
  wire [9:0] _seachx_data_in359;
  wire [9:0] _seachx_data_in360;
  wire [9:0] _seachx_data_in361;
  wire [9:0] _seachx_data_in362;
  wire [9:0] _seachx_data_in363;
  wire [9:0] _seachx_data_in364;
  wire [9:0] _seachx_data_in365;
  wire [9:0] _seachx_data_in366;
  wire [9:0] _seachx_data_in367;
  wire [9:0] _seachx_data_in368;
  wire [9:0] _seachx_data_in369;
  wire [9:0] _seachx_data_in370;
  wire [9:0] _seachx_data_in371;
  wire [9:0] _seachx_data_in372;
  wire [9:0] _seachx_data_in373;
  wire [9:0] _seachx_data_in374;
  wire [9:0] _seachx_data_in375;
  wire [9:0] _seachx_data_in376;
  wire [9:0] _seachx_data_in377;
  wire [9:0] _seachx_data_in378;
  wire [9:0] _seachx_data_in379;
  wire [9:0] _seachx_data_in380;
  wire [9:0] _seachx_data_in381;
  wire [9:0] _seachx_data_in382;
  wire [9:0] _seachx_data_in385;
  wire [9:0] _seachx_data_in386;
  wire [9:0] _seachx_data_in387;
  wire [9:0] _seachx_data_in388;
  wire [9:0] _seachx_data_in389;
  wire [9:0] _seachx_data_in390;
  wire [9:0] _seachx_data_in391;
  wire [9:0] _seachx_data_in392;
  wire [9:0] _seachx_data_in393;
  wire [9:0] _seachx_data_in394;
  wire [9:0] _seachx_data_in395;
  wire [9:0] _seachx_data_in396;
  wire [9:0] _seachx_data_in397;
  wire [9:0] _seachx_data_in398;
  wire [9:0] _seachx_data_in399;
  wire [9:0] _seachx_data_in400;
  wire [9:0] _seachx_data_in401;
  wire [9:0] _seachx_data_in402;
  wire [9:0] _seachx_data_in403;
  wire [9:0] _seachx_data_in404;
  wire [9:0] _seachx_data_in405;
  wire [9:0] _seachx_data_in406;
  wire [9:0] _seachx_data_in407;
  wire [9:0] _seachx_data_in408;
  wire [9:0] _seachx_data_in409;
  wire [9:0] _seachx_data_in410;
  wire [9:0] _seachx_data_in411;
  wire [9:0] _seachx_data_in412;
  wire [9:0] _seachx_data_in413;
  wire [9:0] _seachx_data_in414;
  wire [9:0] _seachx_data_in417;
  wire [9:0] _seachx_data_in418;
  wire [9:0] _seachx_data_in419;
  wire [9:0] _seachx_data_in420;
  wire [9:0] _seachx_data_in421;
  wire [9:0] _seachx_data_in422;
  wire [9:0] _seachx_data_in423;
  wire [9:0] _seachx_data_in424;
  wire [9:0] _seachx_data_in425;
  wire [9:0] _seachx_data_in426;
  wire [9:0] _seachx_data_in427;
  wire [9:0] _seachx_data_in428;
  wire [9:0] _seachx_data_in429;
  wire [9:0] _seachx_data_in430;
  wire [9:0] _seachx_data_in431;
  wire [9:0] _seachx_data_in432;
  wire [9:0] _seachx_data_in433;
  wire [9:0] _seachx_data_in434;
  wire [9:0] _seachx_data_in435;
  wire [9:0] _seachx_data_in436;
  wire [9:0] _seachx_data_in437;
  wire [9:0] _seachx_data_in438;
  wire [9:0] _seachx_data_in439;
  wire [9:0] _seachx_data_in440;
  wire [9:0] _seachx_data_in441;
  wire [9:0] _seachx_data_in442;
  wire [9:0] _seachx_data_in443;
  wire [9:0] _seachx_data_in444;
  wire [9:0] _seachx_data_in445;
  wire [9:0] _seachx_data_in446;
  wire [9:0] _seachx_data_in449;
  wire [9:0] _seachx_data_in450;
  wire [9:0] _seachx_data_in451;
  wire [9:0] _seachx_data_in452;
  wire [9:0] _seachx_data_in453;
  wire [9:0] _seachx_data_in454;
  wire [9:0] _seachx_data_in455;
  wire [9:0] _seachx_data_in456;
  wire [9:0] _seachx_data_in457;
  wire [9:0] _seachx_data_in458;
  wire [9:0] _seachx_data_in459;
  wire [9:0] _seachx_data_in460;
  wire [9:0] _seachx_data_in461;
  wire [9:0] _seachx_data_in462;
  wire [9:0] _seachx_data_in463;
  wire [9:0] _seachx_data_in464;
  wire [9:0] _seachx_data_in465;
  wire [9:0] _seachx_data_in466;
  wire [9:0] _seachx_data_in467;
  wire [9:0] _seachx_data_in468;
  wire [9:0] _seachx_data_in469;
  wire [9:0] _seachx_data_in470;
  wire [9:0] _seachx_data_in471;
  wire [9:0] _seachx_data_in472;
  wire [9:0] _seachx_data_in473;
  wire [9:0] _seachx_data_in474;
  wire [9:0] _seachx_data_in475;
  wire [9:0] _seachx_data_in476;
  wire [9:0] _seachx_data_in477;
  wire [9:0] _seachx_data_in478;
  wire [9:0] _seachx_data_out33;
  wire [9:0] _seachx_data_out34;
  wire [9:0] _seachx_data_out35;
  wire [9:0] _seachx_data_out36;
  wire [9:0] _seachx_data_out37;
  wire [9:0] _seachx_data_out38;
  wire [9:0] _seachx_data_out39;
  wire [9:0] _seachx_data_out40;
  wire [9:0] _seachx_data_out41;
  wire [9:0] _seachx_data_out42;
  wire [9:0] _seachx_data_out43;
  wire [9:0] _seachx_data_out44;
  wire [9:0] _seachx_data_out45;
  wire [9:0] _seachx_data_out46;
  wire [9:0] _seachx_data_out47;
  wire [9:0] _seachx_data_out48;
  wire [9:0] _seachx_data_out49;
  wire [9:0] _seachx_data_out50;
  wire [9:0] _seachx_data_out51;
  wire [9:0] _seachx_data_out52;
  wire [9:0] _seachx_data_out53;
  wire [9:0] _seachx_data_out54;
  wire [9:0] _seachx_data_out55;
  wire [9:0] _seachx_data_out56;
  wire [9:0] _seachx_data_out57;
  wire [9:0] _seachx_data_out58;
  wire [9:0] _seachx_data_out59;
  wire [9:0] _seachx_data_out60;
  wire [9:0] _seachx_data_out61;
  wire [9:0] _seachx_data_out62;
  wire [9:0] _seachx_data_out65;
  wire [9:0] _seachx_data_out66;
  wire [9:0] _seachx_data_out67;
  wire [9:0] _seachx_data_out68;
  wire [9:0] _seachx_data_out69;
  wire [9:0] _seachx_data_out70;
  wire [9:0] _seachx_data_out71;
  wire [9:0] _seachx_data_out72;
  wire [9:0] _seachx_data_out73;
  wire [9:0] _seachx_data_out74;
  wire [9:0] _seachx_data_out75;
  wire [9:0] _seachx_data_out76;
  wire [9:0] _seachx_data_out77;
  wire [9:0] _seachx_data_out78;
  wire [9:0] _seachx_data_out79;
  wire [9:0] _seachx_data_out80;
  wire [9:0] _seachx_data_out81;
  wire [9:0] _seachx_data_out82;
  wire [9:0] _seachx_data_out83;
  wire [9:0] _seachx_data_out84;
  wire [9:0] _seachx_data_out85;
  wire [9:0] _seachx_data_out86;
  wire [9:0] _seachx_data_out87;
  wire [9:0] _seachx_data_out88;
  wire [9:0] _seachx_data_out89;
  wire [9:0] _seachx_data_out90;
  wire [9:0] _seachx_data_out91;
  wire [9:0] _seachx_data_out92;
  wire [9:0] _seachx_data_out93;
  wire [9:0] _seachx_data_out94;
  wire [9:0] _seachx_data_out97;
  wire [9:0] _seachx_data_out98;
  wire [9:0] _seachx_data_out99;
  wire [9:0] _seachx_data_out100;
  wire [9:0] _seachx_data_out101;
  wire [9:0] _seachx_data_out102;
  wire [9:0] _seachx_data_out103;
  wire [9:0] _seachx_data_out104;
  wire [9:0] _seachx_data_out105;
  wire [9:0] _seachx_data_out106;
  wire [9:0] _seachx_data_out107;
  wire [9:0] _seachx_data_out108;
  wire [9:0] _seachx_data_out109;
  wire [9:0] _seachx_data_out110;
  wire [9:0] _seachx_data_out111;
  wire [9:0] _seachx_data_out112;
  wire [9:0] _seachx_data_out113;
  wire [9:0] _seachx_data_out114;
  wire [9:0] _seachx_data_out115;
  wire [9:0] _seachx_data_out116;
  wire [9:0] _seachx_data_out117;
  wire [9:0] _seachx_data_out118;
  wire [9:0] _seachx_data_out119;
  wire [9:0] _seachx_data_out120;
  wire [9:0] _seachx_data_out121;
  wire [9:0] _seachx_data_out122;
  wire [9:0] _seachx_data_out123;
  wire [9:0] _seachx_data_out124;
  wire [9:0] _seachx_data_out125;
  wire [9:0] _seachx_data_out126;
  wire [9:0] _seachx_data_out129;
  wire [9:0] _seachx_data_out130;
  wire [9:0] _seachx_data_out131;
  wire [9:0] _seachx_data_out132;
  wire [9:0] _seachx_data_out133;
  wire [9:0] _seachx_data_out134;
  wire [9:0] _seachx_data_out135;
  wire [9:0] _seachx_data_out136;
  wire [9:0] _seachx_data_out137;
  wire [9:0] _seachx_data_out138;
  wire [9:0] _seachx_data_out139;
  wire [9:0] _seachx_data_out140;
  wire [9:0] _seachx_data_out141;
  wire [9:0] _seachx_data_out142;
  wire [9:0] _seachx_data_out143;
  wire [9:0] _seachx_data_out144;
  wire [9:0] _seachx_data_out145;
  wire [9:0] _seachx_data_out146;
  wire [9:0] _seachx_data_out147;
  wire [9:0] _seachx_data_out148;
  wire [9:0] _seachx_data_out149;
  wire [9:0] _seachx_data_out150;
  wire [9:0] _seachx_data_out151;
  wire [9:0] _seachx_data_out152;
  wire [9:0] _seachx_data_out153;
  wire [9:0] _seachx_data_out154;
  wire [9:0] _seachx_data_out155;
  wire [9:0] _seachx_data_out156;
  wire [9:0] _seachx_data_out157;
  wire [9:0] _seachx_data_out158;
  wire [9:0] _seachx_data_out161;
  wire [9:0] _seachx_data_out162;
  wire [9:0] _seachx_data_out163;
  wire [9:0] _seachx_data_out164;
  wire [9:0] _seachx_data_out165;
  wire [9:0] _seachx_data_out166;
  wire [9:0] _seachx_data_out167;
  wire [9:0] _seachx_data_out168;
  wire [9:0] _seachx_data_out169;
  wire [9:0] _seachx_data_out170;
  wire [9:0] _seachx_data_out171;
  wire [9:0] _seachx_data_out172;
  wire [9:0] _seachx_data_out173;
  wire [9:0] _seachx_data_out174;
  wire [9:0] _seachx_data_out175;
  wire [9:0] _seachx_data_out176;
  wire [9:0] _seachx_data_out177;
  wire [9:0] _seachx_data_out178;
  wire [9:0] _seachx_data_out179;
  wire [9:0] _seachx_data_out180;
  wire [9:0] _seachx_data_out181;
  wire [9:0] _seachx_data_out182;
  wire [9:0] _seachx_data_out183;
  wire [9:0] _seachx_data_out184;
  wire [9:0] _seachx_data_out185;
  wire [9:0] _seachx_data_out186;
  wire [9:0] _seachx_data_out187;
  wire [9:0] _seachx_data_out188;
  wire [9:0] _seachx_data_out189;
  wire [9:0] _seachx_data_out190;
  wire [9:0] _seachx_data_out193;
  wire [9:0] _seachx_data_out194;
  wire [9:0] _seachx_data_out195;
  wire [9:0] _seachx_data_out196;
  wire [9:0] _seachx_data_out197;
  wire [9:0] _seachx_data_out198;
  wire [9:0] _seachx_data_out199;
  wire [9:0] _seachx_data_out200;
  wire [9:0] _seachx_data_out201;
  wire [9:0] _seachx_data_out202;
  wire [9:0] _seachx_data_out203;
  wire [9:0] _seachx_data_out204;
  wire [9:0] _seachx_data_out205;
  wire [9:0] _seachx_data_out206;
  wire [9:0] _seachx_data_out207;
  wire [9:0] _seachx_data_out208;
  wire [9:0] _seachx_data_out209;
  wire [9:0] _seachx_data_out210;
  wire [9:0] _seachx_data_out211;
  wire [9:0] _seachx_data_out212;
  wire [9:0] _seachx_data_out213;
  wire [9:0] _seachx_data_out214;
  wire [9:0] _seachx_data_out215;
  wire [9:0] _seachx_data_out216;
  wire [9:0] _seachx_data_out217;
  wire [9:0] _seachx_data_out218;
  wire [9:0] _seachx_data_out219;
  wire [9:0] _seachx_data_out220;
  wire [9:0] _seachx_data_out221;
  wire [9:0] _seachx_data_out222;
  wire [9:0] _seachx_data_out225;
  wire [9:0] _seachx_data_out226;
  wire [9:0] _seachx_data_out227;
  wire [9:0] _seachx_data_out228;
  wire [9:0] _seachx_data_out229;
  wire [9:0] _seachx_data_out230;
  wire [9:0] _seachx_data_out231;
  wire [9:0] _seachx_data_out232;
  wire [9:0] _seachx_data_out233;
  wire [9:0] _seachx_data_out234;
  wire [9:0] _seachx_data_out235;
  wire [9:0] _seachx_data_out236;
  wire [9:0] _seachx_data_out237;
  wire [9:0] _seachx_data_out238;
  wire [9:0] _seachx_data_out239;
  wire [9:0] _seachx_data_out240;
  wire [9:0] _seachx_data_out241;
  wire [9:0] _seachx_data_out242;
  wire [9:0] _seachx_data_out243;
  wire [9:0] _seachx_data_out244;
  wire [9:0] _seachx_data_out245;
  wire [9:0] _seachx_data_out246;
  wire [9:0] _seachx_data_out247;
  wire [9:0] _seachx_data_out248;
  wire [9:0] _seachx_data_out249;
  wire [9:0] _seachx_data_out250;
  wire [9:0] _seachx_data_out251;
  wire [9:0] _seachx_data_out252;
  wire [9:0] _seachx_data_out253;
  wire [9:0] _seachx_data_out254;
  wire [9:0] _seachx_data_out257;
  wire [9:0] _seachx_data_out258;
  wire [9:0] _seachx_data_out259;
  wire [9:0] _seachx_data_out260;
  wire [9:0] _seachx_data_out261;
  wire [9:0] _seachx_data_out262;
  wire [9:0] _seachx_data_out263;
  wire [9:0] _seachx_data_out264;
  wire [9:0] _seachx_data_out265;
  wire [9:0] _seachx_data_out266;
  wire [9:0] _seachx_data_out267;
  wire [9:0] _seachx_data_out268;
  wire [9:0] _seachx_data_out269;
  wire [9:0] _seachx_data_out270;
  wire [9:0] _seachx_data_out271;
  wire [9:0] _seachx_data_out272;
  wire [9:0] _seachx_data_out273;
  wire [9:0] _seachx_data_out274;
  wire [9:0] _seachx_data_out275;
  wire [9:0] _seachx_data_out276;
  wire [9:0] _seachx_data_out277;
  wire [9:0] _seachx_data_out278;
  wire [9:0] _seachx_data_out279;
  wire [9:0] _seachx_data_out280;
  wire [9:0] _seachx_data_out281;
  wire [9:0] _seachx_data_out282;
  wire [9:0] _seachx_data_out283;
  wire [9:0] _seachx_data_out284;
  wire [9:0] _seachx_data_out285;
  wire [9:0] _seachx_data_out286;
  wire [9:0] _seachx_data_out289;
  wire [9:0] _seachx_data_out290;
  wire [9:0] _seachx_data_out291;
  wire [9:0] _seachx_data_out292;
  wire [9:0] _seachx_data_out293;
  wire [9:0] _seachx_data_out294;
  wire [9:0] _seachx_data_out295;
  wire [9:0] _seachx_data_out296;
  wire [9:0] _seachx_data_out297;
  wire [9:0] _seachx_data_out298;
  wire [9:0] _seachx_data_out299;
  wire [9:0] _seachx_data_out300;
  wire [9:0] _seachx_data_out301;
  wire [9:0] _seachx_data_out302;
  wire [9:0] _seachx_data_out303;
  wire [9:0] _seachx_data_out304;
  wire [9:0] _seachx_data_out305;
  wire [9:0] _seachx_data_out306;
  wire [9:0] _seachx_data_out307;
  wire [9:0] _seachx_data_out308;
  wire [9:0] _seachx_data_out309;
  wire [9:0] _seachx_data_out310;
  wire [9:0] _seachx_data_out311;
  wire [9:0] _seachx_data_out312;
  wire [9:0] _seachx_data_out313;
  wire [9:0] _seachx_data_out314;
  wire [9:0] _seachx_data_out315;
  wire [9:0] _seachx_data_out316;
  wire [9:0] _seachx_data_out317;
  wire [9:0] _seachx_data_out318;
  wire [9:0] _seachx_data_out321;
  wire [9:0] _seachx_data_out322;
  wire [9:0] _seachx_data_out323;
  wire [9:0] _seachx_data_out324;
  wire [9:0] _seachx_data_out325;
  wire [9:0] _seachx_data_out326;
  wire [9:0] _seachx_data_out327;
  wire [9:0] _seachx_data_out328;
  wire [9:0] _seachx_data_out329;
  wire [9:0] _seachx_data_out330;
  wire [9:0] _seachx_data_out331;
  wire [9:0] _seachx_data_out332;
  wire [9:0] _seachx_data_out333;
  wire [9:0] _seachx_data_out334;
  wire [9:0] _seachx_data_out335;
  wire [9:0] _seachx_data_out336;
  wire [9:0] _seachx_data_out337;
  wire [9:0] _seachx_data_out338;
  wire [9:0] _seachx_data_out339;
  wire [9:0] _seachx_data_out340;
  wire [9:0] _seachx_data_out341;
  wire [9:0] _seachx_data_out342;
  wire [9:0] _seachx_data_out343;
  wire [9:0] _seachx_data_out344;
  wire [9:0] _seachx_data_out345;
  wire [9:0] _seachx_data_out346;
  wire [9:0] _seachx_data_out347;
  wire [9:0] _seachx_data_out348;
  wire [9:0] _seachx_data_out349;
  wire [9:0] _seachx_data_out350;
  wire [9:0] _seachx_data_out353;
  wire [9:0] _seachx_data_out354;
  wire [9:0] _seachx_data_out355;
  wire [9:0] _seachx_data_out356;
  wire [9:0] _seachx_data_out357;
  wire [9:0] _seachx_data_out358;
  wire [9:0] _seachx_data_out359;
  wire [9:0] _seachx_data_out360;
  wire [9:0] _seachx_data_out361;
  wire [9:0] _seachx_data_out362;
  wire [9:0] _seachx_data_out363;
  wire [9:0] _seachx_data_out364;
  wire [9:0] _seachx_data_out365;
  wire [9:0] _seachx_data_out366;
  wire [9:0] _seachx_data_out367;
  wire [9:0] _seachx_data_out368;
  wire [9:0] _seachx_data_out369;
  wire [9:0] _seachx_data_out370;
  wire [9:0] _seachx_data_out371;
  wire [9:0] _seachx_data_out372;
  wire [9:0] _seachx_data_out373;
  wire [9:0] _seachx_data_out374;
  wire [9:0] _seachx_data_out375;
  wire [9:0] _seachx_data_out376;
  wire [9:0] _seachx_data_out377;
  wire [9:0] _seachx_data_out378;
  wire [9:0] _seachx_data_out379;
  wire [9:0] _seachx_data_out380;
  wire [9:0] _seachx_data_out381;
  wire [9:0] _seachx_data_out382;
  wire [9:0] _seachx_data_out385;
  wire [9:0] _seachx_data_out386;
  wire [9:0] _seachx_data_out387;
  wire [9:0] _seachx_data_out388;
  wire [9:0] _seachx_data_out389;
  wire [9:0] _seachx_data_out390;
  wire [9:0] _seachx_data_out391;
  wire [9:0] _seachx_data_out392;
  wire [9:0] _seachx_data_out393;
  wire [9:0] _seachx_data_out394;
  wire [9:0] _seachx_data_out395;
  wire [9:0] _seachx_data_out396;
  wire [9:0] _seachx_data_out397;
  wire [9:0] _seachx_data_out398;
  wire [9:0] _seachx_data_out399;
  wire [9:0] _seachx_data_out400;
  wire [9:0] _seachx_data_out401;
  wire [9:0] _seachx_data_out402;
  wire [9:0] _seachx_data_out403;
  wire [9:0] _seachx_data_out404;
  wire [9:0] _seachx_data_out405;
  wire [9:0] _seachx_data_out406;
  wire [9:0] _seachx_data_out407;
  wire [9:0] _seachx_data_out408;
  wire [9:0] _seachx_data_out409;
  wire [9:0] _seachx_data_out410;
  wire [9:0] _seachx_data_out411;
  wire [9:0] _seachx_data_out412;
  wire [9:0] _seachx_data_out413;
  wire [9:0] _seachx_data_out414;
  wire [9:0] _seachx_data_out417;
  wire [9:0] _seachx_data_out418;
  wire [9:0] _seachx_data_out419;
  wire [9:0] _seachx_data_out420;
  wire [9:0] _seachx_data_out421;
  wire [9:0] _seachx_data_out422;
  wire [9:0] _seachx_data_out423;
  wire [9:0] _seachx_data_out424;
  wire [9:0] _seachx_data_out425;
  wire [9:0] _seachx_data_out426;
  wire [9:0] _seachx_data_out427;
  wire [9:0] _seachx_data_out428;
  wire [9:0] _seachx_data_out429;
  wire [9:0] _seachx_data_out430;
  wire [9:0] _seachx_data_out431;
  wire [9:0] _seachx_data_out432;
  wire [9:0] _seachx_data_out433;
  wire [9:0] _seachx_data_out434;
  wire [9:0] _seachx_data_out435;
  wire [9:0] _seachx_data_out436;
  wire [9:0] _seachx_data_out437;
  wire [9:0] _seachx_data_out438;
  wire [9:0] _seachx_data_out439;
  wire [9:0] _seachx_data_out440;
  wire [9:0] _seachx_data_out441;
  wire [9:0] _seachx_data_out442;
  wire [9:0] _seachx_data_out443;
  wire [9:0] _seachx_data_out444;
  wire [9:0] _seachx_data_out445;
  wire [9:0] _seachx_data_out446;
  wire [9:0] _seachx_data_out449;
  wire [9:0] _seachx_data_out450;
  wire [9:0] _seachx_data_out451;
  wire [9:0] _seachx_data_out452;
  wire [9:0] _seachx_data_out453;
  wire [9:0] _seachx_data_out454;
  wire [9:0] _seachx_data_out455;
  wire [9:0] _seachx_data_out456;
  wire [9:0] _seachx_data_out457;
  wire [9:0] _seachx_data_out458;
  wire [9:0] _seachx_data_out459;
  wire [9:0] _seachx_data_out460;
  wire [9:0] _seachx_data_out461;
  wire [9:0] _seachx_data_out462;
  wire [9:0] _seachx_data_out463;
  wire [9:0] _seachx_data_out464;
  wire [9:0] _seachx_data_out465;
  wire [9:0] _seachx_data_out466;
  wire [9:0] _seachx_data_out467;
  wire [9:0] _seachx_data_out468;
  wire [9:0] _seachx_data_out469;
  wire [9:0] _seachx_data_out470;
  wire [9:0] _seachx_data_out471;
  wire [9:0] _seachx_data_out472;
  wire [9:0] _seachx_data_out473;
  wire [9:0] _seachx_data_out474;
  wire [9:0] _seachx_data_out475;
  wire [9:0] _seachx_data_out476;
  wire [9:0] _seachx_data_out477;
  wire [9:0] _seachx_data_out478;
  wire [9:0] _seachx_startplot;
  wire [9:0] _seachx_goalplot;
  wire _seachx_in_do;
  wire _seachx_out_do;
  wire _seachx_out_data;
  wire _seachx_p_reset;
  wire _seachx_m_clock;
  wire [9:0] _kanwa_x_data_in33;
  wire [9:0] _kanwa_x_data_in34;
  wire [9:0] _kanwa_x_data_in35;
  wire [9:0] _kanwa_x_data_in36;
  wire [9:0] _kanwa_x_data_in37;
  wire [9:0] _kanwa_x_data_in38;
  wire [9:0] _kanwa_x_data_in39;
  wire [9:0] _kanwa_x_data_in40;
  wire [9:0] _kanwa_x_data_in41;
  wire [9:0] _kanwa_x_data_in42;
  wire [9:0] _kanwa_x_data_in43;
  wire [9:0] _kanwa_x_data_in44;
  wire [9:0] _kanwa_x_data_in45;
  wire [9:0] _kanwa_x_data_in46;
  wire [9:0] _kanwa_x_data_in47;
  wire [9:0] _kanwa_x_data_in48;
  wire [9:0] _kanwa_x_data_in49;
  wire [9:0] _kanwa_x_data_in50;
  wire [9:0] _kanwa_x_data_in51;
  wire [9:0] _kanwa_x_data_in52;
  wire [9:0] _kanwa_x_data_in53;
  wire [9:0] _kanwa_x_data_in54;
  wire [9:0] _kanwa_x_data_in55;
  wire [9:0] _kanwa_x_data_in56;
  wire [9:0] _kanwa_x_data_in57;
  wire [9:0] _kanwa_x_data_in58;
  wire [9:0] _kanwa_x_data_in59;
  wire [9:0] _kanwa_x_data_in60;
  wire [9:0] _kanwa_x_data_in61;
  wire [9:0] _kanwa_x_data_in62;
  wire [9:0] _kanwa_x_data_in65;
  wire [9:0] _kanwa_x_data_in66;
  wire [9:0] _kanwa_x_data_in67;
  wire [9:0] _kanwa_x_data_in68;
  wire [9:0] _kanwa_x_data_in69;
  wire [9:0] _kanwa_x_data_in70;
  wire [9:0] _kanwa_x_data_in71;
  wire [9:0] _kanwa_x_data_in72;
  wire [9:0] _kanwa_x_data_in73;
  wire [9:0] _kanwa_x_data_in74;
  wire [9:0] _kanwa_x_data_in75;
  wire [9:0] _kanwa_x_data_in76;
  wire [9:0] _kanwa_x_data_in77;
  wire [9:0] _kanwa_x_data_in78;
  wire [9:0] _kanwa_x_data_in79;
  wire [9:0] _kanwa_x_data_in80;
  wire [9:0] _kanwa_x_data_in81;
  wire [9:0] _kanwa_x_data_in82;
  wire [9:0] _kanwa_x_data_in83;
  wire [9:0] _kanwa_x_data_in84;
  wire [9:0] _kanwa_x_data_in85;
  wire [9:0] _kanwa_x_data_in86;
  wire [9:0] _kanwa_x_data_in87;
  wire [9:0] _kanwa_x_data_in88;
  wire [9:0] _kanwa_x_data_in89;
  wire [9:0] _kanwa_x_data_in90;
  wire [9:0] _kanwa_x_data_in91;
  wire [9:0] _kanwa_x_data_in92;
  wire [9:0] _kanwa_x_data_in93;
  wire [9:0] _kanwa_x_data_in94;
  wire [9:0] _kanwa_x_data_in97;
  wire [9:0] _kanwa_x_data_in98;
  wire [9:0] _kanwa_x_data_in99;
  wire [9:0] _kanwa_x_data_in100;
  wire [9:0] _kanwa_x_data_in101;
  wire [9:0] _kanwa_x_data_in102;
  wire [9:0] _kanwa_x_data_in103;
  wire [9:0] _kanwa_x_data_in104;
  wire [9:0] _kanwa_x_data_in105;
  wire [9:0] _kanwa_x_data_in106;
  wire [9:0] _kanwa_x_data_in107;
  wire [9:0] _kanwa_x_data_in108;
  wire [9:0] _kanwa_x_data_in109;
  wire [9:0] _kanwa_x_data_in110;
  wire [9:0] _kanwa_x_data_in111;
  wire [9:0] _kanwa_x_data_in112;
  wire [9:0] _kanwa_x_data_in113;
  wire [9:0] _kanwa_x_data_in114;
  wire [9:0] _kanwa_x_data_in115;
  wire [9:0] _kanwa_x_data_in116;
  wire [9:0] _kanwa_x_data_in117;
  wire [9:0] _kanwa_x_data_in118;
  wire [9:0] _kanwa_x_data_in119;
  wire [9:0] _kanwa_x_data_in120;
  wire [9:0] _kanwa_x_data_in121;
  wire [9:0] _kanwa_x_data_in122;
  wire [9:0] _kanwa_x_data_in123;
  wire [9:0] _kanwa_x_data_in124;
  wire [9:0] _kanwa_x_data_in125;
  wire [9:0] _kanwa_x_data_in126;
  wire [9:0] _kanwa_x_data_in129;
  wire [9:0] _kanwa_x_data_in130;
  wire [9:0] _kanwa_x_data_in131;
  wire [9:0] _kanwa_x_data_in132;
  wire [9:0] _kanwa_x_data_in133;
  wire [9:0] _kanwa_x_data_in134;
  wire [9:0] _kanwa_x_data_in135;
  wire [9:0] _kanwa_x_data_in136;
  wire [9:0] _kanwa_x_data_in137;
  wire [9:0] _kanwa_x_data_in138;
  wire [9:0] _kanwa_x_data_in139;
  wire [9:0] _kanwa_x_data_in140;
  wire [9:0] _kanwa_x_data_in141;
  wire [9:0] _kanwa_x_data_in142;
  wire [9:0] _kanwa_x_data_in143;
  wire [9:0] _kanwa_x_data_in144;
  wire [9:0] _kanwa_x_data_in145;
  wire [9:0] _kanwa_x_data_in146;
  wire [9:0] _kanwa_x_data_in147;
  wire [9:0] _kanwa_x_data_in148;
  wire [9:0] _kanwa_x_data_in149;
  wire [9:0] _kanwa_x_data_in150;
  wire [9:0] _kanwa_x_data_in151;
  wire [9:0] _kanwa_x_data_in152;
  wire [9:0] _kanwa_x_data_in153;
  wire [9:0] _kanwa_x_data_in154;
  wire [9:0] _kanwa_x_data_in155;
  wire [9:0] _kanwa_x_data_in156;
  wire [9:0] _kanwa_x_data_in157;
  wire [9:0] _kanwa_x_data_in158;
  wire [9:0] _kanwa_x_data_in161;
  wire [9:0] _kanwa_x_data_in162;
  wire [9:0] _kanwa_x_data_in163;
  wire [9:0] _kanwa_x_data_in164;
  wire [9:0] _kanwa_x_data_in165;
  wire [9:0] _kanwa_x_data_in166;
  wire [9:0] _kanwa_x_data_in167;
  wire [9:0] _kanwa_x_data_in168;
  wire [9:0] _kanwa_x_data_in169;
  wire [9:0] _kanwa_x_data_in170;
  wire [9:0] _kanwa_x_data_in171;
  wire [9:0] _kanwa_x_data_in172;
  wire [9:0] _kanwa_x_data_in173;
  wire [9:0] _kanwa_x_data_in174;
  wire [9:0] _kanwa_x_data_in175;
  wire [9:0] _kanwa_x_data_in176;
  wire [9:0] _kanwa_x_data_in177;
  wire [9:0] _kanwa_x_data_in178;
  wire [9:0] _kanwa_x_data_in179;
  wire [9:0] _kanwa_x_data_in180;
  wire [9:0] _kanwa_x_data_in181;
  wire [9:0] _kanwa_x_data_in182;
  wire [9:0] _kanwa_x_data_in183;
  wire [9:0] _kanwa_x_data_in184;
  wire [9:0] _kanwa_x_data_in185;
  wire [9:0] _kanwa_x_data_in186;
  wire [9:0] _kanwa_x_data_in187;
  wire [9:0] _kanwa_x_data_in188;
  wire [9:0] _kanwa_x_data_in189;
  wire [9:0] _kanwa_x_data_in190;
  wire [9:0] _kanwa_x_data_in193;
  wire [9:0] _kanwa_x_data_in194;
  wire [9:0] _kanwa_x_data_in195;
  wire [9:0] _kanwa_x_data_in196;
  wire [9:0] _kanwa_x_data_in197;
  wire [9:0] _kanwa_x_data_in198;
  wire [9:0] _kanwa_x_data_in199;
  wire [9:0] _kanwa_x_data_in200;
  wire [9:0] _kanwa_x_data_in201;
  wire [9:0] _kanwa_x_data_in202;
  wire [9:0] _kanwa_x_data_in203;
  wire [9:0] _kanwa_x_data_in204;
  wire [9:0] _kanwa_x_data_in205;
  wire [9:0] _kanwa_x_data_in206;
  wire [9:0] _kanwa_x_data_in207;
  wire [9:0] _kanwa_x_data_in208;
  wire [9:0] _kanwa_x_data_in209;
  wire [9:0] _kanwa_x_data_in210;
  wire [9:0] _kanwa_x_data_in211;
  wire [9:0] _kanwa_x_data_in212;
  wire [9:0] _kanwa_x_data_in213;
  wire [9:0] _kanwa_x_data_in214;
  wire [9:0] _kanwa_x_data_in215;
  wire [9:0] _kanwa_x_data_in216;
  wire [9:0] _kanwa_x_data_in217;
  wire [9:0] _kanwa_x_data_in218;
  wire [9:0] _kanwa_x_data_in219;
  wire [9:0] _kanwa_x_data_in220;
  wire [9:0] _kanwa_x_data_in221;
  wire [9:0] _kanwa_x_data_in222;
  wire [9:0] _kanwa_x_data_in225;
  wire [9:0] _kanwa_x_data_in226;
  wire [9:0] _kanwa_x_data_in227;
  wire [9:0] _kanwa_x_data_in228;
  wire [9:0] _kanwa_x_data_in229;
  wire [9:0] _kanwa_x_data_in230;
  wire [9:0] _kanwa_x_data_in231;
  wire [9:0] _kanwa_x_data_in232;
  wire [9:0] _kanwa_x_data_in233;
  wire [9:0] _kanwa_x_data_in234;
  wire [9:0] _kanwa_x_data_in235;
  wire [9:0] _kanwa_x_data_in236;
  wire [9:0] _kanwa_x_data_in237;
  wire [9:0] _kanwa_x_data_in238;
  wire [9:0] _kanwa_x_data_in239;
  wire [9:0] _kanwa_x_data_in240;
  wire [9:0] _kanwa_x_data_in241;
  wire [9:0] _kanwa_x_data_in242;
  wire [9:0] _kanwa_x_data_in243;
  wire [9:0] _kanwa_x_data_in244;
  wire [9:0] _kanwa_x_data_in245;
  wire [9:0] _kanwa_x_data_in246;
  wire [9:0] _kanwa_x_data_in247;
  wire [9:0] _kanwa_x_data_in248;
  wire [9:0] _kanwa_x_data_in249;
  wire [9:0] _kanwa_x_data_in250;
  wire [9:0] _kanwa_x_data_in251;
  wire [9:0] _kanwa_x_data_in252;
  wire [9:0] _kanwa_x_data_in253;
  wire [9:0] _kanwa_x_data_in254;
  wire [9:0] _kanwa_x_data_in257;
  wire [9:0] _kanwa_x_data_in258;
  wire [9:0] _kanwa_x_data_in259;
  wire [9:0] _kanwa_x_data_in260;
  wire [9:0] _kanwa_x_data_in261;
  wire [9:0] _kanwa_x_data_in262;
  wire [9:0] _kanwa_x_data_in263;
  wire [9:0] _kanwa_x_data_in264;
  wire [9:0] _kanwa_x_data_in265;
  wire [9:0] _kanwa_x_data_in266;
  wire [9:0] _kanwa_x_data_in267;
  wire [9:0] _kanwa_x_data_in268;
  wire [9:0] _kanwa_x_data_in269;
  wire [9:0] _kanwa_x_data_in270;
  wire [9:0] _kanwa_x_data_in271;
  wire [9:0] _kanwa_x_data_in272;
  wire [9:0] _kanwa_x_data_in273;
  wire [9:0] _kanwa_x_data_in274;
  wire [9:0] _kanwa_x_data_in275;
  wire [9:0] _kanwa_x_data_in276;
  wire [9:0] _kanwa_x_data_in277;
  wire [9:0] _kanwa_x_data_in278;
  wire [9:0] _kanwa_x_data_in279;
  wire [9:0] _kanwa_x_data_in280;
  wire [9:0] _kanwa_x_data_in281;
  wire [9:0] _kanwa_x_data_in282;
  wire [9:0] _kanwa_x_data_in283;
  wire [9:0] _kanwa_x_data_in284;
  wire [9:0] _kanwa_x_data_in285;
  wire [9:0] _kanwa_x_data_in286;
  wire [9:0] _kanwa_x_data_in289;
  wire [9:0] _kanwa_x_data_in290;
  wire [9:0] _kanwa_x_data_in291;
  wire [9:0] _kanwa_x_data_in292;
  wire [9:0] _kanwa_x_data_in293;
  wire [9:0] _kanwa_x_data_in294;
  wire [9:0] _kanwa_x_data_in295;
  wire [9:0] _kanwa_x_data_in296;
  wire [9:0] _kanwa_x_data_in297;
  wire [9:0] _kanwa_x_data_in298;
  wire [9:0] _kanwa_x_data_in299;
  wire [9:0] _kanwa_x_data_in300;
  wire [9:0] _kanwa_x_data_in301;
  wire [9:0] _kanwa_x_data_in302;
  wire [9:0] _kanwa_x_data_in303;
  wire [9:0] _kanwa_x_data_in304;
  wire [9:0] _kanwa_x_data_in305;
  wire [9:0] _kanwa_x_data_in306;
  wire [9:0] _kanwa_x_data_in307;
  wire [9:0] _kanwa_x_data_in308;
  wire [9:0] _kanwa_x_data_in309;
  wire [9:0] _kanwa_x_data_in310;
  wire [9:0] _kanwa_x_data_in311;
  wire [9:0] _kanwa_x_data_in312;
  wire [9:0] _kanwa_x_data_in313;
  wire [9:0] _kanwa_x_data_in314;
  wire [9:0] _kanwa_x_data_in315;
  wire [9:0] _kanwa_x_data_in316;
  wire [9:0] _kanwa_x_data_in317;
  wire [9:0] _kanwa_x_data_in318;
  wire [9:0] _kanwa_x_data_in321;
  wire [9:0] _kanwa_x_data_in322;
  wire [9:0] _kanwa_x_data_in323;
  wire [9:0] _kanwa_x_data_in324;
  wire [9:0] _kanwa_x_data_in325;
  wire [9:0] _kanwa_x_data_in326;
  wire [9:0] _kanwa_x_data_in327;
  wire [9:0] _kanwa_x_data_in328;
  wire [9:0] _kanwa_x_data_in329;
  wire [9:0] _kanwa_x_data_in330;
  wire [9:0] _kanwa_x_data_in331;
  wire [9:0] _kanwa_x_data_in332;
  wire [9:0] _kanwa_x_data_in333;
  wire [9:0] _kanwa_x_data_in334;
  wire [9:0] _kanwa_x_data_in335;
  wire [9:0] _kanwa_x_data_in336;
  wire [9:0] _kanwa_x_data_in337;
  wire [9:0] _kanwa_x_data_in338;
  wire [9:0] _kanwa_x_data_in339;
  wire [9:0] _kanwa_x_data_in340;
  wire [9:0] _kanwa_x_data_in341;
  wire [9:0] _kanwa_x_data_in342;
  wire [9:0] _kanwa_x_data_in343;
  wire [9:0] _kanwa_x_data_in344;
  wire [9:0] _kanwa_x_data_in345;
  wire [9:0] _kanwa_x_data_in346;
  wire [9:0] _kanwa_x_data_in347;
  wire [9:0] _kanwa_x_data_in348;
  wire [9:0] _kanwa_x_data_in349;
  wire [9:0] _kanwa_x_data_in350;
  wire [9:0] _kanwa_x_data_in353;
  wire [9:0] _kanwa_x_data_in354;
  wire [9:0] _kanwa_x_data_in355;
  wire [9:0] _kanwa_x_data_in356;
  wire [9:0] _kanwa_x_data_in357;
  wire [9:0] _kanwa_x_data_in358;
  wire [9:0] _kanwa_x_data_in359;
  wire [9:0] _kanwa_x_data_in360;
  wire [9:0] _kanwa_x_data_in361;
  wire [9:0] _kanwa_x_data_in362;
  wire [9:0] _kanwa_x_data_in363;
  wire [9:0] _kanwa_x_data_in364;
  wire [9:0] _kanwa_x_data_in365;
  wire [9:0] _kanwa_x_data_in366;
  wire [9:0] _kanwa_x_data_in367;
  wire [9:0] _kanwa_x_data_in368;
  wire [9:0] _kanwa_x_data_in369;
  wire [9:0] _kanwa_x_data_in370;
  wire [9:0] _kanwa_x_data_in371;
  wire [9:0] _kanwa_x_data_in372;
  wire [9:0] _kanwa_x_data_in373;
  wire [9:0] _kanwa_x_data_in374;
  wire [9:0] _kanwa_x_data_in375;
  wire [9:0] _kanwa_x_data_in376;
  wire [9:0] _kanwa_x_data_in377;
  wire [9:0] _kanwa_x_data_in378;
  wire [9:0] _kanwa_x_data_in379;
  wire [9:0] _kanwa_x_data_in380;
  wire [9:0] _kanwa_x_data_in381;
  wire [9:0] _kanwa_x_data_in382;
  wire [9:0] _kanwa_x_data_in385;
  wire [9:0] _kanwa_x_data_in386;
  wire [9:0] _kanwa_x_data_in387;
  wire [9:0] _kanwa_x_data_in388;
  wire [9:0] _kanwa_x_data_in389;
  wire [9:0] _kanwa_x_data_in390;
  wire [9:0] _kanwa_x_data_in391;
  wire [9:0] _kanwa_x_data_in392;
  wire [9:0] _kanwa_x_data_in393;
  wire [9:0] _kanwa_x_data_in394;
  wire [9:0] _kanwa_x_data_in395;
  wire [9:0] _kanwa_x_data_in396;
  wire [9:0] _kanwa_x_data_in397;
  wire [9:0] _kanwa_x_data_in398;
  wire [9:0] _kanwa_x_data_in399;
  wire [9:0] _kanwa_x_data_in400;
  wire [9:0] _kanwa_x_data_in401;
  wire [9:0] _kanwa_x_data_in402;
  wire [9:0] _kanwa_x_data_in403;
  wire [9:0] _kanwa_x_data_in404;
  wire [9:0] _kanwa_x_data_in405;
  wire [9:0] _kanwa_x_data_in406;
  wire [9:0] _kanwa_x_data_in407;
  wire [9:0] _kanwa_x_data_in408;
  wire [9:0] _kanwa_x_data_in409;
  wire [9:0] _kanwa_x_data_in410;
  wire [9:0] _kanwa_x_data_in411;
  wire [9:0] _kanwa_x_data_in412;
  wire [9:0] _kanwa_x_data_in413;
  wire [9:0] _kanwa_x_data_in414;
  wire [9:0] _kanwa_x_data_in417;
  wire [9:0] _kanwa_x_data_in418;
  wire [9:0] _kanwa_x_data_in419;
  wire [9:0] _kanwa_x_data_in420;
  wire [9:0] _kanwa_x_data_in421;
  wire [9:0] _kanwa_x_data_in422;
  wire [9:0] _kanwa_x_data_in423;
  wire [9:0] _kanwa_x_data_in424;
  wire [9:0] _kanwa_x_data_in425;
  wire [9:0] _kanwa_x_data_in426;
  wire [9:0] _kanwa_x_data_in427;
  wire [9:0] _kanwa_x_data_in428;
  wire [9:0] _kanwa_x_data_in429;
  wire [9:0] _kanwa_x_data_in430;
  wire [9:0] _kanwa_x_data_in431;
  wire [9:0] _kanwa_x_data_in432;
  wire [9:0] _kanwa_x_data_in433;
  wire [9:0] _kanwa_x_data_in434;
  wire [9:0] _kanwa_x_data_in435;
  wire [9:0] _kanwa_x_data_in436;
  wire [9:0] _kanwa_x_data_in437;
  wire [9:0] _kanwa_x_data_in438;
  wire [9:0] _kanwa_x_data_in439;
  wire [9:0] _kanwa_x_data_in440;
  wire [9:0] _kanwa_x_data_in441;
  wire [9:0] _kanwa_x_data_in442;
  wire [9:0] _kanwa_x_data_in443;
  wire [9:0] _kanwa_x_data_in444;
  wire [9:0] _kanwa_x_data_in445;
  wire [9:0] _kanwa_x_data_in446;
  wire [9:0] _kanwa_x_data_in449;
  wire [9:0] _kanwa_x_data_in450;
  wire [9:0] _kanwa_x_data_in451;
  wire [9:0] _kanwa_x_data_in452;
  wire [9:0] _kanwa_x_data_in453;
  wire [9:0] _kanwa_x_data_in454;
  wire [9:0] _kanwa_x_data_in455;
  wire [9:0] _kanwa_x_data_in456;
  wire [9:0] _kanwa_x_data_in457;
  wire [9:0] _kanwa_x_data_in458;
  wire [9:0] _kanwa_x_data_in459;
  wire [9:0] _kanwa_x_data_in460;
  wire [9:0] _kanwa_x_data_in461;
  wire [9:0] _kanwa_x_data_in462;
  wire [9:0] _kanwa_x_data_in463;
  wire [9:0] _kanwa_x_data_in464;
  wire [9:0] _kanwa_x_data_in465;
  wire [9:0] _kanwa_x_data_in466;
  wire [9:0] _kanwa_x_data_in467;
  wire [9:0] _kanwa_x_data_in468;
  wire [9:0] _kanwa_x_data_in469;
  wire [9:0] _kanwa_x_data_in470;
  wire [9:0] _kanwa_x_data_in471;
  wire [9:0] _kanwa_x_data_in472;
  wire [9:0] _kanwa_x_data_in473;
  wire [9:0] _kanwa_x_data_in474;
  wire [9:0] _kanwa_x_data_in475;
  wire [9:0] _kanwa_x_data_in476;
  wire [9:0] _kanwa_x_data_in477;
  wire [9:0] _kanwa_x_data_in478;
  wire [9:0] _kanwa_x_start;
  wire [9:0] _kanwa_x_goal;
  wire [9:0] _kanwa_x_data_out33;
  wire [9:0] _kanwa_x_data_out34;
  wire [9:0] _kanwa_x_data_out35;
  wire [9:0] _kanwa_x_data_out36;
  wire [9:0] _kanwa_x_data_out37;
  wire [9:0] _kanwa_x_data_out38;
  wire [9:0] _kanwa_x_data_out39;
  wire [9:0] _kanwa_x_data_out40;
  wire [9:0] _kanwa_x_data_out41;
  wire [9:0] _kanwa_x_data_out42;
  wire [9:0] _kanwa_x_data_out43;
  wire [9:0] _kanwa_x_data_out44;
  wire [9:0] _kanwa_x_data_out45;
  wire [9:0] _kanwa_x_data_out46;
  wire [9:0] _kanwa_x_data_out47;
  wire [9:0] _kanwa_x_data_out48;
  wire [9:0] _kanwa_x_data_out49;
  wire [9:0] _kanwa_x_data_out50;
  wire [9:0] _kanwa_x_data_out51;
  wire [9:0] _kanwa_x_data_out52;
  wire [9:0] _kanwa_x_data_out53;
  wire [9:0] _kanwa_x_data_out54;
  wire [9:0] _kanwa_x_data_out55;
  wire [9:0] _kanwa_x_data_out56;
  wire [9:0] _kanwa_x_data_out57;
  wire [9:0] _kanwa_x_data_out58;
  wire [9:0] _kanwa_x_data_out59;
  wire [9:0] _kanwa_x_data_out60;
  wire [9:0] _kanwa_x_data_out61;
  wire [9:0] _kanwa_x_data_out62;
  wire [9:0] _kanwa_x_data_out65;
  wire [9:0] _kanwa_x_data_out66;
  wire [9:0] _kanwa_x_data_out67;
  wire [9:0] _kanwa_x_data_out68;
  wire [9:0] _kanwa_x_data_out69;
  wire [9:0] _kanwa_x_data_out70;
  wire [9:0] _kanwa_x_data_out71;
  wire [9:0] _kanwa_x_data_out72;
  wire [9:0] _kanwa_x_data_out73;
  wire [9:0] _kanwa_x_data_out74;
  wire [9:0] _kanwa_x_data_out75;
  wire [9:0] _kanwa_x_data_out76;
  wire [9:0] _kanwa_x_data_out77;
  wire [9:0] _kanwa_x_data_out78;
  wire [9:0] _kanwa_x_data_out79;
  wire [9:0] _kanwa_x_data_out80;
  wire [9:0] _kanwa_x_data_out81;
  wire [9:0] _kanwa_x_data_out82;
  wire [9:0] _kanwa_x_data_out83;
  wire [9:0] _kanwa_x_data_out84;
  wire [9:0] _kanwa_x_data_out85;
  wire [9:0] _kanwa_x_data_out86;
  wire [9:0] _kanwa_x_data_out87;
  wire [9:0] _kanwa_x_data_out88;
  wire [9:0] _kanwa_x_data_out89;
  wire [9:0] _kanwa_x_data_out90;
  wire [9:0] _kanwa_x_data_out91;
  wire [9:0] _kanwa_x_data_out92;
  wire [9:0] _kanwa_x_data_out93;
  wire [9:0] _kanwa_x_data_out94;
  wire [9:0] _kanwa_x_data_out97;
  wire [9:0] _kanwa_x_data_out98;
  wire [9:0] _kanwa_x_data_out99;
  wire [9:0] _kanwa_x_data_out100;
  wire [9:0] _kanwa_x_data_out101;
  wire [9:0] _kanwa_x_data_out102;
  wire [9:0] _kanwa_x_data_out103;
  wire [9:0] _kanwa_x_data_out104;
  wire [9:0] _kanwa_x_data_out105;
  wire [9:0] _kanwa_x_data_out106;
  wire [9:0] _kanwa_x_data_out107;
  wire [9:0] _kanwa_x_data_out108;
  wire [9:0] _kanwa_x_data_out109;
  wire [9:0] _kanwa_x_data_out110;
  wire [9:0] _kanwa_x_data_out111;
  wire [9:0] _kanwa_x_data_out112;
  wire [9:0] _kanwa_x_data_out113;
  wire [9:0] _kanwa_x_data_out114;
  wire [9:0] _kanwa_x_data_out115;
  wire [9:0] _kanwa_x_data_out116;
  wire [9:0] _kanwa_x_data_out117;
  wire [9:0] _kanwa_x_data_out118;
  wire [9:0] _kanwa_x_data_out119;
  wire [9:0] _kanwa_x_data_out120;
  wire [9:0] _kanwa_x_data_out121;
  wire [9:0] _kanwa_x_data_out122;
  wire [9:0] _kanwa_x_data_out123;
  wire [9:0] _kanwa_x_data_out124;
  wire [9:0] _kanwa_x_data_out125;
  wire [9:0] _kanwa_x_data_out126;
  wire [9:0] _kanwa_x_data_out129;
  wire [9:0] _kanwa_x_data_out130;
  wire [9:0] _kanwa_x_data_out131;
  wire [9:0] _kanwa_x_data_out132;
  wire [9:0] _kanwa_x_data_out133;
  wire [9:0] _kanwa_x_data_out134;
  wire [9:0] _kanwa_x_data_out135;
  wire [9:0] _kanwa_x_data_out136;
  wire [9:0] _kanwa_x_data_out137;
  wire [9:0] _kanwa_x_data_out138;
  wire [9:0] _kanwa_x_data_out139;
  wire [9:0] _kanwa_x_data_out140;
  wire [9:0] _kanwa_x_data_out141;
  wire [9:0] _kanwa_x_data_out142;
  wire [9:0] _kanwa_x_data_out143;
  wire [9:0] _kanwa_x_data_out144;
  wire [9:0] _kanwa_x_data_out145;
  wire [9:0] _kanwa_x_data_out146;
  wire [9:0] _kanwa_x_data_out147;
  wire [9:0] _kanwa_x_data_out148;
  wire [9:0] _kanwa_x_data_out149;
  wire [9:0] _kanwa_x_data_out150;
  wire [9:0] _kanwa_x_data_out151;
  wire [9:0] _kanwa_x_data_out152;
  wire [9:0] _kanwa_x_data_out153;
  wire [9:0] _kanwa_x_data_out154;
  wire [9:0] _kanwa_x_data_out155;
  wire [9:0] _kanwa_x_data_out156;
  wire [9:0] _kanwa_x_data_out157;
  wire [9:0] _kanwa_x_data_out158;
  wire [9:0] _kanwa_x_data_out161;
  wire [9:0] _kanwa_x_data_out162;
  wire [9:0] _kanwa_x_data_out163;
  wire [9:0] _kanwa_x_data_out164;
  wire [9:0] _kanwa_x_data_out165;
  wire [9:0] _kanwa_x_data_out166;
  wire [9:0] _kanwa_x_data_out167;
  wire [9:0] _kanwa_x_data_out168;
  wire [9:0] _kanwa_x_data_out169;
  wire [9:0] _kanwa_x_data_out170;
  wire [9:0] _kanwa_x_data_out171;
  wire [9:0] _kanwa_x_data_out172;
  wire [9:0] _kanwa_x_data_out173;
  wire [9:0] _kanwa_x_data_out174;
  wire [9:0] _kanwa_x_data_out175;
  wire [9:0] _kanwa_x_data_out176;
  wire [9:0] _kanwa_x_data_out177;
  wire [9:0] _kanwa_x_data_out178;
  wire [9:0] _kanwa_x_data_out179;
  wire [9:0] _kanwa_x_data_out180;
  wire [9:0] _kanwa_x_data_out181;
  wire [9:0] _kanwa_x_data_out182;
  wire [9:0] _kanwa_x_data_out183;
  wire [9:0] _kanwa_x_data_out184;
  wire [9:0] _kanwa_x_data_out185;
  wire [9:0] _kanwa_x_data_out186;
  wire [9:0] _kanwa_x_data_out187;
  wire [9:0] _kanwa_x_data_out188;
  wire [9:0] _kanwa_x_data_out189;
  wire [9:0] _kanwa_x_data_out190;
  wire [9:0] _kanwa_x_data_out193;
  wire [9:0] _kanwa_x_data_out194;
  wire [9:0] _kanwa_x_data_out195;
  wire [9:0] _kanwa_x_data_out196;
  wire [9:0] _kanwa_x_data_out197;
  wire [9:0] _kanwa_x_data_out198;
  wire [9:0] _kanwa_x_data_out199;
  wire [9:0] _kanwa_x_data_out200;
  wire [9:0] _kanwa_x_data_out201;
  wire [9:0] _kanwa_x_data_out202;
  wire [9:0] _kanwa_x_data_out203;
  wire [9:0] _kanwa_x_data_out204;
  wire [9:0] _kanwa_x_data_out205;
  wire [9:0] _kanwa_x_data_out206;
  wire [9:0] _kanwa_x_data_out207;
  wire [9:0] _kanwa_x_data_out208;
  wire [9:0] _kanwa_x_data_out209;
  wire [9:0] _kanwa_x_data_out210;
  wire [9:0] _kanwa_x_data_out211;
  wire [9:0] _kanwa_x_data_out212;
  wire [9:0] _kanwa_x_data_out213;
  wire [9:0] _kanwa_x_data_out214;
  wire [9:0] _kanwa_x_data_out215;
  wire [9:0] _kanwa_x_data_out216;
  wire [9:0] _kanwa_x_data_out217;
  wire [9:0] _kanwa_x_data_out218;
  wire [9:0] _kanwa_x_data_out219;
  wire [9:0] _kanwa_x_data_out220;
  wire [9:0] _kanwa_x_data_out221;
  wire [9:0] _kanwa_x_data_out222;
  wire [9:0] _kanwa_x_data_out225;
  wire [9:0] _kanwa_x_data_out226;
  wire [9:0] _kanwa_x_data_out227;
  wire [9:0] _kanwa_x_data_out228;
  wire [9:0] _kanwa_x_data_out229;
  wire [9:0] _kanwa_x_data_out230;
  wire [9:0] _kanwa_x_data_out231;
  wire [9:0] _kanwa_x_data_out232;
  wire [9:0] _kanwa_x_data_out233;
  wire [9:0] _kanwa_x_data_out234;
  wire [9:0] _kanwa_x_data_out235;
  wire [9:0] _kanwa_x_data_out236;
  wire [9:0] _kanwa_x_data_out237;
  wire [9:0] _kanwa_x_data_out238;
  wire [9:0] _kanwa_x_data_out239;
  wire [9:0] _kanwa_x_data_out240;
  wire [9:0] _kanwa_x_data_out241;
  wire [9:0] _kanwa_x_data_out242;
  wire [9:0] _kanwa_x_data_out243;
  wire [9:0] _kanwa_x_data_out244;
  wire [9:0] _kanwa_x_data_out245;
  wire [9:0] _kanwa_x_data_out246;
  wire [9:0] _kanwa_x_data_out247;
  wire [9:0] _kanwa_x_data_out248;
  wire [9:0] _kanwa_x_data_out249;
  wire [9:0] _kanwa_x_data_out250;
  wire [9:0] _kanwa_x_data_out251;
  wire [9:0] _kanwa_x_data_out252;
  wire [9:0] _kanwa_x_data_out253;
  wire [9:0] _kanwa_x_data_out254;
  wire [9:0] _kanwa_x_data_out257;
  wire [9:0] _kanwa_x_data_out258;
  wire [9:0] _kanwa_x_data_out259;
  wire [9:0] _kanwa_x_data_out260;
  wire [9:0] _kanwa_x_data_out261;
  wire [9:0] _kanwa_x_data_out262;
  wire [9:0] _kanwa_x_data_out263;
  wire [9:0] _kanwa_x_data_out264;
  wire [9:0] _kanwa_x_data_out265;
  wire [9:0] _kanwa_x_data_out266;
  wire [9:0] _kanwa_x_data_out267;
  wire [9:0] _kanwa_x_data_out268;
  wire [9:0] _kanwa_x_data_out269;
  wire [9:0] _kanwa_x_data_out270;
  wire [9:0] _kanwa_x_data_out271;
  wire [9:0] _kanwa_x_data_out272;
  wire [9:0] _kanwa_x_data_out273;
  wire [9:0] _kanwa_x_data_out274;
  wire [9:0] _kanwa_x_data_out275;
  wire [9:0] _kanwa_x_data_out276;
  wire [9:0] _kanwa_x_data_out277;
  wire [9:0] _kanwa_x_data_out278;
  wire [9:0] _kanwa_x_data_out279;
  wire [9:0] _kanwa_x_data_out280;
  wire [9:0] _kanwa_x_data_out281;
  wire [9:0] _kanwa_x_data_out282;
  wire [9:0] _kanwa_x_data_out283;
  wire [9:0] _kanwa_x_data_out284;
  wire [9:0] _kanwa_x_data_out285;
  wire [9:0] _kanwa_x_data_out286;
  wire [9:0] _kanwa_x_data_out289;
  wire [9:0] _kanwa_x_data_out290;
  wire [9:0] _kanwa_x_data_out291;
  wire [9:0] _kanwa_x_data_out292;
  wire [9:0] _kanwa_x_data_out293;
  wire [9:0] _kanwa_x_data_out294;
  wire [9:0] _kanwa_x_data_out295;
  wire [9:0] _kanwa_x_data_out296;
  wire [9:0] _kanwa_x_data_out297;
  wire [9:0] _kanwa_x_data_out298;
  wire [9:0] _kanwa_x_data_out299;
  wire [9:0] _kanwa_x_data_out300;
  wire [9:0] _kanwa_x_data_out301;
  wire [9:0] _kanwa_x_data_out302;
  wire [9:0] _kanwa_x_data_out303;
  wire [9:0] _kanwa_x_data_out304;
  wire [9:0] _kanwa_x_data_out305;
  wire [9:0] _kanwa_x_data_out306;
  wire [9:0] _kanwa_x_data_out307;
  wire [9:0] _kanwa_x_data_out308;
  wire [9:0] _kanwa_x_data_out309;
  wire [9:0] _kanwa_x_data_out310;
  wire [9:0] _kanwa_x_data_out311;
  wire [9:0] _kanwa_x_data_out312;
  wire [9:0] _kanwa_x_data_out313;
  wire [9:0] _kanwa_x_data_out314;
  wire [9:0] _kanwa_x_data_out315;
  wire [9:0] _kanwa_x_data_out316;
  wire [9:0] _kanwa_x_data_out317;
  wire [9:0] _kanwa_x_data_out318;
  wire [9:0] _kanwa_x_data_out321;
  wire [9:0] _kanwa_x_data_out322;
  wire [9:0] _kanwa_x_data_out323;
  wire [9:0] _kanwa_x_data_out324;
  wire [9:0] _kanwa_x_data_out325;
  wire [9:0] _kanwa_x_data_out326;
  wire [9:0] _kanwa_x_data_out327;
  wire [9:0] _kanwa_x_data_out328;
  wire [9:0] _kanwa_x_data_out329;
  wire [9:0] _kanwa_x_data_out330;
  wire [9:0] _kanwa_x_data_out331;
  wire [9:0] _kanwa_x_data_out332;
  wire [9:0] _kanwa_x_data_out333;
  wire [9:0] _kanwa_x_data_out334;
  wire [9:0] _kanwa_x_data_out335;
  wire [9:0] _kanwa_x_data_out336;
  wire [9:0] _kanwa_x_data_out337;
  wire [9:0] _kanwa_x_data_out338;
  wire [9:0] _kanwa_x_data_out339;
  wire [9:0] _kanwa_x_data_out340;
  wire [9:0] _kanwa_x_data_out341;
  wire [9:0] _kanwa_x_data_out342;
  wire [9:0] _kanwa_x_data_out343;
  wire [9:0] _kanwa_x_data_out344;
  wire [9:0] _kanwa_x_data_out345;
  wire [9:0] _kanwa_x_data_out346;
  wire [9:0] _kanwa_x_data_out347;
  wire [9:0] _kanwa_x_data_out348;
  wire [9:0] _kanwa_x_data_out349;
  wire [9:0] _kanwa_x_data_out350;
  wire [9:0] _kanwa_x_data_out353;
  wire [9:0] _kanwa_x_data_out354;
  wire [9:0] _kanwa_x_data_out355;
  wire [9:0] _kanwa_x_data_out356;
  wire [9:0] _kanwa_x_data_out357;
  wire [9:0] _kanwa_x_data_out358;
  wire [9:0] _kanwa_x_data_out359;
  wire [9:0] _kanwa_x_data_out360;
  wire [9:0] _kanwa_x_data_out361;
  wire [9:0] _kanwa_x_data_out362;
  wire [9:0] _kanwa_x_data_out363;
  wire [9:0] _kanwa_x_data_out364;
  wire [9:0] _kanwa_x_data_out365;
  wire [9:0] _kanwa_x_data_out366;
  wire [9:0] _kanwa_x_data_out367;
  wire [9:0] _kanwa_x_data_out368;
  wire [9:0] _kanwa_x_data_out369;
  wire [9:0] _kanwa_x_data_out370;
  wire [9:0] _kanwa_x_data_out371;
  wire [9:0] _kanwa_x_data_out372;
  wire [9:0] _kanwa_x_data_out373;
  wire [9:0] _kanwa_x_data_out374;
  wire [9:0] _kanwa_x_data_out375;
  wire [9:0] _kanwa_x_data_out376;
  wire [9:0] _kanwa_x_data_out377;
  wire [9:0] _kanwa_x_data_out378;
  wire [9:0] _kanwa_x_data_out379;
  wire [9:0] _kanwa_x_data_out380;
  wire [9:0] _kanwa_x_data_out381;
  wire [9:0] _kanwa_x_data_out382;
  wire [9:0] _kanwa_x_data_out385;
  wire [9:0] _kanwa_x_data_out386;
  wire [9:0] _kanwa_x_data_out387;
  wire [9:0] _kanwa_x_data_out388;
  wire [9:0] _kanwa_x_data_out389;
  wire [9:0] _kanwa_x_data_out390;
  wire [9:0] _kanwa_x_data_out391;
  wire [9:0] _kanwa_x_data_out392;
  wire [9:0] _kanwa_x_data_out393;
  wire [9:0] _kanwa_x_data_out394;
  wire [9:0] _kanwa_x_data_out395;
  wire [9:0] _kanwa_x_data_out396;
  wire [9:0] _kanwa_x_data_out397;
  wire [9:0] _kanwa_x_data_out398;
  wire [9:0] _kanwa_x_data_out399;
  wire [9:0] _kanwa_x_data_out400;
  wire [9:0] _kanwa_x_data_out401;
  wire [9:0] _kanwa_x_data_out402;
  wire [9:0] _kanwa_x_data_out403;
  wire [9:0] _kanwa_x_data_out404;
  wire [9:0] _kanwa_x_data_out405;
  wire [9:0] _kanwa_x_data_out406;
  wire [9:0] _kanwa_x_data_out407;
  wire [9:0] _kanwa_x_data_out408;
  wire [9:0] _kanwa_x_data_out409;
  wire [9:0] _kanwa_x_data_out410;
  wire [9:0] _kanwa_x_data_out411;
  wire [9:0] _kanwa_x_data_out412;
  wire [9:0] _kanwa_x_data_out413;
  wire [9:0] _kanwa_x_data_out414;
  wire [9:0] _kanwa_x_data_out417;
  wire [9:0] _kanwa_x_data_out418;
  wire [9:0] _kanwa_x_data_out419;
  wire [9:0] _kanwa_x_data_out420;
  wire [9:0] _kanwa_x_data_out421;
  wire [9:0] _kanwa_x_data_out422;
  wire [9:0] _kanwa_x_data_out423;
  wire [9:0] _kanwa_x_data_out424;
  wire [9:0] _kanwa_x_data_out425;
  wire [9:0] _kanwa_x_data_out426;
  wire [9:0] _kanwa_x_data_out427;
  wire [9:0] _kanwa_x_data_out428;
  wire [9:0] _kanwa_x_data_out429;
  wire [9:0] _kanwa_x_data_out430;
  wire [9:0] _kanwa_x_data_out431;
  wire [9:0] _kanwa_x_data_out432;
  wire [9:0] _kanwa_x_data_out433;
  wire [9:0] _kanwa_x_data_out434;
  wire [9:0] _kanwa_x_data_out435;
  wire [9:0] _kanwa_x_data_out436;
  wire [9:0] _kanwa_x_data_out437;
  wire [9:0] _kanwa_x_data_out438;
  wire [9:0] _kanwa_x_data_out439;
  wire [9:0] _kanwa_x_data_out440;
  wire [9:0] _kanwa_x_data_out441;
  wire [9:0] _kanwa_x_data_out442;
  wire [9:0] _kanwa_x_data_out443;
  wire [9:0] _kanwa_x_data_out444;
  wire [9:0] _kanwa_x_data_out445;
  wire [9:0] _kanwa_x_data_out446;
  wire [9:0] _kanwa_x_data_out449;
  wire [9:0] _kanwa_x_data_out450;
  wire [9:0] _kanwa_x_data_out451;
  wire [9:0] _kanwa_x_data_out452;
  wire [9:0] _kanwa_x_data_out453;
  wire [9:0] _kanwa_x_data_out454;
  wire [9:0] _kanwa_x_data_out455;
  wire [9:0] _kanwa_x_data_out456;
  wire [9:0] _kanwa_x_data_out457;
  wire [9:0] _kanwa_x_data_out458;
  wire [9:0] _kanwa_x_data_out459;
  wire [9:0] _kanwa_x_data_out460;
  wire [9:0] _kanwa_x_data_out461;
  wire [9:0] _kanwa_x_data_out462;
  wire [9:0] _kanwa_x_data_out463;
  wire [9:0] _kanwa_x_data_out464;
  wire [9:0] _kanwa_x_data_out465;
  wire [9:0] _kanwa_x_data_out466;
  wire [9:0] _kanwa_x_data_out467;
  wire [9:0] _kanwa_x_data_out468;
  wire [9:0] _kanwa_x_data_out469;
  wire [9:0] _kanwa_x_data_out470;
  wire [9:0] _kanwa_x_data_out471;
  wire [9:0] _kanwa_x_data_out472;
  wire [9:0] _kanwa_x_data_out473;
  wire [9:0] _kanwa_x_data_out474;
  wire [9:0] _kanwa_x_data_out475;
  wire [9:0] _kanwa_x_data_out476;
  wire [9:0] _kanwa_x_data_out477;
  wire [9:0] _kanwa_x_data_out478;
  wire _kanwa_x_in_do;
  wire _kanwa_x_out_do;
  wire _kanwa_x_p_reset;
  wire _kanwa_x_m_clock;
  wire [9:0] _kouka_x_data_in33;
  wire [9:0] _kouka_x_data_in34;
  wire [9:0] _kouka_x_data_in35;
  wire [9:0] _kouka_x_data_in36;
  wire [9:0] _kouka_x_data_in37;
  wire [9:0] _kouka_x_data_in38;
  wire [9:0] _kouka_x_data_in39;
  wire [9:0] _kouka_x_data_in40;
  wire [9:0] _kouka_x_data_in41;
  wire [9:0] _kouka_x_data_in42;
  wire [9:0] _kouka_x_data_in43;
  wire [9:0] _kouka_x_data_in44;
  wire [9:0] _kouka_x_data_in45;
  wire [9:0] _kouka_x_data_in46;
  wire [9:0] _kouka_x_data_in47;
  wire [9:0] _kouka_x_data_in48;
  wire [9:0] _kouka_x_data_in49;
  wire [9:0] _kouka_x_data_in50;
  wire [9:0] _kouka_x_data_in51;
  wire [9:0] _kouka_x_data_in52;
  wire [9:0] _kouka_x_data_in53;
  wire [9:0] _kouka_x_data_in54;
  wire [9:0] _kouka_x_data_in55;
  wire [9:0] _kouka_x_data_in56;
  wire [9:0] _kouka_x_data_in57;
  wire [9:0] _kouka_x_data_in58;
  wire [9:0] _kouka_x_data_in59;
  wire [9:0] _kouka_x_data_in60;
  wire [9:0] _kouka_x_data_in61;
  wire [9:0] _kouka_x_data_in62;
  wire [9:0] _kouka_x_data_in65;
  wire [9:0] _kouka_x_data_in66;
  wire [9:0] _kouka_x_data_in67;
  wire [9:0] _kouka_x_data_in68;
  wire [9:0] _kouka_x_data_in69;
  wire [9:0] _kouka_x_data_in70;
  wire [9:0] _kouka_x_data_in71;
  wire [9:0] _kouka_x_data_in72;
  wire [9:0] _kouka_x_data_in73;
  wire [9:0] _kouka_x_data_in74;
  wire [9:0] _kouka_x_data_in75;
  wire [9:0] _kouka_x_data_in76;
  wire [9:0] _kouka_x_data_in77;
  wire [9:0] _kouka_x_data_in78;
  wire [9:0] _kouka_x_data_in79;
  wire [9:0] _kouka_x_data_in80;
  wire [9:0] _kouka_x_data_in81;
  wire [9:0] _kouka_x_data_in82;
  wire [9:0] _kouka_x_data_in83;
  wire [9:0] _kouka_x_data_in84;
  wire [9:0] _kouka_x_data_in85;
  wire [9:0] _kouka_x_data_in86;
  wire [9:0] _kouka_x_data_in87;
  wire [9:0] _kouka_x_data_in88;
  wire [9:0] _kouka_x_data_in89;
  wire [9:0] _kouka_x_data_in90;
  wire [9:0] _kouka_x_data_in91;
  wire [9:0] _kouka_x_data_in92;
  wire [9:0] _kouka_x_data_in93;
  wire [9:0] _kouka_x_data_in94;
  wire [9:0] _kouka_x_data_in97;
  wire [9:0] _kouka_x_data_in98;
  wire [9:0] _kouka_x_data_in99;
  wire [9:0] _kouka_x_data_in100;
  wire [9:0] _kouka_x_data_in101;
  wire [9:0] _kouka_x_data_in102;
  wire [9:0] _kouka_x_data_in103;
  wire [9:0] _kouka_x_data_in104;
  wire [9:0] _kouka_x_data_in105;
  wire [9:0] _kouka_x_data_in106;
  wire [9:0] _kouka_x_data_in107;
  wire [9:0] _kouka_x_data_in108;
  wire [9:0] _kouka_x_data_in109;
  wire [9:0] _kouka_x_data_in110;
  wire [9:0] _kouka_x_data_in111;
  wire [9:0] _kouka_x_data_in112;
  wire [9:0] _kouka_x_data_in113;
  wire [9:0] _kouka_x_data_in114;
  wire [9:0] _kouka_x_data_in115;
  wire [9:0] _kouka_x_data_in116;
  wire [9:0] _kouka_x_data_in117;
  wire [9:0] _kouka_x_data_in118;
  wire [9:0] _kouka_x_data_in119;
  wire [9:0] _kouka_x_data_in120;
  wire [9:0] _kouka_x_data_in121;
  wire [9:0] _kouka_x_data_in122;
  wire [9:0] _kouka_x_data_in123;
  wire [9:0] _kouka_x_data_in124;
  wire [9:0] _kouka_x_data_in125;
  wire [9:0] _kouka_x_data_in126;
  wire [9:0] _kouka_x_data_in129;
  wire [9:0] _kouka_x_data_in130;
  wire [9:0] _kouka_x_data_in131;
  wire [9:0] _kouka_x_data_in132;
  wire [9:0] _kouka_x_data_in133;
  wire [9:0] _kouka_x_data_in134;
  wire [9:0] _kouka_x_data_in135;
  wire [9:0] _kouka_x_data_in136;
  wire [9:0] _kouka_x_data_in137;
  wire [9:0] _kouka_x_data_in138;
  wire [9:0] _kouka_x_data_in139;
  wire [9:0] _kouka_x_data_in140;
  wire [9:0] _kouka_x_data_in141;
  wire [9:0] _kouka_x_data_in142;
  wire [9:0] _kouka_x_data_in143;
  wire [9:0] _kouka_x_data_in144;
  wire [9:0] _kouka_x_data_in145;
  wire [9:0] _kouka_x_data_in146;
  wire [9:0] _kouka_x_data_in147;
  wire [9:0] _kouka_x_data_in148;
  wire [9:0] _kouka_x_data_in149;
  wire [9:0] _kouka_x_data_in150;
  wire [9:0] _kouka_x_data_in151;
  wire [9:0] _kouka_x_data_in152;
  wire [9:0] _kouka_x_data_in153;
  wire [9:0] _kouka_x_data_in154;
  wire [9:0] _kouka_x_data_in155;
  wire [9:0] _kouka_x_data_in156;
  wire [9:0] _kouka_x_data_in157;
  wire [9:0] _kouka_x_data_in158;
  wire [9:0] _kouka_x_data_in161;
  wire [9:0] _kouka_x_data_in162;
  wire [9:0] _kouka_x_data_in163;
  wire [9:0] _kouka_x_data_in164;
  wire [9:0] _kouka_x_data_in165;
  wire [9:0] _kouka_x_data_in166;
  wire [9:0] _kouka_x_data_in167;
  wire [9:0] _kouka_x_data_in168;
  wire [9:0] _kouka_x_data_in169;
  wire [9:0] _kouka_x_data_in170;
  wire [9:0] _kouka_x_data_in171;
  wire [9:0] _kouka_x_data_in172;
  wire [9:0] _kouka_x_data_in173;
  wire [9:0] _kouka_x_data_in174;
  wire [9:0] _kouka_x_data_in175;
  wire [9:0] _kouka_x_data_in176;
  wire [9:0] _kouka_x_data_in177;
  wire [9:0] _kouka_x_data_in178;
  wire [9:0] _kouka_x_data_in179;
  wire [9:0] _kouka_x_data_in180;
  wire [9:0] _kouka_x_data_in181;
  wire [9:0] _kouka_x_data_in182;
  wire [9:0] _kouka_x_data_in183;
  wire [9:0] _kouka_x_data_in184;
  wire [9:0] _kouka_x_data_in185;
  wire [9:0] _kouka_x_data_in186;
  wire [9:0] _kouka_x_data_in187;
  wire [9:0] _kouka_x_data_in188;
  wire [9:0] _kouka_x_data_in189;
  wire [9:0] _kouka_x_data_in190;
  wire [9:0] _kouka_x_data_in193;
  wire [9:0] _kouka_x_data_in194;
  wire [9:0] _kouka_x_data_in195;
  wire [9:0] _kouka_x_data_in196;
  wire [9:0] _kouka_x_data_in197;
  wire [9:0] _kouka_x_data_in198;
  wire [9:0] _kouka_x_data_in199;
  wire [9:0] _kouka_x_data_in200;
  wire [9:0] _kouka_x_data_in201;
  wire [9:0] _kouka_x_data_in202;
  wire [9:0] _kouka_x_data_in203;
  wire [9:0] _kouka_x_data_in204;
  wire [9:0] _kouka_x_data_in205;
  wire [9:0] _kouka_x_data_in206;
  wire [9:0] _kouka_x_data_in207;
  wire [9:0] _kouka_x_data_in208;
  wire [9:0] _kouka_x_data_in209;
  wire [9:0] _kouka_x_data_in210;
  wire [9:0] _kouka_x_data_in211;
  wire [9:0] _kouka_x_data_in212;
  wire [9:0] _kouka_x_data_in213;
  wire [9:0] _kouka_x_data_in214;
  wire [9:0] _kouka_x_data_in215;
  wire [9:0] _kouka_x_data_in216;
  wire [9:0] _kouka_x_data_in217;
  wire [9:0] _kouka_x_data_in218;
  wire [9:0] _kouka_x_data_in219;
  wire [9:0] _kouka_x_data_in220;
  wire [9:0] _kouka_x_data_in221;
  wire [9:0] _kouka_x_data_in222;
  wire [9:0] _kouka_x_data_in225;
  wire [9:0] _kouka_x_data_in226;
  wire [9:0] _kouka_x_data_in227;
  wire [9:0] _kouka_x_data_in228;
  wire [9:0] _kouka_x_data_in229;
  wire [9:0] _kouka_x_data_in230;
  wire [9:0] _kouka_x_data_in231;
  wire [9:0] _kouka_x_data_in232;
  wire [9:0] _kouka_x_data_in233;
  wire [9:0] _kouka_x_data_in234;
  wire [9:0] _kouka_x_data_in235;
  wire [9:0] _kouka_x_data_in236;
  wire [9:0] _kouka_x_data_in237;
  wire [9:0] _kouka_x_data_in238;
  wire [9:0] _kouka_x_data_in239;
  wire [9:0] _kouka_x_data_in240;
  wire [9:0] _kouka_x_data_in241;
  wire [9:0] _kouka_x_data_in242;
  wire [9:0] _kouka_x_data_in243;
  wire [9:0] _kouka_x_data_in244;
  wire [9:0] _kouka_x_data_in245;
  wire [9:0] _kouka_x_data_in246;
  wire [9:0] _kouka_x_data_in247;
  wire [9:0] _kouka_x_data_in248;
  wire [9:0] _kouka_x_data_in249;
  wire [9:0] _kouka_x_data_in250;
  wire [9:0] _kouka_x_data_in251;
  wire [9:0] _kouka_x_data_in252;
  wire [9:0] _kouka_x_data_in253;
  wire [9:0] _kouka_x_data_in254;
  wire [9:0] _kouka_x_data_in257;
  wire [9:0] _kouka_x_data_in258;
  wire [9:0] _kouka_x_data_in259;
  wire [9:0] _kouka_x_data_in260;
  wire [9:0] _kouka_x_data_in261;
  wire [9:0] _kouka_x_data_in262;
  wire [9:0] _kouka_x_data_in263;
  wire [9:0] _kouka_x_data_in264;
  wire [9:0] _kouka_x_data_in265;
  wire [9:0] _kouka_x_data_in266;
  wire [9:0] _kouka_x_data_in267;
  wire [9:0] _kouka_x_data_in268;
  wire [9:0] _kouka_x_data_in269;
  wire [9:0] _kouka_x_data_in270;
  wire [9:0] _kouka_x_data_in271;
  wire [9:0] _kouka_x_data_in272;
  wire [9:0] _kouka_x_data_in273;
  wire [9:0] _kouka_x_data_in274;
  wire [9:0] _kouka_x_data_in275;
  wire [9:0] _kouka_x_data_in276;
  wire [9:0] _kouka_x_data_in277;
  wire [9:0] _kouka_x_data_in278;
  wire [9:0] _kouka_x_data_in279;
  wire [9:0] _kouka_x_data_in280;
  wire [9:0] _kouka_x_data_in281;
  wire [9:0] _kouka_x_data_in282;
  wire [9:0] _kouka_x_data_in283;
  wire [9:0] _kouka_x_data_in284;
  wire [9:0] _kouka_x_data_in285;
  wire [9:0] _kouka_x_data_in286;
  wire [9:0] _kouka_x_data_in289;
  wire [9:0] _kouka_x_data_in290;
  wire [9:0] _kouka_x_data_in291;
  wire [9:0] _kouka_x_data_in292;
  wire [9:0] _kouka_x_data_in293;
  wire [9:0] _kouka_x_data_in294;
  wire [9:0] _kouka_x_data_in295;
  wire [9:0] _kouka_x_data_in296;
  wire [9:0] _kouka_x_data_in297;
  wire [9:0] _kouka_x_data_in298;
  wire [9:0] _kouka_x_data_in299;
  wire [9:0] _kouka_x_data_in300;
  wire [9:0] _kouka_x_data_in301;
  wire [9:0] _kouka_x_data_in302;
  wire [9:0] _kouka_x_data_in303;
  wire [9:0] _kouka_x_data_in304;
  wire [9:0] _kouka_x_data_in305;
  wire [9:0] _kouka_x_data_in306;
  wire [9:0] _kouka_x_data_in307;
  wire [9:0] _kouka_x_data_in308;
  wire [9:0] _kouka_x_data_in309;
  wire [9:0] _kouka_x_data_in310;
  wire [9:0] _kouka_x_data_in311;
  wire [9:0] _kouka_x_data_in312;
  wire [9:0] _kouka_x_data_in313;
  wire [9:0] _kouka_x_data_in314;
  wire [9:0] _kouka_x_data_in315;
  wire [9:0] _kouka_x_data_in316;
  wire [9:0] _kouka_x_data_in317;
  wire [9:0] _kouka_x_data_in318;
  wire [9:0] _kouka_x_data_in321;
  wire [9:0] _kouka_x_data_in322;
  wire [9:0] _kouka_x_data_in323;
  wire [9:0] _kouka_x_data_in324;
  wire [9:0] _kouka_x_data_in325;
  wire [9:0] _kouka_x_data_in326;
  wire [9:0] _kouka_x_data_in327;
  wire [9:0] _kouka_x_data_in328;
  wire [9:0] _kouka_x_data_in329;
  wire [9:0] _kouka_x_data_in330;
  wire [9:0] _kouka_x_data_in331;
  wire [9:0] _kouka_x_data_in332;
  wire [9:0] _kouka_x_data_in333;
  wire [9:0] _kouka_x_data_in334;
  wire [9:0] _kouka_x_data_in335;
  wire [9:0] _kouka_x_data_in336;
  wire [9:0] _kouka_x_data_in337;
  wire [9:0] _kouka_x_data_in338;
  wire [9:0] _kouka_x_data_in339;
  wire [9:0] _kouka_x_data_in340;
  wire [9:0] _kouka_x_data_in341;
  wire [9:0] _kouka_x_data_in342;
  wire [9:0] _kouka_x_data_in343;
  wire [9:0] _kouka_x_data_in344;
  wire [9:0] _kouka_x_data_in345;
  wire [9:0] _kouka_x_data_in346;
  wire [9:0] _kouka_x_data_in347;
  wire [9:0] _kouka_x_data_in348;
  wire [9:0] _kouka_x_data_in349;
  wire [9:0] _kouka_x_data_in350;
  wire [9:0] _kouka_x_data_in353;
  wire [9:0] _kouka_x_data_in354;
  wire [9:0] _kouka_x_data_in355;
  wire [9:0] _kouka_x_data_in356;
  wire [9:0] _kouka_x_data_in357;
  wire [9:0] _kouka_x_data_in358;
  wire [9:0] _kouka_x_data_in359;
  wire [9:0] _kouka_x_data_in360;
  wire [9:0] _kouka_x_data_in361;
  wire [9:0] _kouka_x_data_in362;
  wire [9:0] _kouka_x_data_in363;
  wire [9:0] _kouka_x_data_in364;
  wire [9:0] _kouka_x_data_in365;
  wire [9:0] _kouka_x_data_in366;
  wire [9:0] _kouka_x_data_in367;
  wire [9:0] _kouka_x_data_in368;
  wire [9:0] _kouka_x_data_in369;
  wire [9:0] _kouka_x_data_in370;
  wire [9:0] _kouka_x_data_in371;
  wire [9:0] _kouka_x_data_in372;
  wire [9:0] _kouka_x_data_in373;
  wire [9:0] _kouka_x_data_in374;
  wire [9:0] _kouka_x_data_in375;
  wire [9:0] _kouka_x_data_in376;
  wire [9:0] _kouka_x_data_in377;
  wire [9:0] _kouka_x_data_in378;
  wire [9:0] _kouka_x_data_in379;
  wire [9:0] _kouka_x_data_in380;
  wire [9:0] _kouka_x_data_in381;
  wire [9:0] _kouka_x_data_in382;
  wire [9:0] _kouka_x_data_in385;
  wire [9:0] _kouka_x_data_in386;
  wire [9:0] _kouka_x_data_in387;
  wire [9:0] _kouka_x_data_in388;
  wire [9:0] _kouka_x_data_in389;
  wire [9:0] _kouka_x_data_in390;
  wire [9:0] _kouka_x_data_in391;
  wire [9:0] _kouka_x_data_in392;
  wire [9:0] _kouka_x_data_in393;
  wire [9:0] _kouka_x_data_in394;
  wire [9:0] _kouka_x_data_in395;
  wire [9:0] _kouka_x_data_in396;
  wire [9:0] _kouka_x_data_in397;
  wire [9:0] _kouka_x_data_in398;
  wire [9:0] _kouka_x_data_in399;
  wire [9:0] _kouka_x_data_in400;
  wire [9:0] _kouka_x_data_in401;
  wire [9:0] _kouka_x_data_in402;
  wire [9:0] _kouka_x_data_in403;
  wire [9:0] _kouka_x_data_in404;
  wire [9:0] _kouka_x_data_in405;
  wire [9:0] _kouka_x_data_in406;
  wire [9:0] _kouka_x_data_in407;
  wire [9:0] _kouka_x_data_in408;
  wire [9:0] _kouka_x_data_in409;
  wire [9:0] _kouka_x_data_in410;
  wire [9:0] _kouka_x_data_in411;
  wire [9:0] _kouka_x_data_in412;
  wire [9:0] _kouka_x_data_in413;
  wire [9:0] _kouka_x_data_in414;
  wire [9:0] _kouka_x_data_in417;
  wire [9:0] _kouka_x_data_in418;
  wire [9:0] _kouka_x_data_in419;
  wire [9:0] _kouka_x_data_in420;
  wire [9:0] _kouka_x_data_in421;
  wire [9:0] _kouka_x_data_in422;
  wire [9:0] _kouka_x_data_in423;
  wire [9:0] _kouka_x_data_in424;
  wire [9:0] _kouka_x_data_in425;
  wire [9:0] _kouka_x_data_in426;
  wire [9:0] _kouka_x_data_in427;
  wire [9:0] _kouka_x_data_in428;
  wire [9:0] _kouka_x_data_in429;
  wire [9:0] _kouka_x_data_in430;
  wire [9:0] _kouka_x_data_in431;
  wire [9:0] _kouka_x_data_in432;
  wire [9:0] _kouka_x_data_in433;
  wire [9:0] _kouka_x_data_in434;
  wire [9:0] _kouka_x_data_in435;
  wire [9:0] _kouka_x_data_in436;
  wire [9:0] _kouka_x_data_in437;
  wire [9:0] _kouka_x_data_in438;
  wire [9:0] _kouka_x_data_in439;
  wire [9:0] _kouka_x_data_in440;
  wire [9:0] _kouka_x_data_in441;
  wire [9:0] _kouka_x_data_in442;
  wire [9:0] _kouka_x_data_in443;
  wire [9:0] _kouka_x_data_in444;
  wire [9:0] _kouka_x_data_in445;
  wire [9:0] _kouka_x_data_in446;
  wire [9:0] _kouka_x_data_in449;
  wire [9:0] _kouka_x_data_in450;
  wire [9:0] _kouka_x_data_in451;
  wire [9:0] _kouka_x_data_in452;
  wire [9:0] _kouka_x_data_in453;
  wire [9:0] _kouka_x_data_in454;
  wire [9:0] _kouka_x_data_in455;
  wire [9:0] _kouka_x_data_in456;
  wire [9:0] _kouka_x_data_in457;
  wire [9:0] _kouka_x_data_in458;
  wire [9:0] _kouka_x_data_in459;
  wire [9:0] _kouka_x_data_in460;
  wire [9:0] _kouka_x_data_in461;
  wire [9:0] _kouka_x_data_in462;
  wire [9:0] _kouka_x_data_in463;
  wire [9:0] _kouka_x_data_in464;
  wire [9:0] _kouka_x_data_in465;
  wire [9:0] _kouka_x_data_in466;
  wire [9:0] _kouka_x_data_in467;
  wire [9:0] _kouka_x_data_in468;
  wire [9:0] _kouka_x_data_in469;
  wire [9:0] _kouka_x_data_in470;
  wire [9:0] _kouka_x_data_in471;
  wire [9:0] _kouka_x_data_in472;
  wire [9:0] _kouka_x_data_in473;
  wire [9:0] _kouka_x_data_in474;
  wire [9:0] _kouka_x_data_in475;
  wire [9:0] _kouka_x_data_in476;
  wire [9:0] _kouka_x_data_in477;
  wire [9:0] _kouka_x_data_in478;
  wire [9:0] _kouka_x_start;
  wire [9:0] _kouka_x_goal;
  wire [9:0] _kouka_x_loot_out0;
  wire [9:0] _kouka_x_loot_out1;
  wire [9:0] _kouka_x_loot_out2;
  wire [9:0] _kouka_x_loot_out3;
  wire [9:0] _kouka_x_loot_out4;
  wire [9:0] _kouka_x_loot_out5;
  wire [9:0] _kouka_x_loot_out6;
  wire [9:0] _kouka_x_loot_out7;
  wire [9:0] _kouka_x_loot_out8;
  wire [9:0] _kouka_x_loot_out9;
  wire [9:0] _kouka_x_loot_out10;
  wire [9:0] _kouka_x_loot_out11;
  wire [9:0] _kouka_x_loot_out12;
  wire [9:0] _kouka_x_loot_out13;
  wire [9:0] _kouka_x_loot_out14;
  wire [9:0] _kouka_x_loot_out15;
  wire [9:0] _kouka_x_loot_out16;
  wire [9:0] _kouka_x_loot_out17;
  wire [9:0] _kouka_x_loot_out18;
  wire [9:0] _kouka_x_loot_out19;
  wire [9:0] _kouka_x_loot_out20;
  wire [9:0] _kouka_x_loot_out21;
  wire [9:0] _kouka_x_loot_out22;
  wire [9:0] _kouka_x_loot_out23;
  wire [9:0] _kouka_x_loot_out24;
  wire [9:0] _kouka_x_loot_out25;
  wire [9:0] _kouka_x_loot_out26;
  wire [9:0] _kouka_x_loot_out27;
  wire [9:0] _kouka_x_loot_out28;
  wire [9:0] _kouka_x_loot_out29;
  wire [9:0] _kouka_x_loot_out30;
  wire [9:0] _kouka_x_loot_out31;
  wire [9:0] _kouka_x_loot_out32;
  wire [9:0] _kouka_x_loot_out33;
  wire [9:0] _kouka_x_loot_out34;
  wire [9:0] _kouka_x_loot_out35;
  wire [9:0] _kouka_x_loot_out36;
  wire [9:0] _kouka_x_loot_out37;
  wire [9:0] _kouka_x_loot_out38;
  wire [9:0] _kouka_x_loot_out39;
  wire [9:0] _kouka_x_loot_out40;
  wire [9:0] _kouka_x_loot_out41;
  wire [9:0] _kouka_x_loot_out42;
  wire [9:0] _kouka_x_loot_out43;
  wire [9:0] _kouka_x_loot_out44;
  wire [9:0] _kouka_x_loot_out45;
  wire [9:0] _kouka_x_loot_out46;
  wire [9:0] _kouka_x_loot_out47;
  wire [9:0] _kouka_x_loot_out48;
  wire [9:0] _kouka_x_loot_out49;
  wire [9:0] _kouka_x_loot_out50;
  wire [9:0] _kouka_x_loot_out51;
  wire [9:0] _kouka_x_loot_out52;
  wire [9:0] _kouka_x_loot_out53;
  wire [9:0] _kouka_x_loot_out54;
  wire [9:0] _kouka_x_loot_out55;
  wire [9:0] _kouka_x_loot_out56;
  wire [9:0] _kouka_x_loot_out57;
  wire [9:0] _kouka_x_loot_out58;
  wire [9:0] _kouka_x_loot_out59;
  wire [9:0] _kouka_x_loot_out60;
  wire [9:0] _kouka_x_loot_out61;
  wire [9:0] _kouka_x_loot_out62;
  wire [9:0] _kouka_x_loot_out63;
  wire [9:0] _kouka_x_loot_out64;
  wire [9:0] _kouka_x_loot_out65;
  wire [9:0] _kouka_x_loot_out66;
  wire [9:0] _kouka_x_loot_out67;
  wire [9:0] _kouka_x_loot_out68;
  wire [9:0] _kouka_x_loot_out69;
  wire [9:0] _kouka_x_loot_out70;
  wire [9:0] _kouka_x_loot_out71;
  wire [9:0] _kouka_x_loot_out72;
  wire [9:0] _kouka_x_loot_out73;
  wire [9:0] _kouka_x_loot_out74;
  wire [9:0] _kouka_x_loot_out75;
  wire [9:0] _kouka_x_loot_out76;
  wire [9:0] _kouka_x_loot_out77;
  wire [9:0] _kouka_x_loot_out78;
  wire [9:0] _kouka_x_loot_out79;
  wire [9:0] _kouka_x_loot_out80;
  wire [9:0] _kouka_x_loot_out81;
  wire [9:0] _kouka_x_loot_out82;
  wire [9:0] _kouka_x_loot_out83;
  wire [9:0] _kouka_x_loot_out84;
  wire [9:0] _kouka_x_loot_out85;
  wire [9:0] _kouka_x_loot_out86;
  wire [9:0] _kouka_x_loot_out87;
  wire [9:0] _kouka_x_loot_out88;
  wire [9:0] _kouka_x_loot_out89;
  wire [9:0] _kouka_x_loot_out90;
  wire [9:0] _kouka_x_loot_out91;
  wire [9:0] _kouka_x_loot_out92;
  wire [9:0] _kouka_x_loot_out93;
  wire [9:0] _kouka_x_loot_out94;
  wire [9:0] _kouka_x_loot_out95;
  wire [9:0] _kouka_x_loot_out96;
  wire [9:0] _kouka_x_loot_out97;
  wire [9:0] _kouka_x_loot_out98;
  wire [9:0] _kouka_x_loot_out99;
  wire [9:0] _kouka_x_loot_out100;
  wire [9:0] _kouka_x_loot_out101;
  wire [9:0] _kouka_x_loot_out102;
  wire [9:0] _kouka_x_loot_out103;
  wire [9:0] _kouka_x_loot_out104;
  wire [9:0] _kouka_x_loot_out105;
  wire [9:0] _kouka_x_loot_out106;
  wire [9:0] _kouka_x_loot_out107;
  wire [9:0] _kouka_x_loot_out108;
  wire [9:0] _kouka_x_loot_out109;
  wire [9:0] _kouka_x_loot_out110;
  wire [9:0] _kouka_x_loot_out111;
  wire [9:0] _kouka_x_loot_out112;
  wire [9:0] _kouka_x_loot_out113;
  wire [9:0] _kouka_x_loot_out114;
  wire [9:0] _kouka_x_loot_out115;
  wire [9:0] _kouka_x_loot_out116;
  wire [9:0] _kouka_x_loot_out117;
  wire [9:0] _kouka_x_loot_out118;
  wire [9:0] _kouka_x_loot_out119;
  wire [9:0] _kouka_x_loot_out120;
  wire [9:0] _kouka_x_loot_out121;
  wire [9:0] _kouka_x_loot_out122;
  wire [9:0] _kouka_x_loot_out123;
  wire [9:0] _kouka_x_loot_out124;
  wire [9:0] _kouka_x_loot_out125;
  wire [9:0] _kouka_x_loot_out126;
  wire [9:0] _kouka_x_loot_out127;
  wire [9:0] _kouka_x_loot_out128;
  wire [9:0] _kouka_x_loot_out129;
  wire [9:0] _kouka_x_loot_out130;
  wire [9:0] _kouka_x_loot_out131;
  wire [9:0] _kouka_x_loot_out132;
  wire [9:0] _kouka_x_loot_out133;
  wire [9:0] _kouka_x_loot_out134;
  wire [9:0] _kouka_x_loot_out135;
  wire [9:0] _kouka_x_loot_out136;
  wire [9:0] _kouka_x_loot_out137;
  wire [9:0] _kouka_x_loot_out138;
  wire [9:0] _kouka_x_loot_out139;
  wire [9:0] _kouka_x_loot_out140;
  wire [9:0] _kouka_x_loot_out141;
  wire [9:0] _kouka_x_loot_out142;
  wire [9:0] _kouka_x_loot_out143;
  wire [9:0] _kouka_x_loot_out144;
  wire [9:0] _kouka_x_loot_out145;
  wire [9:0] _kouka_x_loot_out146;
  wire [9:0] _kouka_x_loot_out147;
  wire [9:0] _kouka_x_loot_out148;
  wire [9:0] _kouka_x_loot_out149;
  wire [9:0] _kouka_x_loot_out150;
  wire [9:0] _kouka_x_loot_out151;
  wire [9:0] _kouka_x_loot_out152;
  wire [9:0] _kouka_x_loot_out153;
  wire [9:0] _kouka_x_loot_out154;
  wire [9:0] _kouka_x_loot_out155;
  wire [9:0] _kouka_x_loot_out156;
  wire [9:0] _kouka_x_loot_out157;
  wire [9:0] _kouka_x_loot_out158;
  wire [9:0] _kouka_x_loot_out159;
  wire [9:0] _kouka_x_loot_out160;
  wire [9:0] _kouka_x_loot_out161;
  wire [9:0] _kouka_x_loot_out162;
  wire [9:0] _kouka_x_loot_out163;
  wire [9:0] _kouka_x_loot_out164;
  wire [9:0] _kouka_x_loot_out165;
  wire [9:0] _kouka_x_loot_out166;
  wire [9:0] _kouka_x_loot_out167;
  wire [9:0] _kouka_x_loot_out168;
  wire [9:0] _kouka_x_loot_out169;
  wire [9:0] _kouka_x_loot_out170;
  wire [9:0] _kouka_x_loot_out171;
  wire [9:0] _kouka_x_loot_out172;
  wire [9:0] _kouka_x_loot_out173;
  wire [9:0] _kouka_x_loot_out174;
  wire [9:0] _kouka_x_loot_out175;
  wire [9:0] _kouka_x_loot_out176;
  wire [9:0] _kouka_x_loot_out177;
  wire [9:0] _kouka_x_loot_out178;
  wire [9:0] _kouka_x_loot_out179;
  wire [9:0] _kouka_x_loot_out180;
  wire [9:0] _kouka_x_loot_out181;
  wire [9:0] _kouka_x_loot_out182;
  wire [9:0] _kouka_x_loot_out183;
  wire [9:0] _kouka_x_loot_out184;
  wire [9:0] _kouka_x_loot_out185;
  wire [9:0] _kouka_x_loot_out186;
  wire [9:0] _kouka_x_loot_out187;
  wire [9:0] _kouka_x_loot_out188;
  wire [9:0] _kouka_x_loot_out189;
  wire [9:0] _kouka_x_loot_out190;
  wire [9:0] _kouka_x_loot_out191;
  wire [9:0] _kouka_x_loot_out192;
  wire [9:0] _kouka_x_loot_out193;
  wire [9:0] _kouka_x_loot_out194;
  wire [9:0] _kouka_x_loot_out195;
  wire [9:0] _kouka_x_loot_out196;
  wire [9:0] _kouka_x_loot_out197;
  wire [9:0] _kouka_x_loot_out198;
  wire [9:0] _kouka_x_loot_out199;
  wire [9:0] _kouka_x_loot_out200;
  wire [9:0] _kouka_x_loot_out201;
  wire [9:0] _kouka_x_loot_out202;
  wire [9:0] _kouka_x_loot_out203;
  wire [9:0] _kouka_x_loot_out204;
  wire [9:0] _kouka_x_loot_out205;
  wire [9:0] _kouka_x_loot_out206;
  wire [9:0] _kouka_x_loot_out207;
  wire [9:0] _kouka_x_loot_out208;
  wire [9:0] _kouka_x_loot_out209;
  wire [9:0] _kouka_x_loot_out210;
  wire [9:0] _kouka_x_loot_out211;
  wire [9:0] _kouka_x_loot_out212;
  wire [9:0] _kouka_x_loot_out213;
  wire [9:0] _kouka_x_loot_out214;
  wire [9:0] _kouka_x_loot_out215;
  wire [9:0] _kouka_x_loot_out216;
  wire [9:0] _kouka_x_loot_out217;
  wire [9:0] _kouka_x_loot_out218;
  wire [9:0] _kouka_x_loot_out219;
  wire [9:0] _kouka_x_loot_out220;
  wire [9:0] _kouka_x_loot_out221;
  wire [9:0] _kouka_x_loot_out222;
  wire _kouka_x_in_do;
  wire _kouka_x_out_do;
  wire _kouka_x_p_reset;
  wire _kouka_x_m_clock;
  reg _reg_0;
  wire _net_1;
  wire _net_2;
  wire _net_3;
  wire _net_4;
  wire _net_5;
  wire _net_6;
  wire _net_7;
  wire _net_8;
  wire _net_9;
  wire _net_10;
  wire _net_11;
  wire _net_12;
  wire _net_13;
  wire _net_14;
  wire _net_15;
  wire _net_16;
  wire _net_17;
  wire _net_18;
  wire _net_19;
  wire _net_20;
  wire _net_21;
  wire _net_22;
  wire _net_23;
  wire _net_24;
  wire _net_25;
  wire _net_26;
  wire _net_27;
  wire _net_28;
  wire _net_29;
  wire _net_30;
  wire _net_31;
  wire _net_32;
  wire _net_33;
  wire _net_34;
  wire _net_35;
  wire _net_36;
  wire _net_37;
  wire _net_38;
  wire _net_39;
  wire _net_40;
  wire _net_41;
  wire _net_42;
  wire _net_43;
  wire _net_44;
  wire _net_45;
  wire _net_46;
  wire _net_47;
  wire _net_48;
  wire _net_49;
  wire _net_50;
  wire _net_51;
  wire _net_52;
  wire _net_53;
  wire _net_54;
  wire _net_55;
  wire _net_56;
  wire _net_57;
  wire _net_58;
  wire _net_59;
  wire _net_60;
  wire _net_61;
  wire _net_62;
  wire _net_63;
  wire _net_64;
  wire _net_65;
  wire _net_66;
  wire _net_67;
  wire _net_68;
  wire _net_69;
  wire _net_70;
  wire _net_71;
  wire _net_72;
  wire _net_73;
  wire _net_74;
  wire _net_75;
  wire _net_76;
  wire _net_77;
  wire _net_78;
  wire _net_79;
  wire _net_80;
  wire _net_81;
  wire _net_82;
  wire _net_83;
  wire _net_84;
  wire _net_85;
  wire _net_86;
  wire _net_87;
  wire _net_88;
  wire _net_89;
  wire _net_90;
  wire _net_91;
  wire _net_92;
  wire _net_93;
  wire _net_94;
  wire _net_95;
  wire _net_96;
  wire _net_97;
  wire _net_98;
  wire _net_99;
  wire _net_100;
  wire _net_101;
  wire _net_102;
  wire _net_103;
  wire _net_104;
  wire _net_105;
  wire _net_106;
  wire _net_107;
  wire _net_108;
  wire _net_109;
  wire _net_110;
  wire _net_111;
  wire _net_112;
  wire _net_113;
  wire _net_114;
  wire _net_115;
  wire _net_116;
  wire _net_117;
  wire _net_118;
  wire _net_119;
  wire _net_120;
  wire _net_121;
  wire _net_122;
  wire _net_123;
  wire _net_124;
  wire _net_125;
  wire _net_126;
  wire _net_127;
  wire _net_128;
  wire _net_129;
  wire _net_130;
  wire _net_131;
  wire _net_132;
  wire _net_133;
  wire _net_134;
  wire _net_135;
  wire _net_136;
  wire _net_137;
  wire _net_138;
  wire _net_139;
  wire _net_140;
  wire _net_141;
  wire _net_142;
  wire _net_143;
  wire _net_144;
  wire _net_145;
  wire _net_146;
  wire _net_147;
  wire _net_148;
  wire _net_149;
  wire _net_150;
  wire _net_151;
  wire _net_152;
  wire _net_153;
  wire _net_154;
  wire _net_155;
  wire _net_156;
  wire _net_157;
  wire _net_158;
  wire _net_159;
  wire _net_160;
  wire _net_161;
  wire _net_162;
  wire _net_163;
  wire _net_164;
  wire _net_165;
  wire _net_166;
  wire _net_167;
  wire _net_168;
  wire _net_169;
  wire _net_170;
  wire _net_171;
  wire _net_172;
  wire _net_173;
  wire _net_174;
  wire _net_175;
  wire _net_176;
  wire _net_177;
  wire _net_178;
  wire _net_179;
  wire _net_180;
  wire _net_181;
  wire _net_182;
  wire _net_183;
  wire _net_184;
  wire _net_185;
  wire _net_186;
  wire _net_187;
  wire _net_188;
  wire _net_189;
  wire _net_190;
  wire _net_191;
  wire _net_192;
  wire _net_193;
  wire _net_194;
  wire _net_195;
  wire _net_196;
  wire _net_197;
  wire _net_198;
  wire _net_199;
  wire _net_200;
  wire _net_201;
  wire _net_202;
  wire _net_203;
  wire _net_204;
  wire _net_205;
  wire _net_206;
  wire _net_207;
  wire _net_208;
  wire _net_209;
  wire _net_210;
  wire _net_211;
  wire _net_212;
  wire _net_213;
  wire _net_214;
  wire _net_215;
  wire _net_216;
  wire _net_217;
  wire _net_218;
  wire _net_219;
  wire _net_220;
  wire _net_221;
  wire _net_222;
  wire _net_223;
  wire _net_224;
  wire _net_225;
  wire _net_226;
  wire _net_227;
  wire _net_228;
  wire _net_229;
  wire _net_230;
  wire _net_231;
  wire _net_232;
  wire _net_233;
  wire _net_234;
  wire _net_235;
  wire _net_236;
  wire _net_237;
  wire _net_238;
  wire _net_239;
  wire _net_240;
  wire _net_241;
  wire _net_242;
  wire _net_243;
  wire _net_244;
  wire _net_245;
  wire _net_246;
  wire _net_247;
  wire _net_248;
  wire _net_249;
  wire _net_250;
  wire _net_251;
  wire _net_252;
  wire _net_253;
  wire _net_254;
  wire _net_255;
  wire _net_256;
  wire _net_257;
  wire _net_258;
  wire _net_259;
  wire _net_260;
  wire _net_261;
  wire _net_262;
  wire _net_263;
  wire _net_264;
  wire _net_265;
  wire _net_266;
  wire _net_267;
  wire _net_268;
  wire _net_269;
  wire _net_270;
  wire _net_271;
  wire _net_272;
  wire _net_273;
  wire _net_274;
  wire _net_275;
  wire _net_276;
  wire _net_277;
  wire _net_278;
  wire _net_279;
  wire _net_280;
  wire _net_281;
  wire _net_282;
  wire _net_283;
  wire _net_284;
  wire _net_285;
  wire _net_286;
  wire _net_287;
  wire _net_288;
  wire _net_289;
  wire _net_290;
  wire _net_291;
  wire _net_292;
  wire _net_293;
  wire _net_294;
  wire _net_295;
  wire _net_296;
  wire _net_297;
  wire _net_298;
  wire _net_299;
  wire _net_300;
  wire _net_301;
  wire _net_302;
  wire _net_303;
  wire _net_304;
  wire _net_305;
  wire _net_306;
  wire _net_307;
  wire _net_308;
  wire _net_309;
  wire _net_310;
  wire _net_311;
  wire _net_312;
  wire _net_313;
  wire _net_314;
  wire _net_315;
  wire _net_316;
  wire _net_317;
  wire _net_318;
  wire _net_319;
  wire _net_320;
  wire _net_321;
  wire _net_322;
  wire _net_323;
  wire _net_324;
  wire _net_325;
  wire _net_326;
  wire _net_327;
  wire _net_328;
  wire _net_329;
  wire _net_330;
  wire _net_331;
  wire _net_332;
  wire _net_333;
  wire _net_334;
  wire _net_335;
  wire _net_336;
  wire _net_337;
  wire _net_338;
  wire _net_339;
  wire _net_340;
  wire _net_341;
  wire _net_342;
  wire _net_343;
  wire _net_344;
  wire _net_345;
  wire _net_346;
  wire _net_347;
  wire _net_348;
  wire _net_349;
  wire _net_350;
  wire _net_351;
  wire _net_352;
  wire _net_353;
  wire _net_354;
  wire _net_355;
  wire _net_356;
  wire _net_357;
  wire _net_358;
  wire _net_359;
  wire _net_360;
  wire _net_361;
  wire _net_362;
  wire _net_363;
  wire _net_364;
  wire _net_365;
  wire _net_366;
  wire _net_367;
  wire _net_368;
  wire _net_369;
  wire _net_370;
  wire _net_371;
  wire _net_372;
  wire _net_373;
  wire _net_374;
  wire _net_375;
  wire _net_376;
  wire _net_377;
  wire _net_378;
  wire _net_379;
  wire _net_380;
  wire _net_381;
  wire _net_382;
  wire _net_383;
  wire _net_384;
  wire _net_385;
  wire _net_386;
  wire _net_387;
  wire _net_388;
  wire _net_389;
  wire _net_390;
  wire _net_391;
  wire _net_392;
  wire _net_393;
  wire _net_394;
  wire _net_395;
  wire _net_396;
  wire _net_397;
  wire _net_398;
  wire _net_399;
  wire _net_400;
  wire _net_401;
  wire _net_402;
  wire _net_403;
  wire _net_404;
  wire _net_405;
  wire _net_406;
  wire _net_407;
  wire _net_408;
  wire _net_409;
  wire _net_410;
  wire _net_411;
  wire _net_412;
  wire _net_413;
  wire _net_414;
  wire _net_415;
  wire _net_416;
  wire _net_417;
  wire _net_418;
  wire _net_419;
  wire _net_420;
  wire _net_421;
kouka kouka_x (.m_clock(m_clock), .p_reset( p_reset), .out_do(_kouka_x_out_do), .in_do(_kouka_x_in_do), .loot_out0(_kouka_x_loot_out0), .loot_out1(_kouka_x_loot_out1), .loot_out2(_kouka_x_loot_out2), .loot_out3(_kouka_x_loot_out3), .loot_out4(_kouka_x_loot_out4), .loot_out5(_kouka_x_loot_out5), .loot_out6(_kouka_x_loot_out6), .loot_out7(_kouka_x_loot_out7), .loot_out8(_kouka_x_loot_out8), .loot_out9(_kouka_x_loot_out9), .loot_out10(_kouka_x_loot_out10), .loot_out11(_kouka_x_loot_out11), .loot_out12(_kouka_x_loot_out12), .loot_out13(_kouka_x_loot_out13), .loot_out14(_kouka_x_loot_out14), .loot_out15(_kouka_x_loot_out15), .loot_out16(_kouka_x_loot_out16), .loot_out17(_kouka_x_loot_out17), .loot_out18(_kouka_x_loot_out18), .loot_out19(_kouka_x_loot_out19), .loot_out20(_kouka_x_loot_out20), .loot_out21(_kouka_x_loot_out21), .loot_out22(_kouka_x_loot_out22), .loot_out23(_kouka_x_loot_out23), .loot_out24(_kouka_x_loot_out24), .loot_out25(_kouka_x_loot_out25), .loot_out26(_kouka_x_loot_out26), .loot_out27(_kouka_x_loot_out27), .loot_out28(_kouka_x_loot_out28), .loot_out29(_kouka_x_loot_out29), .loot_out30(_kouka_x_loot_out30), .loot_out31(_kouka_x_loot_out31), .loot_out32(_kouka_x_loot_out32), .loot_out33(_kouka_x_loot_out33), .loot_out34(_kouka_x_loot_out34), .loot_out35(_kouka_x_loot_out35), .loot_out36(_kouka_x_loot_out36), .loot_out37(_kouka_x_loot_out37), .loot_out38(_kouka_x_loot_out38), .loot_out39(_kouka_x_loot_out39), .loot_out40(_kouka_x_loot_out40), .loot_out41(_kouka_x_loot_out41), .loot_out42(_kouka_x_loot_out42), .loot_out43(_kouka_x_loot_out43), .loot_out44(_kouka_x_loot_out44), .loot_out45(_kouka_x_loot_out45), .loot_out46(_kouka_x_loot_out46), .loot_out47(_kouka_x_loot_out47), .loot_out48(_kouka_x_loot_out48), .loot_out49(_kouka_x_loot_out49), .loot_out50(_kouka_x_loot_out50), .loot_out51(_kouka_x_loot_out51), .loot_out52(_kouka_x_loot_out52), .loot_out53(_kouka_x_loot_out53), .loot_out54(_kouka_x_loot_out54), .loot_out55(_kouka_x_loot_out55), .loot_out56(_kouka_x_loot_out56), .loot_out57(_kouka_x_loot_out57), .loot_out58(_kouka_x_loot_out58), .loot_out59(_kouka_x_loot_out59), .loot_out60(_kouka_x_loot_out60), .loot_out61(_kouka_x_loot_out61), .loot_out62(_kouka_x_loot_out62), .loot_out63(_kouka_x_loot_out63), .loot_out64(_kouka_x_loot_out64), .loot_out65(_kouka_x_loot_out65), .loot_out66(_kouka_x_loot_out66), .loot_out67(_kouka_x_loot_out67), .loot_out68(_kouka_x_loot_out68), .loot_out69(_kouka_x_loot_out69), .loot_out70(_kouka_x_loot_out70), .loot_out71(_kouka_x_loot_out71), .loot_out72(_kouka_x_loot_out72), .loot_out73(_kouka_x_loot_out73), .loot_out74(_kouka_x_loot_out74), .loot_out75(_kouka_x_loot_out75), .loot_out76(_kouka_x_loot_out76), .loot_out77(_kouka_x_loot_out77), .loot_out78(_kouka_x_loot_out78), .loot_out79(_kouka_x_loot_out79), .loot_out80(_kouka_x_loot_out80), .loot_out81(_kouka_x_loot_out81), .loot_out82(_kouka_x_loot_out82), .loot_out83(_kouka_x_loot_out83), .loot_out84(_kouka_x_loot_out84), .loot_out85(_kouka_x_loot_out85), .loot_out86(_kouka_x_loot_out86), .loot_out87(_kouka_x_loot_out87), .loot_out88(_kouka_x_loot_out88), .loot_out89(_kouka_x_loot_out89), .loot_out90(_kouka_x_loot_out90), .loot_out91(_kouka_x_loot_out91), .loot_out92(_kouka_x_loot_out92), .loot_out93(_kouka_x_loot_out93), .loot_out94(_kouka_x_loot_out94), .loot_out95(_kouka_x_loot_out95), .loot_out96(_kouka_x_loot_out96), .loot_out97(_kouka_x_loot_out97), .loot_out98(_kouka_x_loot_out98), .loot_out99(_kouka_x_loot_out99), .loot_out100(_kouka_x_loot_out100), .loot_out101(_kouka_x_loot_out101), .loot_out102(_kouka_x_loot_out102), .loot_out103(_kouka_x_loot_out103), .loot_out104(_kouka_x_loot_out104), .loot_out105(_kouka_x_loot_out105), .loot_out106(_kouka_x_loot_out106), .loot_out107(_kouka_x_loot_out107), .loot_out108(_kouka_x_loot_out108), .loot_out109(_kouka_x_loot_out109), .loot_out110(_kouka_x_loot_out110), .loot_out111(_kouka_x_loot_out111), .loot_out112(_kouka_x_loot_out112), .loot_out113(_kouka_x_loot_out113), .loot_out114(_kouka_x_loot_out114), .loot_out115(_kouka_x_loot_out115), .loot_out116(_kouka_x_loot_out116), .loot_out117(_kouka_x_loot_out117), .loot_out118(_kouka_x_loot_out118), .loot_out119(_kouka_x_loot_out119), .loot_out120(_kouka_x_loot_out120), .loot_out121(_kouka_x_loot_out121), .loot_out122(_kouka_x_loot_out122), .loot_out123(_kouka_x_loot_out123), .loot_out124(_kouka_x_loot_out124), .loot_out125(_kouka_x_loot_out125), .loot_out126(_kouka_x_loot_out126), .loot_out127(_kouka_x_loot_out127), .loot_out128(_kouka_x_loot_out128), .loot_out129(_kouka_x_loot_out129), .loot_out130(_kouka_x_loot_out130), .loot_out131(_kouka_x_loot_out131), .loot_out132(_kouka_x_loot_out132), .loot_out133(_kouka_x_loot_out133), .loot_out134(_kouka_x_loot_out134), .loot_out135(_kouka_x_loot_out135), .loot_out136(_kouka_x_loot_out136), .loot_out137(_kouka_x_loot_out137), .loot_out138(_kouka_x_loot_out138), .loot_out139(_kouka_x_loot_out139), .loot_out140(_kouka_x_loot_out140), .loot_out141(_kouka_x_loot_out141), .loot_out142(_kouka_x_loot_out142), .loot_out143(_kouka_x_loot_out143), .loot_out144(_kouka_x_loot_out144), .loot_out145(_kouka_x_loot_out145), .loot_out146(_kouka_x_loot_out146), .loot_out147(_kouka_x_loot_out147), .loot_out148(_kouka_x_loot_out148), .loot_out149(_kouka_x_loot_out149), .loot_out150(_kouka_x_loot_out150), .loot_out151(_kouka_x_loot_out151), .loot_out152(_kouka_x_loot_out152), .loot_out153(_kouka_x_loot_out153), .loot_out154(_kouka_x_loot_out154), .loot_out155(_kouka_x_loot_out155), .loot_out156(_kouka_x_loot_out156), .loot_out157(_kouka_x_loot_out157), .loot_out158(_kouka_x_loot_out158), .loot_out159(_kouka_x_loot_out159), .loot_out160(_kouka_x_loot_out160), .loot_out161(_kouka_x_loot_out161), .loot_out162(_kouka_x_loot_out162), .loot_out163(_kouka_x_loot_out163), .loot_out164(_kouka_x_loot_out164), .loot_out165(_kouka_x_loot_out165), .loot_out166(_kouka_x_loot_out166), .loot_out167(_kouka_x_loot_out167), .loot_out168(_kouka_x_loot_out168), .loot_out169(_kouka_x_loot_out169), .loot_out170(_kouka_x_loot_out170), .loot_out171(_kouka_x_loot_out171), .loot_out172(_kouka_x_loot_out172), .loot_out173(_kouka_x_loot_out173), .loot_out174(_kouka_x_loot_out174), .loot_out175(_kouka_x_loot_out175), .loot_out176(_kouka_x_loot_out176), .loot_out177(_kouka_x_loot_out177), .loot_out178(_kouka_x_loot_out178), .loot_out179(_kouka_x_loot_out179), .loot_out180(_kouka_x_loot_out180), .loot_out181(_kouka_x_loot_out181), .loot_out182(_kouka_x_loot_out182), .loot_out183(_kouka_x_loot_out183), .loot_out184(_kouka_x_loot_out184), .loot_out185(_kouka_x_loot_out185), .loot_out186(_kouka_x_loot_out186), .loot_out187(_kouka_x_loot_out187), .loot_out188(_kouka_x_loot_out188), .loot_out189(_kouka_x_loot_out189), .loot_out190(_kouka_x_loot_out190), .loot_out191(_kouka_x_loot_out191), .loot_out192(_kouka_x_loot_out192), .loot_out193(_kouka_x_loot_out193), .loot_out194(_kouka_x_loot_out194), .loot_out195(_kouka_x_loot_out195), .loot_out196(_kouka_x_loot_out196), .loot_out197(_kouka_x_loot_out197), .loot_out198(_kouka_x_loot_out198), .loot_out199(_kouka_x_loot_out199), .loot_out200(_kouka_x_loot_out200), .loot_out201(_kouka_x_loot_out201), .loot_out202(_kouka_x_loot_out202), .loot_out203(_kouka_x_loot_out203), .loot_out204(_kouka_x_loot_out204), .loot_out205(_kouka_x_loot_out205), .loot_out206(_kouka_x_loot_out206), .loot_out207(_kouka_x_loot_out207), .loot_out208(_kouka_x_loot_out208), .loot_out209(_kouka_x_loot_out209), .loot_out210(_kouka_x_loot_out210), .loot_out211(_kouka_x_loot_out211), .loot_out212(_kouka_x_loot_out212), .loot_out213(_kouka_x_loot_out213), .loot_out214(_kouka_x_loot_out214), .loot_out215(_kouka_x_loot_out215), .loot_out216(_kouka_x_loot_out216), .loot_out217(_kouka_x_loot_out217), .loot_out218(_kouka_x_loot_out218), .loot_out219(_kouka_x_loot_out219), .loot_out220(_kouka_x_loot_out220), .loot_out221(_kouka_x_loot_out221), .loot_out222(_kouka_x_loot_out222), .data_in33(_kouka_x_data_in33), .data_in34(_kouka_x_data_in34), .data_in35(_kouka_x_data_in35), .data_in36(_kouka_x_data_in36), .data_in37(_kouka_x_data_in37), .data_in38(_kouka_x_data_in38), .data_in39(_kouka_x_data_in39), .data_in40(_kouka_x_data_in40), .data_in41(_kouka_x_data_in41), .data_in42(_kouka_x_data_in42), .data_in43(_kouka_x_data_in43), .data_in44(_kouka_x_data_in44), .data_in45(_kouka_x_data_in45), .data_in46(_kouka_x_data_in46), .data_in47(_kouka_x_data_in47), .data_in48(_kouka_x_data_in48), .data_in49(_kouka_x_data_in49), .data_in50(_kouka_x_data_in50), .data_in51(_kouka_x_data_in51), .data_in52(_kouka_x_data_in52), .data_in53(_kouka_x_data_in53), .data_in54(_kouka_x_data_in54), .data_in55(_kouka_x_data_in55), .data_in56(_kouka_x_data_in56), .data_in57(_kouka_x_data_in57), .data_in58(_kouka_x_data_in58), .data_in59(_kouka_x_data_in59), .data_in60(_kouka_x_data_in60), .data_in61(_kouka_x_data_in61), .data_in62(_kouka_x_data_in62), .data_in65(_kouka_x_data_in65), .data_in66(_kouka_x_data_in66), .data_in67(_kouka_x_data_in67), .data_in68(_kouka_x_data_in68), .data_in69(_kouka_x_data_in69), .data_in70(_kouka_x_data_in70), .data_in71(_kouka_x_data_in71), .data_in72(_kouka_x_data_in72), .data_in73(_kouka_x_data_in73), .data_in74(_kouka_x_data_in74), .data_in75(_kouka_x_data_in75), .data_in76(_kouka_x_data_in76), .data_in77(_kouka_x_data_in77), .data_in78(_kouka_x_data_in78), .data_in79(_kouka_x_data_in79), .data_in80(_kouka_x_data_in80), .data_in81(_kouka_x_data_in81), .data_in82(_kouka_x_data_in82), .data_in83(_kouka_x_data_in83), .data_in84(_kouka_x_data_in84), .data_in85(_kouka_x_data_in85), .data_in86(_kouka_x_data_in86), .data_in87(_kouka_x_data_in87), .data_in88(_kouka_x_data_in88), .data_in89(_kouka_x_data_in89), .data_in90(_kouka_x_data_in90), .data_in91(_kouka_x_data_in91), .data_in92(_kouka_x_data_in92), .data_in93(_kouka_x_data_in93), .data_in94(_kouka_x_data_in94), .data_in97(_kouka_x_data_in97), .data_in98(_kouka_x_data_in98), .data_in99(_kouka_x_data_in99), .data_in100(_kouka_x_data_in100), .data_in101(_kouka_x_data_in101), .data_in102(_kouka_x_data_in102), .data_in103(_kouka_x_data_in103), .data_in104(_kouka_x_data_in104), .data_in105(_kouka_x_data_in105), .data_in106(_kouka_x_data_in106), .data_in107(_kouka_x_data_in107), .data_in108(_kouka_x_data_in108), .data_in109(_kouka_x_data_in109), .data_in110(_kouka_x_data_in110), .data_in111(_kouka_x_data_in111), .data_in112(_kouka_x_data_in112), .data_in113(_kouka_x_data_in113), .data_in114(_kouka_x_data_in114), .data_in115(_kouka_x_data_in115), .data_in116(_kouka_x_data_in116), .data_in117(_kouka_x_data_in117), .data_in118(_kouka_x_data_in118), .data_in119(_kouka_x_data_in119), .data_in120(_kouka_x_data_in120), .data_in121(_kouka_x_data_in121), .data_in122(_kouka_x_data_in122), .data_in123(_kouka_x_data_in123), .data_in124(_kouka_x_data_in124), .data_in125(_kouka_x_data_in125), .data_in126(_kouka_x_data_in126), .data_in129(_kouka_x_data_in129), .data_in130(_kouka_x_data_in130), .data_in131(_kouka_x_data_in131), .data_in132(_kouka_x_data_in132), .data_in133(_kouka_x_data_in133), .data_in134(_kouka_x_data_in134), .data_in135(_kouka_x_data_in135), .data_in136(_kouka_x_data_in136), .data_in137(_kouka_x_data_in137), .data_in138(_kouka_x_data_in138), .data_in139(_kouka_x_data_in139), .data_in140(_kouka_x_data_in140), .data_in141(_kouka_x_data_in141), .data_in142(_kouka_x_data_in142), .data_in143(_kouka_x_data_in143), .data_in144(_kouka_x_data_in144), .data_in145(_kouka_x_data_in145), .data_in146(_kouka_x_data_in146), .data_in147(_kouka_x_data_in147), .data_in148(_kouka_x_data_in148), .data_in149(_kouka_x_data_in149), .data_in150(_kouka_x_data_in150), .data_in151(_kouka_x_data_in151), .data_in152(_kouka_x_data_in152), .data_in153(_kouka_x_data_in153), .data_in154(_kouka_x_data_in154), .data_in155(_kouka_x_data_in155), .data_in156(_kouka_x_data_in156), .data_in157(_kouka_x_data_in157), .data_in158(_kouka_x_data_in158), .data_in161(_kouka_x_data_in161), .data_in162(_kouka_x_data_in162), .data_in163(_kouka_x_data_in163), .data_in164(_kouka_x_data_in164), .data_in165(_kouka_x_data_in165), .data_in166(_kouka_x_data_in166), .data_in167(_kouka_x_data_in167), .data_in168(_kouka_x_data_in168), .data_in169(_kouka_x_data_in169), .data_in170(_kouka_x_data_in170), .data_in171(_kouka_x_data_in171), .data_in172(_kouka_x_data_in172), .data_in173(_kouka_x_data_in173), .data_in174(_kouka_x_data_in174), .data_in175(_kouka_x_data_in175), .data_in176(_kouka_x_data_in176), .data_in177(_kouka_x_data_in177), .data_in178(_kouka_x_data_in178), .data_in179(_kouka_x_data_in179), .data_in180(_kouka_x_data_in180), .data_in181(_kouka_x_data_in181), .data_in182(_kouka_x_data_in182), .data_in183(_kouka_x_data_in183), .data_in184(_kouka_x_data_in184), .data_in185(_kouka_x_data_in185), .data_in186(_kouka_x_data_in186), .data_in187(_kouka_x_data_in187), .data_in188(_kouka_x_data_in188), .data_in189(_kouka_x_data_in189), .data_in190(_kouka_x_data_in190), .data_in193(_kouka_x_data_in193), .data_in194(_kouka_x_data_in194), .data_in195(_kouka_x_data_in195), .data_in196(_kouka_x_data_in196), .data_in197(_kouka_x_data_in197), .data_in198(_kouka_x_data_in198), .data_in199(_kouka_x_data_in199), .data_in200(_kouka_x_data_in200), .data_in201(_kouka_x_data_in201), .data_in202(_kouka_x_data_in202), .data_in203(_kouka_x_data_in203), .data_in204(_kouka_x_data_in204), .data_in205(_kouka_x_data_in205), .data_in206(_kouka_x_data_in206), .data_in207(_kouka_x_data_in207), .data_in208(_kouka_x_data_in208), .data_in209(_kouka_x_data_in209), .data_in210(_kouka_x_data_in210), .data_in211(_kouka_x_data_in211), .data_in212(_kouka_x_data_in212), .data_in213(_kouka_x_data_in213), .data_in214(_kouka_x_data_in214), .data_in215(_kouka_x_data_in215), .data_in216(_kouka_x_data_in216), .data_in217(_kouka_x_data_in217), .data_in218(_kouka_x_data_in218), .data_in219(_kouka_x_data_in219), .data_in220(_kouka_x_data_in220), .data_in221(_kouka_x_data_in221), .data_in222(_kouka_x_data_in222), .data_in225(_kouka_x_data_in225), .data_in226(_kouka_x_data_in226), .data_in227(_kouka_x_data_in227), .data_in228(_kouka_x_data_in228), .data_in229(_kouka_x_data_in229), .data_in230(_kouka_x_data_in230), .data_in231(_kouka_x_data_in231), .data_in232(_kouka_x_data_in232), .data_in233(_kouka_x_data_in233), .data_in234(_kouka_x_data_in234), .data_in235(_kouka_x_data_in235), .data_in236(_kouka_x_data_in236), .data_in237(_kouka_x_data_in237), .data_in238(_kouka_x_data_in238), .data_in239(_kouka_x_data_in239), .data_in240(_kouka_x_data_in240), .data_in241(_kouka_x_data_in241), .data_in242(_kouka_x_data_in242), .data_in243(_kouka_x_data_in243), .data_in244(_kouka_x_data_in244), .data_in245(_kouka_x_data_in245), .data_in246(_kouka_x_data_in246), .data_in247(_kouka_x_data_in247), .data_in248(_kouka_x_data_in248), .data_in249(_kouka_x_data_in249), .data_in250(_kouka_x_data_in250), .data_in251(_kouka_x_data_in251), .data_in252(_kouka_x_data_in252), .data_in253(_kouka_x_data_in253), .data_in254(_kouka_x_data_in254), .data_in257(_kouka_x_data_in257), .data_in258(_kouka_x_data_in258), .data_in259(_kouka_x_data_in259), .data_in260(_kouka_x_data_in260), .data_in261(_kouka_x_data_in261), .data_in262(_kouka_x_data_in262), .data_in263(_kouka_x_data_in263), .data_in264(_kouka_x_data_in264), .data_in265(_kouka_x_data_in265), .data_in266(_kouka_x_data_in266), .data_in267(_kouka_x_data_in267), .data_in268(_kouka_x_data_in268), .data_in269(_kouka_x_data_in269), .data_in270(_kouka_x_data_in270), .data_in271(_kouka_x_data_in271), .data_in272(_kouka_x_data_in272), .data_in273(_kouka_x_data_in273), .data_in274(_kouka_x_data_in274), .data_in275(_kouka_x_data_in275), .data_in276(_kouka_x_data_in276), .data_in277(_kouka_x_data_in277), .data_in278(_kouka_x_data_in278), .data_in279(_kouka_x_data_in279), .data_in280(_kouka_x_data_in280), .data_in281(_kouka_x_data_in281), .data_in282(_kouka_x_data_in282), .data_in283(_kouka_x_data_in283), .data_in284(_kouka_x_data_in284), .data_in285(_kouka_x_data_in285), .data_in286(_kouka_x_data_in286), .data_in289(_kouka_x_data_in289), .data_in290(_kouka_x_data_in290), .data_in291(_kouka_x_data_in291), .data_in292(_kouka_x_data_in292), .data_in293(_kouka_x_data_in293), .data_in294(_kouka_x_data_in294), .data_in295(_kouka_x_data_in295), .data_in296(_kouka_x_data_in296), .data_in297(_kouka_x_data_in297), .data_in298(_kouka_x_data_in298), .data_in299(_kouka_x_data_in299), .data_in300(_kouka_x_data_in300), .data_in301(_kouka_x_data_in301), .data_in302(_kouka_x_data_in302), .data_in303(_kouka_x_data_in303), .data_in304(_kouka_x_data_in304), .data_in305(_kouka_x_data_in305), .data_in306(_kouka_x_data_in306), .data_in307(_kouka_x_data_in307), .data_in308(_kouka_x_data_in308), .data_in309(_kouka_x_data_in309), .data_in310(_kouka_x_data_in310), .data_in311(_kouka_x_data_in311), .data_in312(_kouka_x_data_in312), .data_in313(_kouka_x_data_in313), .data_in314(_kouka_x_data_in314), .data_in315(_kouka_x_data_in315), .data_in316(_kouka_x_data_in316), .data_in317(_kouka_x_data_in317), .data_in318(_kouka_x_data_in318), .data_in321(_kouka_x_data_in321), .data_in322(_kouka_x_data_in322), .data_in323(_kouka_x_data_in323), .data_in324(_kouka_x_data_in324), .data_in325(_kouka_x_data_in325), .data_in326(_kouka_x_data_in326), .data_in327(_kouka_x_data_in327), .data_in328(_kouka_x_data_in328), .data_in329(_kouka_x_data_in329), .data_in330(_kouka_x_data_in330), .data_in331(_kouka_x_data_in331), .data_in332(_kouka_x_data_in332), .data_in333(_kouka_x_data_in333), .data_in334(_kouka_x_data_in334), .data_in335(_kouka_x_data_in335), .data_in336(_kouka_x_data_in336), .data_in337(_kouka_x_data_in337), .data_in338(_kouka_x_data_in338), .data_in339(_kouka_x_data_in339), .data_in340(_kouka_x_data_in340), .data_in341(_kouka_x_data_in341), .data_in342(_kouka_x_data_in342), .data_in343(_kouka_x_data_in343), .data_in344(_kouka_x_data_in344), .data_in345(_kouka_x_data_in345), .data_in346(_kouka_x_data_in346), .data_in347(_kouka_x_data_in347), .data_in348(_kouka_x_data_in348), .data_in349(_kouka_x_data_in349), .data_in350(_kouka_x_data_in350), .data_in353(_kouka_x_data_in353), .data_in354(_kouka_x_data_in354), .data_in355(_kouka_x_data_in355), .data_in356(_kouka_x_data_in356), .data_in357(_kouka_x_data_in357), .data_in358(_kouka_x_data_in358), .data_in359(_kouka_x_data_in359), .data_in360(_kouka_x_data_in360), .data_in361(_kouka_x_data_in361), .data_in362(_kouka_x_data_in362), .data_in363(_kouka_x_data_in363), .data_in364(_kouka_x_data_in364), .data_in365(_kouka_x_data_in365), .data_in366(_kouka_x_data_in366), .data_in367(_kouka_x_data_in367), .data_in368(_kouka_x_data_in368), .data_in369(_kouka_x_data_in369), .data_in370(_kouka_x_data_in370), .data_in371(_kouka_x_data_in371), .data_in372(_kouka_x_data_in372), .data_in373(_kouka_x_data_in373), .data_in374(_kouka_x_data_in374), .data_in375(_kouka_x_data_in375), .data_in376(_kouka_x_data_in376), .data_in377(_kouka_x_data_in377), .data_in378(_kouka_x_data_in378), .data_in379(_kouka_x_data_in379), .data_in380(_kouka_x_data_in380), .data_in381(_kouka_x_data_in381), .data_in382(_kouka_x_data_in382), .data_in385(_kouka_x_data_in385), .data_in386(_kouka_x_data_in386), .data_in387(_kouka_x_data_in387), .data_in388(_kouka_x_data_in388), .data_in389(_kouka_x_data_in389), .data_in390(_kouka_x_data_in390), .data_in391(_kouka_x_data_in391), .data_in392(_kouka_x_data_in392), .data_in393(_kouka_x_data_in393), .data_in394(_kouka_x_data_in394), .data_in395(_kouka_x_data_in395), .data_in396(_kouka_x_data_in396), .data_in397(_kouka_x_data_in397), .data_in398(_kouka_x_data_in398), .data_in399(_kouka_x_data_in399), .data_in400(_kouka_x_data_in400), .data_in401(_kouka_x_data_in401), .data_in402(_kouka_x_data_in402), .data_in403(_kouka_x_data_in403), .data_in404(_kouka_x_data_in404), .data_in405(_kouka_x_data_in405), .data_in406(_kouka_x_data_in406), .data_in407(_kouka_x_data_in407), .data_in408(_kouka_x_data_in408), .data_in409(_kouka_x_data_in409), .data_in410(_kouka_x_data_in410), .data_in411(_kouka_x_data_in411), .data_in412(_kouka_x_data_in412), .data_in413(_kouka_x_data_in413), .data_in414(_kouka_x_data_in414), .data_in417(_kouka_x_data_in417), .data_in418(_kouka_x_data_in418), .data_in419(_kouka_x_data_in419), .data_in420(_kouka_x_data_in420), .data_in421(_kouka_x_data_in421), .data_in422(_kouka_x_data_in422), .data_in423(_kouka_x_data_in423), .data_in424(_kouka_x_data_in424), .data_in425(_kouka_x_data_in425), .data_in426(_kouka_x_data_in426), .data_in427(_kouka_x_data_in427), .data_in428(_kouka_x_data_in428), .data_in429(_kouka_x_data_in429), .data_in430(_kouka_x_data_in430), .data_in431(_kouka_x_data_in431), .data_in432(_kouka_x_data_in432), .data_in433(_kouka_x_data_in433), .data_in434(_kouka_x_data_in434), .data_in435(_kouka_x_data_in435), .data_in436(_kouka_x_data_in436), .data_in437(_kouka_x_data_in437), .data_in438(_kouka_x_data_in438), .data_in439(_kouka_x_data_in439), .data_in440(_kouka_x_data_in440), .data_in441(_kouka_x_data_in441), .data_in442(_kouka_x_data_in442), .data_in443(_kouka_x_data_in443), .data_in444(_kouka_x_data_in444), .data_in445(_kouka_x_data_in445), .data_in446(_kouka_x_data_in446), .data_in449(_kouka_x_data_in449), .data_in450(_kouka_x_data_in450), .data_in451(_kouka_x_data_in451), .data_in452(_kouka_x_data_in452), .data_in453(_kouka_x_data_in453), .data_in454(_kouka_x_data_in454), .data_in455(_kouka_x_data_in455), .data_in456(_kouka_x_data_in456), .data_in457(_kouka_x_data_in457), .data_in458(_kouka_x_data_in458), .data_in459(_kouka_x_data_in459), .data_in460(_kouka_x_data_in460), .data_in461(_kouka_x_data_in461), .data_in462(_kouka_x_data_in462), .data_in463(_kouka_x_data_in463), .data_in464(_kouka_x_data_in464), .data_in465(_kouka_x_data_in465), .data_in466(_kouka_x_data_in466), .data_in467(_kouka_x_data_in467), .data_in468(_kouka_x_data_in468), .data_in469(_kouka_x_data_in469), .data_in470(_kouka_x_data_in470), .data_in471(_kouka_x_data_in471), .data_in472(_kouka_x_data_in472), .data_in473(_kouka_x_data_in473), .data_in474(_kouka_x_data_in474), .data_in475(_kouka_x_data_in475), .data_in476(_kouka_x_data_in476), .data_in477(_kouka_x_data_in477), .data_in478(_kouka_x_data_in478), .start(_kouka_x_start), .goal(_kouka_x_goal));
kanwa kanwa_x (.m_clock(m_clock), .p_reset( p_reset), .out_do(_kanwa_x_out_do), .in_do(_kanwa_x_in_do), .data_out33(_kanwa_x_data_out33), .data_out34(_kanwa_x_data_out34), .data_out35(_kanwa_x_data_out35), .data_out36(_kanwa_x_data_out36), .data_out37(_kanwa_x_data_out37), .data_out38(_kanwa_x_data_out38), .data_out39(_kanwa_x_data_out39), .data_out40(_kanwa_x_data_out40), .data_out41(_kanwa_x_data_out41), .data_out42(_kanwa_x_data_out42), .data_out43(_kanwa_x_data_out43), .data_out44(_kanwa_x_data_out44), .data_out45(_kanwa_x_data_out45), .data_out46(_kanwa_x_data_out46), .data_out47(_kanwa_x_data_out47), .data_out48(_kanwa_x_data_out48), .data_out49(_kanwa_x_data_out49), .data_out50(_kanwa_x_data_out50), .data_out51(_kanwa_x_data_out51), .data_out52(_kanwa_x_data_out52), .data_out53(_kanwa_x_data_out53), .data_out54(_kanwa_x_data_out54), .data_out55(_kanwa_x_data_out55), .data_out56(_kanwa_x_data_out56), .data_out57(_kanwa_x_data_out57), .data_out58(_kanwa_x_data_out58), .data_out59(_kanwa_x_data_out59), .data_out60(_kanwa_x_data_out60), .data_out61(_kanwa_x_data_out61), .data_out62(_kanwa_x_data_out62), .data_out65(_kanwa_x_data_out65), .data_out66(_kanwa_x_data_out66), .data_out67(_kanwa_x_data_out67), .data_out68(_kanwa_x_data_out68), .data_out69(_kanwa_x_data_out69), .data_out70(_kanwa_x_data_out70), .data_out71(_kanwa_x_data_out71), .data_out72(_kanwa_x_data_out72), .data_out73(_kanwa_x_data_out73), .data_out74(_kanwa_x_data_out74), .data_out75(_kanwa_x_data_out75), .data_out76(_kanwa_x_data_out76), .data_out77(_kanwa_x_data_out77), .data_out78(_kanwa_x_data_out78), .data_out79(_kanwa_x_data_out79), .data_out80(_kanwa_x_data_out80), .data_out81(_kanwa_x_data_out81), .data_out82(_kanwa_x_data_out82), .data_out83(_kanwa_x_data_out83), .data_out84(_kanwa_x_data_out84), .data_out85(_kanwa_x_data_out85), .data_out86(_kanwa_x_data_out86), .data_out87(_kanwa_x_data_out87), .data_out88(_kanwa_x_data_out88), .data_out89(_kanwa_x_data_out89), .data_out90(_kanwa_x_data_out90), .data_out91(_kanwa_x_data_out91), .data_out92(_kanwa_x_data_out92), .data_out93(_kanwa_x_data_out93), .data_out94(_kanwa_x_data_out94), .data_out97(_kanwa_x_data_out97), .data_out98(_kanwa_x_data_out98), .data_out99(_kanwa_x_data_out99), .data_out100(_kanwa_x_data_out100), .data_out101(_kanwa_x_data_out101), .data_out102(_kanwa_x_data_out102), .data_out103(_kanwa_x_data_out103), .data_out104(_kanwa_x_data_out104), .data_out105(_kanwa_x_data_out105), .data_out106(_kanwa_x_data_out106), .data_out107(_kanwa_x_data_out107), .data_out108(_kanwa_x_data_out108), .data_out109(_kanwa_x_data_out109), .data_out110(_kanwa_x_data_out110), .data_out111(_kanwa_x_data_out111), .data_out112(_kanwa_x_data_out112), .data_out113(_kanwa_x_data_out113), .data_out114(_kanwa_x_data_out114), .data_out115(_kanwa_x_data_out115), .data_out116(_kanwa_x_data_out116), .data_out117(_kanwa_x_data_out117), .data_out118(_kanwa_x_data_out118), .data_out119(_kanwa_x_data_out119), .data_out120(_kanwa_x_data_out120), .data_out121(_kanwa_x_data_out121), .data_out122(_kanwa_x_data_out122), .data_out123(_kanwa_x_data_out123), .data_out124(_kanwa_x_data_out124), .data_out125(_kanwa_x_data_out125), .data_out126(_kanwa_x_data_out126), .data_out129(_kanwa_x_data_out129), .data_out130(_kanwa_x_data_out130), .data_out131(_kanwa_x_data_out131), .data_out132(_kanwa_x_data_out132), .data_out133(_kanwa_x_data_out133), .data_out134(_kanwa_x_data_out134), .data_out135(_kanwa_x_data_out135), .data_out136(_kanwa_x_data_out136), .data_out137(_kanwa_x_data_out137), .data_out138(_kanwa_x_data_out138), .data_out139(_kanwa_x_data_out139), .data_out140(_kanwa_x_data_out140), .data_out141(_kanwa_x_data_out141), .data_out142(_kanwa_x_data_out142), .data_out143(_kanwa_x_data_out143), .data_out144(_kanwa_x_data_out144), .data_out145(_kanwa_x_data_out145), .data_out146(_kanwa_x_data_out146), .data_out147(_kanwa_x_data_out147), .data_out148(_kanwa_x_data_out148), .data_out149(_kanwa_x_data_out149), .data_out150(_kanwa_x_data_out150), .data_out151(_kanwa_x_data_out151), .data_out152(_kanwa_x_data_out152), .data_out153(_kanwa_x_data_out153), .data_out154(_kanwa_x_data_out154), .data_out155(_kanwa_x_data_out155), .data_out156(_kanwa_x_data_out156), .data_out157(_kanwa_x_data_out157), .data_out158(_kanwa_x_data_out158), .data_out161(_kanwa_x_data_out161), .data_out162(_kanwa_x_data_out162), .data_out163(_kanwa_x_data_out163), .data_out164(_kanwa_x_data_out164), .data_out165(_kanwa_x_data_out165), .data_out166(_kanwa_x_data_out166), .data_out167(_kanwa_x_data_out167), .data_out168(_kanwa_x_data_out168), .data_out169(_kanwa_x_data_out169), .data_out170(_kanwa_x_data_out170), .data_out171(_kanwa_x_data_out171), .data_out172(_kanwa_x_data_out172), .data_out173(_kanwa_x_data_out173), .data_out174(_kanwa_x_data_out174), .data_out175(_kanwa_x_data_out175), .data_out176(_kanwa_x_data_out176), .data_out177(_kanwa_x_data_out177), .data_out178(_kanwa_x_data_out178), .data_out179(_kanwa_x_data_out179), .data_out180(_kanwa_x_data_out180), .data_out181(_kanwa_x_data_out181), .data_out182(_kanwa_x_data_out182), .data_out183(_kanwa_x_data_out183), .data_out184(_kanwa_x_data_out184), .data_out185(_kanwa_x_data_out185), .data_out186(_kanwa_x_data_out186), .data_out187(_kanwa_x_data_out187), .data_out188(_kanwa_x_data_out188), .data_out189(_kanwa_x_data_out189), .data_out190(_kanwa_x_data_out190), .data_out193(_kanwa_x_data_out193), .data_out194(_kanwa_x_data_out194), .data_out195(_kanwa_x_data_out195), .data_out196(_kanwa_x_data_out196), .data_out197(_kanwa_x_data_out197), .data_out198(_kanwa_x_data_out198), .data_out199(_kanwa_x_data_out199), .data_out200(_kanwa_x_data_out200), .data_out201(_kanwa_x_data_out201), .data_out202(_kanwa_x_data_out202), .data_out203(_kanwa_x_data_out203), .data_out204(_kanwa_x_data_out204), .data_out205(_kanwa_x_data_out205), .data_out206(_kanwa_x_data_out206), .data_out207(_kanwa_x_data_out207), .data_out208(_kanwa_x_data_out208), .data_out209(_kanwa_x_data_out209), .data_out210(_kanwa_x_data_out210), .data_out211(_kanwa_x_data_out211), .data_out212(_kanwa_x_data_out212), .data_out213(_kanwa_x_data_out213), .data_out214(_kanwa_x_data_out214), .data_out215(_kanwa_x_data_out215), .data_out216(_kanwa_x_data_out216), .data_out217(_kanwa_x_data_out217), .data_out218(_kanwa_x_data_out218), .data_out219(_kanwa_x_data_out219), .data_out220(_kanwa_x_data_out220), .data_out221(_kanwa_x_data_out221), .data_out222(_kanwa_x_data_out222), .data_out225(_kanwa_x_data_out225), .data_out226(_kanwa_x_data_out226), .data_out227(_kanwa_x_data_out227), .data_out228(_kanwa_x_data_out228), .data_out229(_kanwa_x_data_out229), .data_out230(_kanwa_x_data_out230), .data_out231(_kanwa_x_data_out231), .data_out232(_kanwa_x_data_out232), .data_out233(_kanwa_x_data_out233), .data_out234(_kanwa_x_data_out234), .data_out235(_kanwa_x_data_out235), .data_out236(_kanwa_x_data_out236), .data_out237(_kanwa_x_data_out237), .data_out238(_kanwa_x_data_out238), .data_out239(_kanwa_x_data_out239), .data_out240(_kanwa_x_data_out240), .data_out241(_kanwa_x_data_out241), .data_out242(_kanwa_x_data_out242), .data_out243(_kanwa_x_data_out243), .data_out244(_kanwa_x_data_out244), .data_out245(_kanwa_x_data_out245), .data_out246(_kanwa_x_data_out246), .data_out247(_kanwa_x_data_out247), .data_out248(_kanwa_x_data_out248), .data_out249(_kanwa_x_data_out249), .data_out250(_kanwa_x_data_out250), .data_out251(_kanwa_x_data_out251), .data_out252(_kanwa_x_data_out252), .data_out253(_kanwa_x_data_out253), .data_out254(_kanwa_x_data_out254), .data_out257(_kanwa_x_data_out257), .data_out258(_kanwa_x_data_out258), .data_out259(_kanwa_x_data_out259), .data_out260(_kanwa_x_data_out260), .data_out261(_kanwa_x_data_out261), .data_out262(_kanwa_x_data_out262), .data_out263(_kanwa_x_data_out263), .data_out264(_kanwa_x_data_out264), .data_out265(_kanwa_x_data_out265), .data_out266(_kanwa_x_data_out266), .data_out267(_kanwa_x_data_out267), .data_out268(_kanwa_x_data_out268), .data_out269(_kanwa_x_data_out269), .data_out270(_kanwa_x_data_out270), .data_out271(_kanwa_x_data_out271), .data_out272(_kanwa_x_data_out272), .data_out273(_kanwa_x_data_out273), .data_out274(_kanwa_x_data_out274), .data_out275(_kanwa_x_data_out275), .data_out276(_kanwa_x_data_out276), .data_out277(_kanwa_x_data_out277), .data_out278(_kanwa_x_data_out278), .data_out279(_kanwa_x_data_out279), .data_out280(_kanwa_x_data_out280), .data_out281(_kanwa_x_data_out281), .data_out282(_kanwa_x_data_out282), .data_out283(_kanwa_x_data_out283), .data_out284(_kanwa_x_data_out284), .data_out285(_kanwa_x_data_out285), .data_out286(_kanwa_x_data_out286), .data_out289(_kanwa_x_data_out289), .data_out290(_kanwa_x_data_out290), .data_out291(_kanwa_x_data_out291), .data_out292(_kanwa_x_data_out292), .data_out293(_kanwa_x_data_out293), .data_out294(_kanwa_x_data_out294), .data_out295(_kanwa_x_data_out295), .data_out296(_kanwa_x_data_out296), .data_out297(_kanwa_x_data_out297), .data_out298(_kanwa_x_data_out298), .data_out299(_kanwa_x_data_out299), .data_out300(_kanwa_x_data_out300), .data_out301(_kanwa_x_data_out301), .data_out302(_kanwa_x_data_out302), .data_out303(_kanwa_x_data_out303), .data_out304(_kanwa_x_data_out304), .data_out305(_kanwa_x_data_out305), .data_out306(_kanwa_x_data_out306), .data_out307(_kanwa_x_data_out307), .data_out308(_kanwa_x_data_out308), .data_out309(_kanwa_x_data_out309), .data_out310(_kanwa_x_data_out310), .data_out311(_kanwa_x_data_out311), .data_out312(_kanwa_x_data_out312), .data_out313(_kanwa_x_data_out313), .data_out314(_kanwa_x_data_out314), .data_out315(_kanwa_x_data_out315), .data_out316(_kanwa_x_data_out316), .data_out317(_kanwa_x_data_out317), .data_out318(_kanwa_x_data_out318), .data_out321(_kanwa_x_data_out321), .data_out322(_kanwa_x_data_out322), .data_out323(_kanwa_x_data_out323), .data_out324(_kanwa_x_data_out324), .data_out325(_kanwa_x_data_out325), .data_out326(_kanwa_x_data_out326), .data_out327(_kanwa_x_data_out327), .data_out328(_kanwa_x_data_out328), .data_out329(_kanwa_x_data_out329), .data_out330(_kanwa_x_data_out330), .data_out331(_kanwa_x_data_out331), .data_out332(_kanwa_x_data_out332), .data_out333(_kanwa_x_data_out333), .data_out334(_kanwa_x_data_out334), .data_out335(_kanwa_x_data_out335), .data_out336(_kanwa_x_data_out336), .data_out337(_kanwa_x_data_out337), .data_out338(_kanwa_x_data_out338), .data_out339(_kanwa_x_data_out339), .data_out340(_kanwa_x_data_out340), .data_out341(_kanwa_x_data_out341), .data_out342(_kanwa_x_data_out342), .data_out343(_kanwa_x_data_out343), .data_out344(_kanwa_x_data_out344), .data_out345(_kanwa_x_data_out345), .data_out346(_kanwa_x_data_out346), .data_out347(_kanwa_x_data_out347), .data_out348(_kanwa_x_data_out348), .data_out349(_kanwa_x_data_out349), .data_out350(_kanwa_x_data_out350), .data_out353(_kanwa_x_data_out353), .data_out354(_kanwa_x_data_out354), .data_out355(_kanwa_x_data_out355), .data_out356(_kanwa_x_data_out356), .data_out357(_kanwa_x_data_out357), .data_out358(_kanwa_x_data_out358), .data_out359(_kanwa_x_data_out359), .data_out360(_kanwa_x_data_out360), .data_out361(_kanwa_x_data_out361), .data_out362(_kanwa_x_data_out362), .data_out363(_kanwa_x_data_out363), .data_out364(_kanwa_x_data_out364), .data_out365(_kanwa_x_data_out365), .data_out366(_kanwa_x_data_out366), .data_out367(_kanwa_x_data_out367), .data_out368(_kanwa_x_data_out368), .data_out369(_kanwa_x_data_out369), .data_out370(_kanwa_x_data_out370), .data_out371(_kanwa_x_data_out371), .data_out372(_kanwa_x_data_out372), .data_out373(_kanwa_x_data_out373), .data_out374(_kanwa_x_data_out374), .data_out375(_kanwa_x_data_out375), .data_out376(_kanwa_x_data_out376), .data_out377(_kanwa_x_data_out377), .data_out378(_kanwa_x_data_out378), .data_out379(_kanwa_x_data_out379), .data_out380(_kanwa_x_data_out380), .data_out381(_kanwa_x_data_out381), .data_out382(_kanwa_x_data_out382), .data_out385(_kanwa_x_data_out385), .data_out386(_kanwa_x_data_out386), .data_out387(_kanwa_x_data_out387), .data_out388(_kanwa_x_data_out388), .data_out389(_kanwa_x_data_out389), .data_out390(_kanwa_x_data_out390), .data_out391(_kanwa_x_data_out391), .data_out392(_kanwa_x_data_out392), .data_out393(_kanwa_x_data_out393), .data_out394(_kanwa_x_data_out394), .data_out395(_kanwa_x_data_out395), .data_out396(_kanwa_x_data_out396), .data_out397(_kanwa_x_data_out397), .data_out398(_kanwa_x_data_out398), .data_out399(_kanwa_x_data_out399), .data_out400(_kanwa_x_data_out400), .data_out401(_kanwa_x_data_out401), .data_out402(_kanwa_x_data_out402), .data_out403(_kanwa_x_data_out403), .data_out404(_kanwa_x_data_out404), .data_out405(_kanwa_x_data_out405), .data_out406(_kanwa_x_data_out406), .data_out407(_kanwa_x_data_out407), .data_out408(_kanwa_x_data_out408), .data_out409(_kanwa_x_data_out409), .data_out410(_kanwa_x_data_out410), .data_out411(_kanwa_x_data_out411), .data_out412(_kanwa_x_data_out412), .data_out413(_kanwa_x_data_out413), .data_out414(_kanwa_x_data_out414), .data_out417(_kanwa_x_data_out417), .data_out418(_kanwa_x_data_out418), .data_out419(_kanwa_x_data_out419), .data_out420(_kanwa_x_data_out420), .data_out421(_kanwa_x_data_out421), .data_out422(_kanwa_x_data_out422), .data_out423(_kanwa_x_data_out423), .data_out424(_kanwa_x_data_out424), .data_out425(_kanwa_x_data_out425), .data_out426(_kanwa_x_data_out426), .data_out427(_kanwa_x_data_out427), .data_out428(_kanwa_x_data_out428), .data_out429(_kanwa_x_data_out429), .data_out430(_kanwa_x_data_out430), .data_out431(_kanwa_x_data_out431), .data_out432(_kanwa_x_data_out432), .data_out433(_kanwa_x_data_out433), .data_out434(_kanwa_x_data_out434), .data_out435(_kanwa_x_data_out435), .data_out436(_kanwa_x_data_out436), .data_out437(_kanwa_x_data_out437), .data_out438(_kanwa_x_data_out438), .data_out439(_kanwa_x_data_out439), .data_out440(_kanwa_x_data_out440), .data_out441(_kanwa_x_data_out441), .data_out442(_kanwa_x_data_out442), .data_out443(_kanwa_x_data_out443), .data_out444(_kanwa_x_data_out444), .data_out445(_kanwa_x_data_out445), .data_out446(_kanwa_x_data_out446), .data_out449(_kanwa_x_data_out449), .data_out450(_kanwa_x_data_out450), .data_out451(_kanwa_x_data_out451), .data_out452(_kanwa_x_data_out452), .data_out453(_kanwa_x_data_out453), .data_out454(_kanwa_x_data_out454), .data_out455(_kanwa_x_data_out455), .data_out456(_kanwa_x_data_out456), .data_out457(_kanwa_x_data_out457), .data_out458(_kanwa_x_data_out458), .data_out459(_kanwa_x_data_out459), .data_out460(_kanwa_x_data_out460), .data_out461(_kanwa_x_data_out461), .data_out462(_kanwa_x_data_out462), .data_out463(_kanwa_x_data_out463), .data_out464(_kanwa_x_data_out464), .data_out465(_kanwa_x_data_out465), .data_out466(_kanwa_x_data_out466), .data_out467(_kanwa_x_data_out467), .data_out468(_kanwa_x_data_out468), .data_out469(_kanwa_x_data_out469), .data_out470(_kanwa_x_data_out470), .data_out471(_kanwa_x_data_out471), .data_out472(_kanwa_x_data_out472), .data_out473(_kanwa_x_data_out473), .data_out474(_kanwa_x_data_out474), .data_out475(_kanwa_x_data_out475), .data_out476(_kanwa_x_data_out476), .data_out477(_kanwa_x_data_out477), .data_out478(_kanwa_x_data_out478), .data_in33(_kanwa_x_data_in33), .data_in34(_kanwa_x_data_in34), .data_in35(_kanwa_x_data_in35), .data_in36(_kanwa_x_data_in36), .data_in37(_kanwa_x_data_in37), .data_in38(_kanwa_x_data_in38), .data_in39(_kanwa_x_data_in39), .data_in40(_kanwa_x_data_in40), .data_in41(_kanwa_x_data_in41), .data_in42(_kanwa_x_data_in42), .data_in43(_kanwa_x_data_in43), .data_in44(_kanwa_x_data_in44), .data_in45(_kanwa_x_data_in45), .data_in46(_kanwa_x_data_in46), .data_in47(_kanwa_x_data_in47), .data_in48(_kanwa_x_data_in48), .data_in49(_kanwa_x_data_in49), .data_in50(_kanwa_x_data_in50), .data_in51(_kanwa_x_data_in51), .data_in52(_kanwa_x_data_in52), .data_in53(_kanwa_x_data_in53), .data_in54(_kanwa_x_data_in54), .data_in55(_kanwa_x_data_in55), .data_in56(_kanwa_x_data_in56), .data_in57(_kanwa_x_data_in57), .data_in58(_kanwa_x_data_in58), .data_in59(_kanwa_x_data_in59), .data_in60(_kanwa_x_data_in60), .data_in61(_kanwa_x_data_in61), .data_in62(_kanwa_x_data_in62), .data_in65(_kanwa_x_data_in65), .data_in66(_kanwa_x_data_in66), .data_in67(_kanwa_x_data_in67), .data_in68(_kanwa_x_data_in68), .data_in69(_kanwa_x_data_in69), .data_in70(_kanwa_x_data_in70), .data_in71(_kanwa_x_data_in71), .data_in72(_kanwa_x_data_in72), .data_in73(_kanwa_x_data_in73), .data_in74(_kanwa_x_data_in74), .data_in75(_kanwa_x_data_in75), .data_in76(_kanwa_x_data_in76), .data_in77(_kanwa_x_data_in77), .data_in78(_kanwa_x_data_in78), .data_in79(_kanwa_x_data_in79), .data_in80(_kanwa_x_data_in80), .data_in81(_kanwa_x_data_in81), .data_in82(_kanwa_x_data_in82), .data_in83(_kanwa_x_data_in83), .data_in84(_kanwa_x_data_in84), .data_in85(_kanwa_x_data_in85), .data_in86(_kanwa_x_data_in86), .data_in87(_kanwa_x_data_in87), .data_in88(_kanwa_x_data_in88), .data_in89(_kanwa_x_data_in89), .data_in90(_kanwa_x_data_in90), .data_in91(_kanwa_x_data_in91), .data_in92(_kanwa_x_data_in92), .data_in93(_kanwa_x_data_in93), .data_in94(_kanwa_x_data_in94), .data_in97(_kanwa_x_data_in97), .data_in98(_kanwa_x_data_in98), .data_in99(_kanwa_x_data_in99), .data_in100(_kanwa_x_data_in100), .data_in101(_kanwa_x_data_in101), .data_in102(_kanwa_x_data_in102), .data_in103(_kanwa_x_data_in103), .data_in104(_kanwa_x_data_in104), .data_in105(_kanwa_x_data_in105), .data_in106(_kanwa_x_data_in106), .data_in107(_kanwa_x_data_in107), .data_in108(_kanwa_x_data_in108), .data_in109(_kanwa_x_data_in109), .data_in110(_kanwa_x_data_in110), .data_in111(_kanwa_x_data_in111), .data_in112(_kanwa_x_data_in112), .data_in113(_kanwa_x_data_in113), .data_in114(_kanwa_x_data_in114), .data_in115(_kanwa_x_data_in115), .data_in116(_kanwa_x_data_in116), .data_in117(_kanwa_x_data_in117), .data_in118(_kanwa_x_data_in118), .data_in119(_kanwa_x_data_in119), .data_in120(_kanwa_x_data_in120), .data_in121(_kanwa_x_data_in121), .data_in122(_kanwa_x_data_in122), .data_in123(_kanwa_x_data_in123), .data_in124(_kanwa_x_data_in124), .data_in125(_kanwa_x_data_in125), .data_in126(_kanwa_x_data_in126), .data_in129(_kanwa_x_data_in129), .data_in130(_kanwa_x_data_in130), .data_in131(_kanwa_x_data_in131), .data_in132(_kanwa_x_data_in132), .data_in133(_kanwa_x_data_in133), .data_in134(_kanwa_x_data_in134), .data_in135(_kanwa_x_data_in135), .data_in136(_kanwa_x_data_in136), .data_in137(_kanwa_x_data_in137), .data_in138(_kanwa_x_data_in138), .data_in139(_kanwa_x_data_in139), .data_in140(_kanwa_x_data_in140), .data_in141(_kanwa_x_data_in141), .data_in142(_kanwa_x_data_in142), .data_in143(_kanwa_x_data_in143), .data_in144(_kanwa_x_data_in144), .data_in145(_kanwa_x_data_in145), .data_in146(_kanwa_x_data_in146), .data_in147(_kanwa_x_data_in147), .data_in148(_kanwa_x_data_in148), .data_in149(_kanwa_x_data_in149), .data_in150(_kanwa_x_data_in150), .data_in151(_kanwa_x_data_in151), .data_in152(_kanwa_x_data_in152), .data_in153(_kanwa_x_data_in153), .data_in154(_kanwa_x_data_in154), .data_in155(_kanwa_x_data_in155), .data_in156(_kanwa_x_data_in156), .data_in157(_kanwa_x_data_in157), .data_in158(_kanwa_x_data_in158), .data_in161(_kanwa_x_data_in161), .data_in162(_kanwa_x_data_in162), .data_in163(_kanwa_x_data_in163), .data_in164(_kanwa_x_data_in164), .data_in165(_kanwa_x_data_in165), .data_in166(_kanwa_x_data_in166), .data_in167(_kanwa_x_data_in167), .data_in168(_kanwa_x_data_in168), .data_in169(_kanwa_x_data_in169), .data_in170(_kanwa_x_data_in170), .data_in171(_kanwa_x_data_in171), .data_in172(_kanwa_x_data_in172), .data_in173(_kanwa_x_data_in173), .data_in174(_kanwa_x_data_in174), .data_in175(_kanwa_x_data_in175), .data_in176(_kanwa_x_data_in176), .data_in177(_kanwa_x_data_in177), .data_in178(_kanwa_x_data_in178), .data_in179(_kanwa_x_data_in179), .data_in180(_kanwa_x_data_in180), .data_in181(_kanwa_x_data_in181), .data_in182(_kanwa_x_data_in182), .data_in183(_kanwa_x_data_in183), .data_in184(_kanwa_x_data_in184), .data_in185(_kanwa_x_data_in185), .data_in186(_kanwa_x_data_in186), .data_in187(_kanwa_x_data_in187), .data_in188(_kanwa_x_data_in188), .data_in189(_kanwa_x_data_in189), .data_in190(_kanwa_x_data_in190), .data_in193(_kanwa_x_data_in193), .data_in194(_kanwa_x_data_in194), .data_in195(_kanwa_x_data_in195), .data_in196(_kanwa_x_data_in196), .data_in197(_kanwa_x_data_in197), .data_in198(_kanwa_x_data_in198), .data_in199(_kanwa_x_data_in199), .data_in200(_kanwa_x_data_in200), .data_in201(_kanwa_x_data_in201), .data_in202(_kanwa_x_data_in202), .data_in203(_kanwa_x_data_in203), .data_in204(_kanwa_x_data_in204), .data_in205(_kanwa_x_data_in205), .data_in206(_kanwa_x_data_in206), .data_in207(_kanwa_x_data_in207), .data_in208(_kanwa_x_data_in208), .data_in209(_kanwa_x_data_in209), .data_in210(_kanwa_x_data_in210), .data_in211(_kanwa_x_data_in211), .data_in212(_kanwa_x_data_in212), .data_in213(_kanwa_x_data_in213), .data_in214(_kanwa_x_data_in214), .data_in215(_kanwa_x_data_in215), .data_in216(_kanwa_x_data_in216), .data_in217(_kanwa_x_data_in217), .data_in218(_kanwa_x_data_in218), .data_in219(_kanwa_x_data_in219), .data_in220(_kanwa_x_data_in220), .data_in221(_kanwa_x_data_in221), .data_in222(_kanwa_x_data_in222), .data_in225(_kanwa_x_data_in225), .data_in226(_kanwa_x_data_in226), .data_in227(_kanwa_x_data_in227), .data_in228(_kanwa_x_data_in228), .data_in229(_kanwa_x_data_in229), .data_in230(_kanwa_x_data_in230), .data_in231(_kanwa_x_data_in231), .data_in232(_kanwa_x_data_in232), .data_in233(_kanwa_x_data_in233), .data_in234(_kanwa_x_data_in234), .data_in235(_kanwa_x_data_in235), .data_in236(_kanwa_x_data_in236), .data_in237(_kanwa_x_data_in237), .data_in238(_kanwa_x_data_in238), .data_in239(_kanwa_x_data_in239), .data_in240(_kanwa_x_data_in240), .data_in241(_kanwa_x_data_in241), .data_in242(_kanwa_x_data_in242), .data_in243(_kanwa_x_data_in243), .data_in244(_kanwa_x_data_in244), .data_in245(_kanwa_x_data_in245), .data_in246(_kanwa_x_data_in246), .data_in247(_kanwa_x_data_in247), .data_in248(_kanwa_x_data_in248), .data_in249(_kanwa_x_data_in249), .data_in250(_kanwa_x_data_in250), .data_in251(_kanwa_x_data_in251), .data_in252(_kanwa_x_data_in252), .data_in253(_kanwa_x_data_in253), .data_in254(_kanwa_x_data_in254), .data_in257(_kanwa_x_data_in257), .data_in258(_kanwa_x_data_in258), .data_in259(_kanwa_x_data_in259), .data_in260(_kanwa_x_data_in260), .data_in261(_kanwa_x_data_in261), .data_in262(_kanwa_x_data_in262), .data_in263(_kanwa_x_data_in263), .data_in264(_kanwa_x_data_in264), .data_in265(_kanwa_x_data_in265), .data_in266(_kanwa_x_data_in266), .data_in267(_kanwa_x_data_in267), .data_in268(_kanwa_x_data_in268), .data_in269(_kanwa_x_data_in269), .data_in270(_kanwa_x_data_in270), .data_in271(_kanwa_x_data_in271), .data_in272(_kanwa_x_data_in272), .data_in273(_kanwa_x_data_in273), .data_in274(_kanwa_x_data_in274), .data_in275(_kanwa_x_data_in275), .data_in276(_kanwa_x_data_in276), .data_in277(_kanwa_x_data_in277), .data_in278(_kanwa_x_data_in278), .data_in279(_kanwa_x_data_in279), .data_in280(_kanwa_x_data_in280), .data_in281(_kanwa_x_data_in281), .data_in282(_kanwa_x_data_in282), .data_in283(_kanwa_x_data_in283), .data_in284(_kanwa_x_data_in284), .data_in285(_kanwa_x_data_in285), .data_in286(_kanwa_x_data_in286), .data_in289(_kanwa_x_data_in289), .data_in290(_kanwa_x_data_in290), .data_in291(_kanwa_x_data_in291), .data_in292(_kanwa_x_data_in292), .data_in293(_kanwa_x_data_in293), .data_in294(_kanwa_x_data_in294), .data_in295(_kanwa_x_data_in295), .data_in296(_kanwa_x_data_in296), .data_in297(_kanwa_x_data_in297), .data_in298(_kanwa_x_data_in298), .data_in299(_kanwa_x_data_in299), .data_in300(_kanwa_x_data_in300), .data_in301(_kanwa_x_data_in301), .data_in302(_kanwa_x_data_in302), .data_in303(_kanwa_x_data_in303), .data_in304(_kanwa_x_data_in304), .data_in305(_kanwa_x_data_in305), .data_in306(_kanwa_x_data_in306), .data_in307(_kanwa_x_data_in307), .data_in308(_kanwa_x_data_in308), .data_in309(_kanwa_x_data_in309), .data_in310(_kanwa_x_data_in310), .data_in311(_kanwa_x_data_in311), .data_in312(_kanwa_x_data_in312), .data_in313(_kanwa_x_data_in313), .data_in314(_kanwa_x_data_in314), .data_in315(_kanwa_x_data_in315), .data_in316(_kanwa_x_data_in316), .data_in317(_kanwa_x_data_in317), .data_in318(_kanwa_x_data_in318), .data_in321(_kanwa_x_data_in321), .data_in322(_kanwa_x_data_in322), .data_in323(_kanwa_x_data_in323), .data_in324(_kanwa_x_data_in324), .data_in325(_kanwa_x_data_in325), .data_in326(_kanwa_x_data_in326), .data_in327(_kanwa_x_data_in327), .data_in328(_kanwa_x_data_in328), .data_in329(_kanwa_x_data_in329), .data_in330(_kanwa_x_data_in330), .data_in331(_kanwa_x_data_in331), .data_in332(_kanwa_x_data_in332), .data_in333(_kanwa_x_data_in333), .data_in334(_kanwa_x_data_in334), .data_in335(_kanwa_x_data_in335), .data_in336(_kanwa_x_data_in336), .data_in337(_kanwa_x_data_in337), .data_in338(_kanwa_x_data_in338), .data_in339(_kanwa_x_data_in339), .data_in340(_kanwa_x_data_in340), .data_in341(_kanwa_x_data_in341), .data_in342(_kanwa_x_data_in342), .data_in343(_kanwa_x_data_in343), .data_in344(_kanwa_x_data_in344), .data_in345(_kanwa_x_data_in345), .data_in346(_kanwa_x_data_in346), .data_in347(_kanwa_x_data_in347), .data_in348(_kanwa_x_data_in348), .data_in349(_kanwa_x_data_in349), .data_in350(_kanwa_x_data_in350), .data_in353(_kanwa_x_data_in353), .data_in354(_kanwa_x_data_in354), .data_in355(_kanwa_x_data_in355), .data_in356(_kanwa_x_data_in356), .data_in357(_kanwa_x_data_in357), .data_in358(_kanwa_x_data_in358), .data_in359(_kanwa_x_data_in359), .data_in360(_kanwa_x_data_in360), .data_in361(_kanwa_x_data_in361), .data_in362(_kanwa_x_data_in362), .data_in363(_kanwa_x_data_in363), .data_in364(_kanwa_x_data_in364), .data_in365(_kanwa_x_data_in365), .data_in366(_kanwa_x_data_in366), .data_in367(_kanwa_x_data_in367), .data_in368(_kanwa_x_data_in368), .data_in369(_kanwa_x_data_in369), .data_in370(_kanwa_x_data_in370), .data_in371(_kanwa_x_data_in371), .data_in372(_kanwa_x_data_in372), .data_in373(_kanwa_x_data_in373), .data_in374(_kanwa_x_data_in374), .data_in375(_kanwa_x_data_in375), .data_in376(_kanwa_x_data_in376), .data_in377(_kanwa_x_data_in377), .data_in378(_kanwa_x_data_in378), .data_in379(_kanwa_x_data_in379), .data_in380(_kanwa_x_data_in380), .data_in381(_kanwa_x_data_in381), .data_in382(_kanwa_x_data_in382), .data_in385(_kanwa_x_data_in385), .data_in386(_kanwa_x_data_in386), .data_in387(_kanwa_x_data_in387), .data_in388(_kanwa_x_data_in388), .data_in389(_kanwa_x_data_in389), .data_in390(_kanwa_x_data_in390), .data_in391(_kanwa_x_data_in391), .data_in392(_kanwa_x_data_in392), .data_in393(_kanwa_x_data_in393), .data_in394(_kanwa_x_data_in394), .data_in395(_kanwa_x_data_in395), .data_in396(_kanwa_x_data_in396), .data_in397(_kanwa_x_data_in397), .data_in398(_kanwa_x_data_in398), .data_in399(_kanwa_x_data_in399), .data_in400(_kanwa_x_data_in400), .data_in401(_kanwa_x_data_in401), .data_in402(_kanwa_x_data_in402), .data_in403(_kanwa_x_data_in403), .data_in404(_kanwa_x_data_in404), .data_in405(_kanwa_x_data_in405), .data_in406(_kanwa_x_data_in406), .data_in407(_kanwa_x_data_in407), .data_in408(_kanwa_x_data_in408), .data_in409(_kanwa_x_data_in409), .data_in410(_kanwa_x_data_in410), .data_in411(_kanwa_x_data_in411), .data_in412(_kanwa_x_data_in412), .data_in413(_kanwa_x_data_in413), .data_in414(_kanwa_x_data_in414), .data_in417(_kanwa_x_data_in417), .data_in418(_kanwa_x_data_in418), .data_in419(_kanwa_x_data_in419), .data_in420(_kanwa_x_data_in420), .data_in421(_kanwa_x_data_in421), .data_in422(_kanwa_x_data_in422), .data_in423(_kanwa_x_data_in423), .data_in424(_kanwa_x_data_in424), .data_in425(_kanwa_x_data_in425), .data_in426(_kanwa_x_data_in426), .data_in427(_kanwa_x_data_in427), .data_in428(_kanwa_x_data_in428), .data_in429(_kanwa_x_data_in429), .data_in430(_kanwa_x_data_in430), .data_in431(_kanwa_x_data_in431), .data_in432(_kanwa_x_data_in432), .data_in433(_kanwa_x_data_in433), .data_in434(_kanwa_x_data_in434), .data_in435(_kanwa_x_data_in435), .data_in436(_kanwa_x_data_in436), .data_in437(_kanwa_x_data_in437), .data_in438(_kanwa_x_data_in438), .data_in439(_kanwa_x_data_in439), .data_in440(_kanwa_x_data_in440), .data_in441(_kanwa_x_data_in441), .data_in442(_kanwa_x_data_in442), .data_in443(_kanwa_x_data_in443), .data_in444(_kanwa_x_data_in444), .data_in445(_kanwa_x_data_in445), .data_in446(_kanwa_x_data_in446), .data_in449(_kanwa_x_data_in449), .data_in450(_kanwa_x_data_in450), .data_in451(_kanwa_x_data_in451), .data_in452(_kanwa_x_data_in452), .data_in453(_kanwa_x_data_in453), .data_in454(_kanwa_x_data_in454), .data_in455(_kanwa_x_data_in455), .data_in456(_kanwa_x_data_in456), .data_in457(_kanwa_x_data_in457), .data_in458(_kanwa_x_data_in458), .data_in459(_kanwa_x_data_in459), .data_in460(_kanwa_x_data_in460), .data_in461(_kanwa_x_data_in461), .data_in462(_kanwa_x_data_in462), .data_in463(_kanwa_x_data_in463), .data_in464(_kanwa_x_data_in464), .data_in465(_kanwa_x_data_in465), .data_in466(_kanwa_x_data_in466), .data_in467(_kanwa_x_data_in467), .data_in468(_kanwa_x_data_in468), .data_in469(_kanwa_x_data_in469), .data_in470(_kanwa_x_data_in470), .data_in471(_kanwa_x_data_in471), .data_in472(_kanwa_x_data_in472), .data_in473(_kanwa_x_data_in473), .data_in474(_kanwa_x_data_in474), .data_in475(_kanwa_x_data_in475), .data_in476(_kanwa_x_data_in476), .data_in477(_kanwa_x_data_in477), .data_in478(_kanwa_x_data_in478), .start(_kanwa_x_start), .goal(_kanwa_x_goal));
seach seachx (.m_clock(m_clock), .p_reset( p_reset), .out_data(_seachx_out_data), .out_do(_seachx_out_do), .in_do(_seachx_in_do), .startplot(_seachx_startplot), .goalplot(_seachx_goalplot), .data_out33(_seachx_data_out33), .data_out34(_seachx_data_out34), .data_out35(_seachx_data_out35), .data_out36(_seachx_data_out36), .data_out37(_seachx_data_out37), .data_out38(_seachx_data_out38), .data_out39(_seachx_data_out39), .data_out40(_seachx_data_out40), .data_out41(_seachx_data_out41), .data_out42(_seachx_data_out42), .data_out43(_seachx_data_out43), .data_out44(_seachx_data_out44), .data_out45(_seachx_data_out45), .data_out46(_seachx_data_out46), .data_out47(_seachx_data_out47), .data_out48(_seachx_data_out48), .data_out49(_seachx_data_out49), .data_out50(_seachx_data_out50), .data_out51(_seachx_data_out51), .data_out52(_seachx_data_out52), .data_out53(_seachx_data_out53), .data_out54(_seachx_data_out54), .data_out55(_seachx_data_out55), .data_out56(_seachx_data_out56), .data_out57(_seachx_data_out57), .data_out58(_seachx_data_out58), .data_out59(_seachx_data_out59), .data_out60(_seachx_data_out60), .data_out61(_seachx_data_out61), .data_out62(_seachx_data_out62), .data_out65(_seachx_data_out65), .data_out66(_seachx_data_out66), .data_out67(_seachx_data_out67), .data_out68(_seachx_data_out68), .data_out69(_seachx_data_out69), .data_out70(_seachx_data_out70), .data_out71(_seachx_data_out71), .data_out72(_seachx_data_out72), .data_out73(_seachx_data_out73), .data_out74(_seachx_data_out74), .data_out75(_seachx_data_out75), .data_out76(_seachx_data_out76), .data_out77(_seachx_data_out77), .data_out78(_seachx_data_out78), .data_out79(_seachx_data_out79), .data_out80(_seachx_data_out80), .data_out81(_seachx_data_out81), .data_out82(_seachx_data_out82), .data_out83(_seachx_data_out83), .data_out84(_seachx_data_out84), .data_out85(_seachx_data_out85), .data_out86(_seachx_data_out86), .data_out87(_seachx_data_out87), .data_out88(_seachx_data_out88), .data_out89(_seachx_data_out89), .data_out90(_seachx_data_out90), .data_out91(_seachx_data_out91), .data_out92(_seachx_data_out92), .data_out93(_seachx_data_out93), .data_out94(_seachx_data_out94), .data_out97(_seachx_data_out97), .data_out98(_seachx_data_out98), .data_out99(_seachx_data_out99), .data_out100(_seachx_data_out100), .data_out101(_seachx_data_out101), .data_out102(_seachx_data_out102), .data_out103(_seachx_data_out103), .data_out104(_seachx_data_out104), .data_out105(_seachx_data_out105), .data_out106(_seachx_data_out106), .data_out107(_seachx_data_out107), .data_out108(_seachx_data_out108), .data_out109(_seachx_data_out109), .data_out110(_seachx_data_out110), .data_out111(_seachx_data_out111), .data_out112(_seachx_data_out112), .data_out113(_seachx_data_out113), .data_out114(_seachx_data_out114), .data_out115(_seachx_data_out115), .data_out116(_seachx_data_out116), .data_out117(_seachx_data_out117), .data_out118(_seachx_data_out118), .data_out119(_seachx_data_out119), .data_out120(_seachx_data_out120), .data_out121(_seachx_data_out121), .data_out122(_seachx_data_out122), .data_out123(_seachx_data_out123), .data_out124(_seachx_data_out124), .data_out125(_seachx_data_out125), .data_out126(_seachx_data_out126), .data_out129(_seachx_data_out129), .data_out130(_seachx_data_out130), .data_out131(_seachx_data_out131), .data_out132(_seachx_data_out132), .data_out133(_seachx_data_out133), .data_out134(_seachx_data_out134), .data_out135(_seachx_data_out135), .data_out136(_seachx_data_out136), .data_out137(_seachx_data_out137), .data_out138(_seachx_data_out138), .data_out139(_seachx_data_out139), .data_out140(_seachx_data_out140), .data_out141(_seachx_data_out141), .data_out142(_seachx_data_out142), .data_out143(_seachx_data_out143), .data_out144(_seachx_data_out144), .data_out145(_seachx_data_out145), .data_out146(_seachx_data_out146), .data_out147(_seachx_data_out147), .data_out148(_seachx_data_out148), .data_out149(_seachx_data_out149), .data_out150(_seachx_data_out150), .data_out151(_seachx_data_out151), .data_out152(_seachx_data_out152), .data_out153(_seachx_data_out153), .data_out154(_seachx_data_out154), .data_out155(_seachx_data_out155), .data_out156(_seachx_data_out156), .data_out157(_seachx_data_out157), .data_out158(_seachx_data_out158), .data_out161(_seachx_data_out161), .data_out162(_seachx_data_out162), .data_out163(_seachx_data_out163), .data_out164(_seachx_data_out164), .data_out165(_seachx_data_out165), .data_out166(_seachx_data_out166), .data_out167(_seachx_data_out167), .data_out168(_seachx_data_out168), .data_out169(_seachx_data_out169), .data_out170(_seachx_data_out170), .data_out171(_seachx_data_out171), .data_out172(_seachx_data_out172), .data_out173(_seachx_data_out173), .data_out174(_seachx_data_out174), .data_out175(_seachx_data_out175), .data_out176(_seachx_data_out176), .data_out177(_seachx_data_out177), .data_out178(_seachx_data_out178), .data_out179(_seachx_data_out179), .data_out180(_seachx_data_out180), .data_out181(_seachx_data_out181), .data_out182(_seachx_data_out182), .data_out183(_seachx_data_out183), .data_out184(_seachx_data_out184), .data_out185(_seachx_data_out185), .data_out186(_seachx_data_out186), .data_out187(_seachx_data_out187), .data_out188(_seachx_data_out188), .data_out189(_seachx_data_out189), .data_out190(_seachx_data_out190), .data_out193(_seachx_data_out193), .data_out194(_seachx_data_out194), .data_out195(_seachx_data_out195), .data_out196(_seachx_data_out196), .data_out197(_seachx_data_out197), .data_out198(_seachx_data_out198), .data_out199(_seachx_data_out199), .data_out200(_seachx_data_out200), .data_out201(_seachx_data_out201), .data_out202(_seachx_data_out202), .data_out203(_seachx_data_out203), .data_out204(_seachx_data_out204), .data_out205(_seachx_data_out205), .data_out206(_seachx_data_out206), .data_out207(_seachx_data_out207), .data_out208(_seachx_data_out208), .data_out209(_seachx_data_out209), .data_out210(_seachx_data_out210), .data_out211(_seachx_data_out211), .data_out212(_seachx_data_out212), .data_out213(_seachx_data_out213), .data_out214(_seachx_data_out214), .data_out215(_seachx_data_out215), .data_out216(_seachx_data_out216), .data_out217(_seachx_data_out217), .data_out218(_seachx_data_out218), .data_out219(_seachx_data_out219), .data_out220(_seachx_data_out220), .data_out221(_seachx_data_out221), .data_out222(_seachx_data_out222), .data_out225(_seachx_data_out225), .data_out226(_seachx_data_out226), .data_out227(_seachx_data_out227), .data_out228(_seachx_data_out228), .data_out229(_seachx_data_out229), .data_out230(_seachx_data_out230), .data_out231(_seachx_data_out231), .data_out232(_seachx_data_out232), .data_out233(_seachx_data_out233), .data_out234(_seachx_data_out234), .data_out235(_seachx_data_out235), .data_out236(_seachx_data_out236), .data_out237(_seachx_data_out237), .data_out238(_seachx_data_out238), .data_out239(_seachx_data_out239), .data_out240(_seachx_data_out240), .data_out241(_seachx_data_out241), .data_out242(_seachx_data_out242), .data_out243(_seachx_data_out243), .data_out244(_seachx_data_out244), .data_out245(_seachx_data_out245), .data_out246(_seachx_data_out246), .data_out247(_seachx_data_out247), .data_out248(_seachx_data_out248), .data_out249(_seachx_data_out249), .data_out250(_seachx_data_out250), .data_out251(_seachx_data_out251), .data_out252(_seachx_data_out252), .data_out253(_seachx_data_out253), .data_out254(_seachx_data_out254), .data_out257(_seachx_data_out257), .data_out258(_seachx_data_out258), .data_out259(_seachx_data_out259), .data_out260(_seachx_data_out260), .data_out261(_seachx_data_out261), .data_out262(_seachx_data_out262), .data_out263(_seachx_data_out263), .data_out264(_seachx_data_out264), .data_out265(_seachx_data_out265), .data_out266(_seachx_data_out266), .data_out267(_seachx_data_out267), .data_out268(_seachx_data_out268), .data_out269(_seachx_data_out269), .data_out270(_seachx_data_out270), .data_out271(_seachx_data_out271), .data_out272(_seachx_data_out272), .data_out273(_seachx_data_out273), .data_out274(_seachx_data_out274), .data_out275(_seachx_data_out275), .data_out276(_seachx_data_out276), .data_out277(_seachx_data_out277), .data_out278(_seachx_data_out278), .data_out279(_seachx_data_out279), .data_out280(_seachx_data_out280), .data_out281(_seachx_data_out281), .data_out282(_seachx_data_out282), .data_out283(_seachx_data_out283), .data_out284(_seachx_data_out284), .data_out285(_seachx_data_out285), .data_out286(_seachx_data_out286), .data_out289(_seachx_data_out289), .data_out290(_seachx_data_out290), .data_out291(_seachx_data_out291), .data_out292(_seachx_data_out292), .data_out293(_seachx_data_out293), .data_out294(_seachx_data_out294), .data_out295(_seachx_data_out295), .data_out296(_seachx_data_out296), .data_out297(_seachx_data_out297), .data_out298(_seachx_data_out298), .data_out299(_seachx_data_out299), .data_out300(_seachx_data_out300), .data_out301(_seachx_data_out301), .data_out302(_seachx_data_out302), .data_out303(_seachx_data_out303), .data_out304(_seachx_data_out304), .data_out305(_seachx_data_out305), .data_out306(_seachx_data_out306), .data_out307(_seachx_data_out307), .data_out308(_seachx_data_out308), .data_out309(_seachx_data_out309), .data_out310(_seachx_data_out310), .data_out311(_seachx_data_out311), .data_out312(_seachx_data_out312), .data_out313(_seachx_data_out313), .data_out314(_seachx_data_out314), .data_out315(_seachx_data_out315), .data_out316(_seachx_data_out316), .data_out317(_seachx_data_out317), .data_out318(_seachx_data_out318), .data_out321(_seachx_data_out321), .data_out322(_seachx_data_out322), .data_out323(_seachx_data_out323), .data_out324(_seachx_data_out324), .data_out325(_seachx_data_out325), .data_out326(_seachx_data_out326), .data_out327(_seachx_data_out327), .data_out328(_seachx_data_out328), .data_out329(_seachx_data_out329), .data_out330(_seachx_data_out330), .data_out331(_seachx_data_out331), .data_out332(_seachx_data_out332), .data_out333(_seachx_data_out333), .data_out334(_seachx_data_out334), .data_out335(_seachx_data_out335), .data_out336(_seachx_data_out336), .data_out337(_seachx_data_out337), .data_out338(_seachx_data_out338), .data_out339(_seachx_data_out339), .data_out340(_seachx_data_out340), .data_out341(_seachx_data_out341), .data_out342(_seachx_data_out342), .data_out343(_seachx_data_out343), .data_out344(_seachx_data_out344), .data_out345(_seachx_data_out345), .data_out346(_seachx_data_out346), .data_out347(_seachx_data_out347), .data_out348(_seachx_data_out348), .data_out349(_seachx_data_out349), .data_out350(_seachx_data_out350), .data_out353(_seachx_data_out353), .data_out354(_seachx_data_out354), .data_out355(_seachx_data_out355), .data_out356(_seachx_data_out356), .data_out357(_seachx_data_out357), .data_out358(_seachx_data_out358), .data_out359(_seachx_data_out359), .data_out360(_seachx_data_out360), .data_out361(_seachx_data_out361), .data_out362(_seachx_data_out362), .data_out363(_seachx_data_out363), .data_out364(_seachx_data_out364), .data_out365(_seachx_data_out365), .data_out366(_seachx_data_out366), .data_out367(_seachx_data_out367), .data_out368(_seachx_data_out368), .data_out369(_seachx_data_out369), .data_out370(_seachx_data_out370), .data_out371(_seachx_data_out371), .data_out372(_seachx_data_out372), .data_out373(_seachx_data_out373), .data_out374(_seachx_data_out374), .data_out375(_seachx_data_out375), .data_out376(_seachx_data_out376), .data_out377(_seachx_data_out377), .data_out378(_seachx_data_out378), .data_out379(_seachx_data_out379), .data_out380(_seachx_data_out380), .data_out381(_seachx_data_out381), .data_out382(_seachx_data_out382), .data_out385(_seachx_data_out385), .data_out386(_seachx_data_out386), .data_out387(_seachx_data_out387), .data_out388(_seachx_data_out388), .data_out389(_seachx_data_out389), .data_out390(_seachx_data_out390), .data_out391(_seachx_data_out391), .data_out392(_seachx_data_out392), .data_out393(_seachx_data_out393), .data_out394(_seachx_data_out394), .data_out395(_seachx_data_out395), .data_out396(_seachx_data_out396), .data_out397(_seachx_data_out397), .data_out398(_seachx_data_out398), .data_out399(_seachx_data_out399), .data_out400(_seachx_data_out400), .data_out401(_seachx_data_out401), .data_out402(_seachx_data_out402), .data_out403(_seachx_data_out403), .data_out404(_seachx_data_out404), .data_out405(_seachx_data_out405), .data_out406(_seachx_data_out406), .data_out407(_seachx_data_out407), .data_out408(_seachx_data_out408), .data_out409(_seachx_data_out409), .data_out410(_seachx_data_out410), .data_out411(_seachx_data_out411), .data_out412(_seachx_data_out412), .data_out413(_seachx_data_out413), .data_out414(_seachx_data_out414), .data_out417(_seachx_data_out417), .data_out418(_seachx_data_out418), .data_out419(_seachx_data_out419), .data_out420(_seachx_data_out420), .data_out421(_seachx_data_out421), .data_out422(_seachx_data_out422), .data_out423(_seachx_data_out423), .data_out424(_seachx_data_out424), .data_out425(_seachx_data_out425), .data_out426(_seachx_data_out426), .data_out427(_seachx_data_out427), .data_out428(_seachx_data_out428), .data_out429(_seachx_data_out429), .data_out430(_seachx_data_out430), .data_out431(_seachx_data_out431), .data_out432(_seachx_data_out432), .data_out433(_seachx_data_out433), .data_out434(_seachx_data_out434), .data_out435(_seachx_data_out435), .data_out436(_seachx_data_out436), .data_out437(_seachx_data_out437), .data_out438(_seachx_data_out438), .data_out439(_seachx_data_out439), .data_out440(_seachx_data_out440), .data_out441(_seachx_data_out441), .data_out442(_seachx_data_out442), .data_out443(_seachx_data_out443), .data_out444(_seachx_data_out444), .data_out445(_seachx_data_out445), .data_out446(_seachx_data_out446), .data_out449(_seachx_data_out449), .data_out450(_seachx_data_out450), .data_out451(_seachx_data_out451), .data_out452(_seachx_data_out452), .data_out453(_seachx_data_out453), .data_out454(_seachx_data_out454), .data_out455(_seachx_data_out455), .data_out456(_seachx_data_out456), .data_out457(_seachx_data_out457), .data_out458(_seachx_data_out458), .data_out459(_seachx_data_out459), .data_out460(_seachx_data_out460), .data_out461(_seachx_data_out461), .data_out462(_seachx_data_out462), .data_out463(_seachx_data_out463), .data_out464(_seachx_data_out464), .data_out465(_seachx_data_out465), .data_out466(_seachx_data_out466), .data_out467(_seachx_data_out467), .data_out468(_seachx_data_out468), .data_out469(_seachx_data_out469), .data_out470(_seachx_data_out470), .data_out471(_seachx_data_out471), .data_out472(_seachx_data_out472), .data_out473(_seachx_data_out473), .data_out474(_seachx_data_out474), .data_out475(_seachx_data_out475), .data_out476(_seachx_data_out476), .data_out477(_seachx_data_out477), .data_out478(_seachx_data_out478), .data_in33(_seachx_data_in33), .data_in34(_seachx_data_in34), .data_in35(_seachx_data_in35), .data_in36(_seachx_data_in36), .data_in37(_seachx_data_in37), .data_in38(_seachx_data_in38), .data_in39(_seachx_data_in39), .data_in40(_seachx_data_in40), .data_in41(_seachx_data_in41), .data_in42(_seachx_data_in42), .data_in43(_seachx_data_in43), .data_in44(_seachx_data_in44), .data_in45(_seachx_data_in45), .data_in46(_seachx_data_in46), .data_in47(_seachx_data_in47), .data_in48(_seachx_data_in48), .data_in49(_seachx_data_in49), .data_in50(_seachx_data_in50), .data_in51(_seachx_data_in51), .data_in52(_seachx_data_in52), .data_in53(_seachx_data_in53), .data_in54(_seachx_data_in54), .data_in55(_seachx_data_in55), .data_in56(_seachx_data_in56), .data_in57(_seachx_data_in57), .data_in58(_seachx_data_in58), .data_in59(_seachx_data_in59), .data_in60(_seachx_data_in60), .data_in61(_seachx_data_in61), .data_in62(_seachx_data_in62), .data_in65(_seachx_data_in65), .data_in66(_seachx_data_in66), .data_in67(_seachx_data_in67), .data_in68(_seachx_data_in68), .data_in69(_seachx_data_in69), .data_in70(_seachx_data_in70), .data_in71(_seachx_data_in71), .data_in72(_seachx_data_in72), .data_in73(_seachx_data_in73), .data_in74(_seachx_data_in74), .data_in75(_seachx_data_in75), .data_in76(_seachx_data_in76), .data_in77(_seachx_data_in77), .data_in78(_seachx_data_in78), .data_in79(_seachx_data_in79), .data_in80(_seachx_data_in80), .data_in81(_seachx_data_in81), .data_in82(_seachx_data_in82), .data_in83(_seachx_data_in83), .data_in84(_seachx_data_in84), .data_in85(_seachx_data_in85), .data_in86(_seachx_data_in86), .data_in87(_seachx_data_in87), .data_in88(_seachx_data_in88), .data_in89(_seachx_data_in89), .data_in90(_seachx_data_in90), .data_in91(_seachx_data_in91), .data_in92(_seachx_data_in92), .data_in93(_seachx_data_in93), .data_in94(_seachx_data_in94), .data_in97(_seachx_data_in97), .data_in98(_seachx_data_in98), .data_in99(_seachx_data_in99), .data_in100(_seachx_data_in100), .data_in101(_seachx_data_in101), .data_in102(_seachx_data_in102), .data_in103(_seachx_data_in103), .data_in104(_seachx_data_in104), .data_in105(_seachx_data_in105), .data_in106(_seachx_data_in106), .data_in107(_seachx_data_in107), .data_in108(_seachx_data_in108), .data_in109(_seachx_data_in109), .data_in110(_seachx_data_in110), .data_in111(_seachx_data_in111), .data_in112(_seachx_data_in112), .data_in113(_seachx_data_in113), .data_in114(_seachx_data_in114), .data_in115(_seachx_data_in115), .data_in116(_seachx_data_in116), .data_in117(_seachx_data_in117), .data_in118(_seachx_data_in118), .data_in119(_seachx_data_in119), .data_in120(_seachx_data_in120), .data_in121(_seachx_data_in121), .data_in122(_seachx_data_in122), .data_in123(_seachx_data_in123), .data_in124(_seachx_data_in124), .data_in125(_seachx_data_in125), .data_in126(_seachx_data_in126), .data_in129(_seachx_data_in129), .data_in130(_seachx_data_in130), .data_in131(_seachx_data_in131), .data_in132(_seachx_data_in132), .data_in133(_seachx_data_in133), .data_in134(_seachx_data_in134), .data_in135(_seachx_data_in135), .data_in136(_seachx_data_in136), .data_in137(_seachx_data_in137), .data_in138(_seachx_data_in138), .data_in139(_seachx_data_in139), .data_in140(_seachx_data_in140), .data_in141(_seachx_data_in141), .data_in142(_seachx_data_in142), .data_in143(_seachx_data_in143), .data_in144(_seachx_data_in144), .data_in145(_seachx_data_in145), .data_in146(_seachx_data_in146), .data_in147(_seachx_data_in147), .data_in148(_seachx_data_in148), .data_in149(_seachx_data_in149), .data_in150(_seachx_data_in150), .data_in151(_seachx_data_in151), .data_in152(_seachx_data_in152), .data_in153(_seachx_data_in153), .data_in154(_seachx_data_in154), .data_in155(_seachx_data_in155), .data_in156(_seachx_data_in156), .data_in157(_seachx_data_in157), .data_in158(_seachx_data_in158), .data_in161(_seachx_data_in161), .data_in162(_seachx_data_in162), .data_in163(_seachx_data_in163), .data_in164(_seachx_data_in164), .data_in165(_seachx_data_in165), .data_in166(_seachx_data_in166), .data_in167(_seachx_data_in167), .data_in168(_seachx_data_in168), .data_in169(_seachx_data_in169), .data_in170(_seachx_data_in170), .data_in171(_seachx_data_in171), .data_in172(_seachx_data_in172), .data_in173(_seachx_data_in173), .data_in174(_seachx_data_in174), .data_in175(_seachx_data_in175), .data_in176(_seachx_data_in176), .data_in177(_seachx_data_in177), .data_in178(_seachx_data_in178), .data_in179(_seachx_data_in179), .data_in180(_seachx_data_in180), .data_in181(_seachx_data_in181), .data_in182(_seachx_data_in182), .data_in183(_seachx_data_in183), .data_in184(_seachx_data_in184), .data_in185(_seachx_data_in185), .data_in186(_seachx_data_in186), .data_in187(_seachx_data_in187), .data_in188(_seachx_data_in188), .data_in189(_seachx_data_in189), .data_in190(_seachx_data_in190), .data_in193(_seachx_data_in193), .data_in194(_seachx_data_in194), .data_in195(_seachx_data_in195), .data_in196(_seachx_data_in196), .data_in197(_seachx_data_in197), .data_in198(_seachx_data_in198), .data_in199(_seachx_data_in199), .data_in200(_seachx_data_in200), .data_in201(_seachx_data_in201), .data_in202(_seachx_data_in202), .data_in203(_seachx_data_in203), .data_in204(_seachx_data_in204), .data_in205(_seachx_data_in205), .data_in206(_seachx_data_in206), .data_in207(_seachx_data_in207), .data_in208(_seachx_data_in208), .data_in209(_seachx_data_in209), .data_in210(_seachx_data_in210), .data_in211(_seachx_data_in211), .data_in212(_seachx_data_in212), .data_in213(_seachx_data_in213), .data_in214(_seachx_data_in214), .data_in215(_seachx_data_in215), .data_in216(_seachx_data_in216), .data_in217(_seachx_data_in217), .data_in218(_seachx_data_in218), .data_in219(_seachx_data_in219), .data_in220(_seachx_data_in220), .data_in221(_seachx_data_in221), .data_in222(_seachx_data_in222), .data_in225(_seachx_data_in225), .data_in226(_seachx_data_in226), .data_in227(_seachx_data_in227), .data_in228(_seachx_data_in228), .data_in229(_seachx_data_in229), .data_in230(_seachx_data_in230), .data_in231(_seachx_data_in231), .data_in232(_seachx_data_in232), .data_in233(_seachx_data_in233), .data_in234(_seachx_data_in234), .data_in235(_seachx_data_in235), .data_in236(_seachx_data_in236), .data_in237(_seachx_data_in237), .data_in238(_seachx_data_in238), .data_in239(_seachx_data_in239), .data_in240(_seachx_data_in240), .data_in241(_seachx_data_in241), .data_in242(_seachx_data_in242), .data_in243(_seachx_data_in243), .data_in244(_seachx_data_in244), .data_in245(_seachx_data_in245), .data_in246(_seachx_data_in246), .data_in247(_seachx_data_in247), .data_in248(_seachx_data_in248), .data_in249(_seachx_data_in249), .data_in250(_seachx_data_in250), .data_in251(_seachx_data_in251), .data_in252(_seachx_data_in252), .data_in253(_seachx_data_in253), .data_in254(_seachx_data_in254), .data_in257(_seachx_data_in257), .data_in258(_seachx_data_in258), .data_in259(_seachx_data_in259), .data_in260(_seachx_data_in260), .data_in261(_seachx_data_in261), .data_in262(_seachx_data_in262), .data_in263(_seachx_data_in263), .data_in264(_seachx_data_in264), .data_in265(_seachx_data_in265), .data_in266(_seachx_data_in266), .data_in267(_seachx_data_in267), .data_in268(_seachx_data_in268), .data_in269(_seachx_data_in269), .data_in270(_seachx_data_in270), .data_in271(_seachx_data_in271), .data_in272(_seachx_data_in272), .data_in273(_seachx_data_in273), .data_in274(_seachx_data_in274), .data_in275(_seachx_data_in275), .data_in276(_seachx_data_in276), .data_in277(_seachx_data_in277), .data_in278(_seachx_data_in278), .data_in279(_seachx_data_in279), .data_in280(_seachx_data_in280), .data_in281(_seachx_data_in281), .data_in282(_seachx_data_in282), .data_in283(_seachx_data_in283), .data_in284(_seachx_data_in284), .data_in285(_seachx_data_in285), .data_in286(_seachx_data_in286), .data_in289(_seachx_data_in289), .data_in290(_seachx_data_in290), .data_in291(_seachx_data_in291), .data_in292(_seachx_data_in292), .data_in293(_seachx_data_in293), .data_in294(_seachx_data_in294), .data_in295(_seachx_data_in295), .data_in296(_seachx_data_in296), .data_in297(_seachx_data_in297), .data_in298(_seachx_data_in298), .data_in299(_seachx_data_in299), .data_in300(_seachx_data_in300), .data_in301(_seachx_data_in301), .data_in302(_seachx_data_in302), .data_in303(_seachx_data_in303), .data_in304(_seachx_data_in304), .data_in305(_seachx_data_in305), .data_in306(_seachx_data_in306), .data_in307(_seachx_data_in307), .data_in308(_seachx_data_in308), .data_in309(_seachx_data_in309), .data_in310(_seachx_data_in310), .data_in311(_seachx_data_in311), .data_in312(_seachx_data_in312), .data_in313(_seachx_data_in313), .data_in314(_seachx_data_in314), .data_in315(_seachx_data_in315), .data_in316(_seachx_data_in316), .data_in317(_seachx_data_in317), .data_in318(_seachx_data_in318), .data_in321(_seachx_data_in321), .data_in322(_seachx_data_in322), .data_in323(_seachx_data_in323), .data_in324(_seachx_data_in324), .data_in325(_seachx_data_in325), .data_in326(_seachx_data_in326), .data_in327(_seachx_data_in327), .data_in328(_seachx_data_in328), .data_in329(_seachx_data_in329), .data_in330(_seachx_data_in330), .data_in331(_seachx_data_in331), .data_in332(_seachx_data_in332), .data_in333(_seachx_data_in333), .data_in334(_seachx_data_in334), .data_in335(_seachx_data_in335), .data_in336(_seachx_data_in336), .data_in337(_seachx_data_in337), .data_in338(_seachx_data_in338), .data_in339(_seachx_data_in339), .data_in340(_seachx_data_in340), .data_in341(_seachx_data_in341), .data_in342(_seachx_data_in342), .data_in343(_seachx_data_in343), .data_in344(_seachx_data_in344), .data_in345(_seachx_data_in345), .data_in346(_seachx_data_in346), .data_in347(_seachx_data_in347), .data_in348(_seachx_data_in348), .data_in349(_seachx_data_in349), .data_in350(_seachx_data_in350), .data_in353(_seachx_data_in353), .data_in354(_seachx_data_in354), .data_in355(_seachx_data_in355), .data_in356(_seachx_data_in356), .data_in357(_seachx_data_in357), .data_in358(_seachx_data_in358), .data_in359(_seachx_data_in359), .data_in360(_seachx_data_in360), .data_in361(_seachx_data_in361), .data_in362(_seachx_data_in362), .data_in363(_seachx_data_in363), .data_in364(_seachx_data_in364), .data_in365(_seachx_data_in365), .data_in366(_seachx_data_in366), .data_in367(_seachx_data_in367), .data_in368(_seachx_data_in368), .data_in369(_seachx_data_in369), .data_in370(_seachx_data_in370), .data_in371(_seachx_data_in371), .data_in372(_seachx_data_in372), .data_in373(_seachx_data_in373), .data_in374(_seachx_data_in374), .data_in375(_seachx_data_in375), .data_in376(_seachx_data_in376), .data_in377(_seachx_data_in377), .data_in378(_seachx_data_in378), .data_in379(_seachx_data_in379), .data_in380(_seachx_data_in380), .data_in381(_seachx_data_in381), .data_in382(_seachx_data_in382), .data_in385(_seachx_data_in385), .data_in386(_seachx_data_in386), .data_in387(_seachx_data_in387), .data_in388(_seachx_data_in388), .data_in389(_seachx_data_in389), .data_in390(_seachx_data_in390), .data_in391(_seachx_data_in391), .data_in392(_seachx_data_in392), .data_in393(_seachx_data_in393), .data_in394(_seachx_data_in394), .data_in395(_seachx_data_in395), .data_in396(_seachx_data_in396), .data_in397(_seachx_data_in397), .data_in398(_seachx_data_in398), .data_in399(_seachx_data_in399), .data_in400(_seachx_data_in400), .data_in401(_seachx_data_in401), .data_in402(_seachx_data_in402), .data_in403(_seachx_data_in403), .data_in404(_seachx_data_in404), .data_in405(_seachx_data_in405), .data_in406(_seachx_data_in406), .data_in407(_seachx_data_in407), .data_in408(_seachx_data_in408), .data_in409(_seachx_data_in409), .data_in410(_seachx_data_in410), .data_in411(_seachx_data_in411), .data_in412(_seachx_data_in412), .data_in413(_seachx_data_in413), .data_in414(_seachx_data_in414), .data_in417(_seachx_data_in417), .data_in418(_seachx_data_in418), .data_in419(_seachx_data_in419), .data_in420(_seachx_data_in420), .data_in421(_seachx_data_in421), .data_in422(_seachx_data_in422), .data_in423(_seachx_data_in423), .data_in424(_seachx_data_in424), .data_in425(_seachx_data_in425), .data_in426(_seachx_data_in426), .data_in427(_seachx_data_in427), .data_in428(_seachx_data_in428), .data_in429(_seachx_data_in429), .data_in430(_seachx_data_in430), .data_in431(_seachx_data_in431), .data_in432(_seachx_data_in432), .data_in433(_seachx_data_in433), .data_in434(_seachx_data_in434), .data_in435(_seachx_data_in435), .data_in436(_seachx_data_in436), .data_in437(_seachx_data_in437), .data_in438(_seachx_data_in438), .data_in439(_seachx_data_in439), .data_in440(_seachx_data_in440), .data_in441(_seachx_data_in441), .data_in442(_seachx_data_in442), .data_in443(_seachx_data_in443), .data_in444(_seachx_data_in444), .data_in445(_seachx_data_in445), .data_in446(_seachx_data_in446), .data_in449(_seachx_data_in449), .data_in450(_seachx_data_in450), .data_in451(_seachx_data_in451), .data_in452(_seachx_data_in452), .data_in453(_seachx_data_in453), .data_in454(_seachx_data_in454), .data_in455(_seachx_data_in455), .data_in456(_seachx_data_in456), .data_in457(_seachx_data_in457), .data_in458(_seachx_data_in458), .data_in459(_seachx_data_in459), .data_in460(_seachx_data_in460), .data_in461(_seachx_data_in461), .data_in462(_seachx_data_in462), .data_in463(_seachx_data_in463), .data_in464(_seachx_data_in464), .data_in465(_seachx_data_in465), .data_in466(_seachx_data_in466), .data_in467(_seachx_data_in467), .data_in468(_seachx_data_in468), .data_in469(_seachx_data_in469), .data_in470(_seachx_data_in470), .data_in471(_seachx_data_in471), .data_in472(_seachx_data_in472), .data_in473(_seachx_data_in473), .data_in474(_seachx_data_in474), .data_in475(_seachx_data_in475), .data_in476(_seachx_data_in476), .data_in477(_seachx_data_in477), .data_in478(_seachx_data_in478));

   assign  _seachx_data_in33 = map_value_arg33;
   assign  _seachx_data_in34 = map_value_arg34;
   assign  _seachx_data_in35 = map_value_arg35;
   assign  _seachx_data_in36 = map_value_arg36;
   assign  _seachx_data_in37 = map_value_arg37;
   assign  _seachx_data_in38 = map_value_arg38;
   assign  _seachx_data_in39 = map_value_arg39;
   assign  _seachx_data_in40 = map_value_arg40;
   assign  _seachx_data_in41 = map_value_arg41;
   assign  _seachx_data_in42 = map_value_arg42;
   assign  _seachx_data_in43 = map_value_arg43;
   assign  _seachx_data_in44 = map_value_arg44;
   assign  _seachx_data_in45 = map_value_arg45;
   assign  _seachx_data_in46 = map_value_arg46;
   assign  _seachx_data_in47 = map_value_arg47;
   assign  _seachx_data_in48 = map_value_arg48;
   assign  _seachx_data_in49 = map_value_arg49;
   assign  _seachx_data_in50 = map_value_arg50;
   assign  _seachx_data_in51 = map_value_arg51;
   assign  _seachx_data_in52 = map_value_arg52;
   assign  _seachx_data_in53 = map_value_arg53;
   assign  _seachx_data_in54 = map_value_arg54;
   assign  _seachx_data_in55 = map_value_arg55;
   assign  _seachx_data_in56 = map_value_arg56;
   assign  _seachx_data_in57 = map_value_arg57;
   assign  _seachx_data_in58 = map_value_arg58;
   assign  _seachx_data_in59 = map_value_arg59;
   assign  _seachx_data_in60 = map_value_arg60;
   assign  _seachx_data_in61 = map_value_arg61;
   assign  _seachx_data_in62 = map_value_arg62;
   assign  _seachx_data_in65 = map_value_arg65;
   assign  _seachx_data_in66 = map_value_arg66;
   assign  _seachx_data_in67 = map_value_arg67;
   assign  _seachx_data_in68 = map_value_arg68;
   assign  _seachx_data_in69 = map_value_arg69;
   assign  _seachx_data_in70 = map_value_arg70;
   assign  _seachx_data_in71 = map_value_arg71;
   assign  _seachx_data_in72 = map_value_arg72;
   assign  _seachx_data_in73 = map_value_arg73;
   assign  _seachx_data_in74 = map_value_arg74;
   assign  _seachx_data_in75 = map_value_arg75;
   assign  _seachx_data_in76 = map_value_arg76;
   assign  _seachx_data_in77 = map_value_arg77;
   assign  _seachx_data_in78 = map_value_arg78;
   assign  _seachx_data_in79 = map_value_arg79;
   assign  _seachx_data_in80 = map_value_arg80;
   assign  _seachx_data_in81 = map_value_arg81;
   assign  _seachx_data_in82 = map_value_arg82;
   assign  _seachx_data_in83 = map_value_arg83;
   assign  _seachx_data_in84 = map_value_arg84;
   assign  _seachx_data_in85 = map_value_arg85;
   assign  _seachx_data_in86 = map_value_arg86;
   assign  _seachx_data_in87 = map_value_arg87;
   assign  _seachx_data_in88 = map_value_arg88;
   assign  _seachx_data_in89 = map_value_arg89;
   assign  _seachx_data_in90 = map_value_arg90;
   assign  _seachx_data_in91 = map_value_arg91;
   assign  _seachx_data_in92 = map_value_arg92;
   assign  _seachx_data_in93 = map_value_arg93;
   assign  _seachx_data_in94 = map_value_arg94;
   assign  _seachx_data_in97 = map_value_arg97;
   assign  _seachx_data_in98 = map_value_arg98;
   assign  _seachx_data_in99 = map_value_arg99;
   assign  _seachx_data_in100 = map_value_arg100;
   assign  _seachx_data_in101 = map_value_arg101;
   assign  _seachx_data_in102 = map_value_arg102;
   assign  _seachx_data_in103 = map_value_arg103;
   assign  _seachx_data_in104 = map_value_arg104;
   assign  _seachx_data_in105 = map_value_arg105;
   assign  _seachx_data_in106 = map_value_arg106;
   assign  _seachx_data_in107 = map_value_arg107;
   assign  _seachx_data_in108 = map_value_arg108;
   assign  _seachx_data_in109 = map_value_arg109;
   assign  _seachx_data_in110 = map_value_arg110;
   assign  _seachx_data_in111 = map_value_arg111;
   assign  _seachx_data_in112 = map_value_arg112;
   assign  _seachx_data_in113 = map_value_arg113;
   assign  _seachx_data_in114 = map_value_arg114;
   assign  _seachx_data_in115 = map_value_arg115;
   assign  _seachx_data_in116 = map_value_arg116;
   assign  _seachx_data_in117 = map_value_arg117;
   assign  _seachx_data_in118 = map_value_arg118;
   assign  _seachx_data_in119 = map_value_arg119;
   assign  _seachx_data_in120 = map_value_arg120;
   assign  _seachx_data_in121 = map_value_arg121;
   assign  _seachx_data_in122 = map_value_arg122;
   assign  _seachx_data_in123 = map_value_arg123;
   assign  _seachx_data_in124 = map_value_arg124;
   assign  _seachx_data_in125 = map_value_arg125;
   assign  _seachx_data_in126 = map_value_arg126;
   assign  _seachx_data_in129 = map_value_arg129;
   assign  _seachx_data_in130 = map_value_arg130;
   assign  _seachx_data_in131 = map_value_arg131;
   assign  _seachx_data_in132 = map_value_arg132;
   assign  _seachx_data_in133 = map_value_arg133;
   assign  _seachx_data_in134 = map_value_arg134;
   assign  _seachx_data_in135 = map_value_arg135;
   assign  _seachx_data_in136 = map_value_arg136;
   assign  _seachx_data_in137 = map_value_arg137;
   assign  _seachx_data_in138 = map_value_arg138;
   assign  _seachx_data_in139 = map_value_arg139;
   assign  _seachx_data_in140 = map_value_arg140;
   assign  _seachx_data_in141 = map_value_arg141;
   assign  _seachx_data_in142 = map_value_arg142;
   assign  _seachx_data_in143 = map_value_arg143;
   assign  _seachx_data_in144 = map_value_arg144;
   assign  _seachx_data_in145 = map_value_arg145;
   assign  _seachx_data_in146 = map_value_arg146;
   assign  _seachx_data_in147 = map_value_arg147;
   assign  _seachx_data_in148 = map_value_arg148;
   assign  _seachx_data_in149 = map_value_arg149;
   assign  _seachx_data_in150 = map_value_arg150;
   assign  _seachx_data_in151 = map_value_arg151;
   assign  _seachx_data_in152 = map_value_arg152;
   assign  _seachx_data_in153 = map_value_arg153;
   assign  _seachx_data_in154 = map_value_arg154;
   assign  _seachx_data_in155 = map_value_arg155;
   assign  _seachx_data_in156 = map_value_arg156;
   assign  _seachx_data_in157 = map_value_arg157;
   assign  _seachx_data_in158 = map_value_arg158;
   assign  _seachx_data_in161 = map_value_arg161;
   assign  _seachx_data_in162 = map_value_arg162;
   assign  _seachx_data_in163 = map_value_arg163;
   assign  _seachx_data_in164 = map_value_arg164;
   assign  _seachx_data_in165 = map_value_arg165;
   assign  _seachx_data_in166 = map_value_arg166;
   assign  _seachx_data_in167 = map_value_arg167;
   assign  _seachx_data_in168 = map_value_arg168;
   assign  _seachx_data_in169 = map_value_arg169;
   assign  _seachx_data_in170 = map_value_arg170;
   assign  _seachx_data_in171 = map_value_arg171;
   assign  _seachx_data_in172 = map_value_arg172;
   assign  _seachx_data_in173 = map_value_arg173;
   assign  _seachx_data_in174 = map_value_arg174;
   assign  _seachx_data_in175 = map_value_arg175;
   assign  _seachx_data_in176 = map_value_arg176;
   assign  _seachx_data_in177 = map_value_arg177;
   assign  _seachx_data_in178 = map_value_arg178;
   assign  _seachx_data_in179 = map_value_arg179;
   assign  _seachx_data_in180 = map_value_arg180;
   assign  _seachx_data_in181 = map_value_arg181;
   assign  _seachx_data_in182 = map_value_arg182;
   assign  _seachx_data_in183 = map_value_arg183;
   assign  _seachx_data_in184 = map_value_arg184;
   assign  _seachx_data_in185 = map_value_arg185;
   assign  _seachx_data_in186 = map_value_arg186;
   assign  _seachx_data_in187 = map_value_arg187;
   assign  _seachx_data_in188 = map_value_arg188;
   assign  _seachx_data_in189 = map_value_arg189;
   assign  _seachx_data_in190 = map_value_arg190;
   assign  _seachx_data_in193 = map_value_arg193;
   assign  _seachx_data_in194 = map_value_arg194;
   assign  _seachx_data_in195 = map_value_arg195;
   assign  _seachx_data_in196 = map_value_arg196;
   assign  _seachx_data_in197 = map_value_arg197;
   assign  _seachx_data_in198 = map_value_arg198;
   assign  _seachx_data_in199 = map_value_arg199;
   assign  _seachx_data_in200 = map_value_arg200;
   assign  _seachx_data_in201 = map_value_arg201;
   assign  _seachx_data_in202 = map_value_arg202;
   assign  _seachx_data_in203 = map_value_arg203;
   assign  _seachx_data_in204 = map_value_arg204;
   assign  _seachx_data_in205 = map_value_arg205;
   assign  _seachx_data_in206 = map_value_arg206;
   assign  _seachx_data_in207 = map_value_arg207;
   assign  _seachx_data_in208 = map_value_arg208;
   assign  _seachx_data_in209 = map_value_arg209;
   assign  _seachx_data_in210 = map_value_arg210;
   assign  _seachx_data_in211 = map_value_arg211;
   assign  _seachx_data_in212 = map_value_arg212;
   assign  _seachx_data_in213 = map_value_arg213;
   assign  _seachx_data_in214 = map_value_arg214;
   assign  _seachx_data_in215 = map_value_arg215;
   assign  _seachx_data_in216 = map_value_arg216;
   assign  _seachx_data_in217 = map_value_arg217;
   assign  _seachx_data_in218 = map_value_arg218;
   assign  _seachx_data_in219 = map_value_arg219;
   assign  _seachx_data_in220 = map_value_arg220;
   assign  _seachx_data_in221 = map_value_arg221;
   assign  _seachx_data_in222 = map_value_arg222;
   assign  _seachx_data_in225 = map_value_arg225;
   assign  _seachx_data_in226 = map_value_arg226;
   assign  _seachx_data_in227 = map_value_arg227;
   assign  _seachx_data_in228 = map_value_arg228;
   assign  _seachx_data_in229 = map_value_arg229;
   assign  _seachx_data_in230 = map_value_arg230;
   assign  _seachx_data_in231 = map_value_arg231;
   assign  _seachx_data_in232 = map_value_arg232;
   assign  _seachx_data_in233 = map_value_arg233;
   assign  _seachx_data_in234 = map_value_arg234;
   assign  _seachx_data_in235 = map_value_arg235;
   assign  _seachx_data_in236 = map_value_arg236;
   assign  _seachx_data_in237 = map_value_arg237;
   assign  _seachx_data_in238 = map_value_arg238;
   assign  _seachx_data_in239 = map_value_arg239;
   assign  _seachx_data_in240 = map_value_arg240;
   assign  _seachx_data_in241 = map_value_arg241;
   assign  _seachx_data_in242 = map_value_arg242;
   assign  _seachx_data_in243 = map_value_arg243;
   assign  _seachx_data_in244 = map_value_arg244;
   assign  _seachx_data_in245 = map_value_arg245;
   assign  _seachx_data_in246 = map_value_arg246;
   assign  _seachx_data_in247 = map_value_arg247;
   assign  _seachx_data_in248 = map_value_arg248;
   assign  _seachx_data_in249 = map_value_arg249;
   assign  _seachx_data_in250 = map_value_arg250;
   assign  _seachx_data_in251 = map_value_arg251;
   assign  _seachx_data_in252 = map_value_arg252;
   assign  _seachx_data_in253 = map_value_arg253;
   assign  _seachx_data_in254 = map_value_arg254;
   assign  _seachx_data_in257 = map_value_arg257;
   assign  _seachx_data_in258 = map_value_arg258;
   assign  _seachx_data_in259 = map_value_arg259;
   assign  _seachx_data_in260 = map_value_arg260;
   assign  _seachx_data_in261 = map_value_arg261;
   assign  _seachx_data_in262 = map_value_arg262;
   assign  _seachx_data_in263 = map_value_arg263;
   assign  _seachx_data_in264 = map_value_arg264;
   assign  _seachx_data_in265 = map_value_arg265;
   assign  _seachx_data_in266 = map_value_arg266;
   assign  _seachx_data_in267 = map_value_arg267;
   assign  _seachx_data_in268 = map_value_arg268;
   assign  _seachx_data_in269 = map_value_arg269;
   assign  _seachx_data_in270 = map_value_arg270;
   assign  _seachx_data_in271 = map_value_arg271;
   assign  _seachx_data_in272 = map_value_arg272;
   assign  _seachx_data_in273 = map_value_arg273;
   assign  _seachx_data_in274 = map_value_arg274;
   assign  _seachx_data_in275 = map_value_arg275;
   assign  _seachx_data_in276 = map_value_arg276;
   assign  _seachx_data_in277 = map_value_arg277;
   assign  _seachx_data_in278 = map_value_arg278;
   assign  _seachx_data_in279 = map_value_arg279;
   assign  _seachx_data_in280 = map_value_arg280;
   assign  _seachx_data_in281 = map_value_arg281;
   assign  _seachx_data_in282 = map_value_arg282;
   assign  _seachx_data_in283 = map_value_arg283;
   assign  _seachx_data_in284 = map_value_arg284;
   assign  _seachx_data_in285 = map_value_arg285;
   assign  _seachx_data_in286 = map_value_arg286;
   assign  _seachx_data_in289 = map_value_arg289;
   assign  _seachx_data_in290 = map_value_arg290;
   assign  _seachx_data_in291 = map_value_arg291;
   assign  _seachx_data_in292 = map_value_arg292;
   assign  _seachx_data_in293 = map_value_arg293;
   assign  _seachx_data_in294 = map_value_arg294;
   assign  _seachx_data_in295 = map_value_arg295;
   assign  _seachx_data_in296 = map_value_arg296;
   assign  _seachx_data_in297 = map_value_arg297;
   assign  _seachx_data_in298 = map_value_arg298;
   assign  _seachx_data_in299 = map_value_arg299;
   assign  _seachx_data_in300 = map_value_arg300;
   assign  _seachx_data_in301 = map_value_arg301;
   assign  _seachx_data_in302 = map_value_arg302;
   assign  _seachx_data_in303 = map_value_arg303;
   assign  _seachx_data_in304 = map_value_arg304;
   assign  _seachx_data_in305 = map_value_arg305;
   assign  _seachx_data_in306 = map_value_arg306;
   assign  _seachx_data_in307 = map_value_arg307;
   assign  _seachx_data_in308 = map_value_arg308;
   assign  _seachx_data_in309 = map_value_arg309;
   assign  _seachx_data_in310 = map_value_arg310;
   assign  _seachx_data_in311 = map_value_arg311;
   assign  _seachx_data_in312 = map_value_arg312;
   assign  _seachx_data_in313 = map_value_arg313;
   assign  _seachx_data_in314 = map_value_arg314;
   assign  _seachx_data_in315 = map_value_arg315;
   assign  _seachx_data_in316 = map_value_arg316;
   assign  _seachx_data_in317 = map_value_arg317;
   assign  _seachx_data_in318 = map_value_arg318;
   assign  _seachx_data_in321 = map_value_arg321;
   assign  _seachx_data_in322 = map_value_arg322;
   assign  _seachx_data_in323 = map_value_arg323;
   assign  _seachx_data_in324 = map_value_arg324;
   assign  _seachx_data_in325 = map_value_arg325;
   assign  _seachx_data_in326 = map_value_arg326;
   assign  _seachx_data_in327 = map_value_arg327;
   assign  _seachx_data_in328 = map_value_arg328;
   assign  _seachx_data_in329 = map_value_arg329;
   assign  _seachx_data_in330 = map_value_arg330;
   assign  _seachx_data_in331 = map_value_arg331;
   assign  _seachx_data_in332 = map_value_arg332;
   assign  _seachx_data_in333 = map_value_arg333;
   assign  _seachx_data_in334 = map_value_arg334;
   assign  _seachx_data_in335 = map_value_arg335;
   assign  _seachx_data_in336 = map_value_arg336;
   assign  _seachx_data_in337 = map_value_arg337;
   assign  _seachx_data_in338 = map_value_arg338;
   assign  _seachx_data_in339 = map_value_arg339;
   assign  _seachx_data_in340 = map_value_arg340;
   assign  _seachx_data_in341 = map_value_arg341;
   assign  _seachx_data_in342 = map_value_arg342;
   assign  _seachx_data_in343 = map_value_arg343;
   assign  _seachx_data_in344 = map_value_arg344;
   assign  _seachx_data_in345 = map_value_arg345;
   assign  _seachx_data_in346 = map_value_arg346;
   assign  _seachx_data_in347 = map_value_arg347;
   assign  _seachx_data_in348 = map_value_arg348;
   assign  _seachx_data_in349 = map_value_arg349;
   assign  _seachx_data_in350 = map_value_arg350;
   assign  _seachx_data_in353 = map_value_arg353;
   assign  _seachx_data_in354 = map_value_arg354;
   assign  _seachx_data_in355 = map_value_arg355;
   assign  _seachx_data_in356 = map_value_arg356;
   assign  _seachx_data_in357 = map_value_arg357;
   assign  _seachx_data_in358 = map_value_arg358;
   assign  _seachx_data_in359 = map_value_arg359;
   assign  _seachx_data_in360 = map_value_arg360;
   assign  _seachx_data_in361 = map_value_arg361;
   assign  _seachx_data_in362 = map_value_arg362;
   assign  _seachx_data_in363 = map_value_arg363;
   assign  _seachx_data_in364 = map_value_arg364;
   assign  _seachx_data_in365 = map_value_arg365;
   assign  _seachx_data_in366 = map_value_arg366;
   assign  _seachx_data_in367 = map_value_arg367;
   assign  _seachx_data_in368 = map_value_arg368;
   assign  _seachx_data_in369 = map_value_arg369;
   assign  _seachx_data_in370 = map_value_arg370;
   assign  _seachx_data_in371 = map_value_arg371;
   assign  _seachx_data_in372 = map_value_arg372;
   assign  _seachx_data_in373 = map_value_arg373;
   assign  _seachx_data_in374 = map_value_arg374;
   assign  _seachx_data_in375 = map_value_arg375;
   assign  _seachx_data_in376 = map_value_arg376;
   assign  _seachx_data_in377 = map_value_arg377;
   assign  _seachx_data_in378 = map_value_arg378;
   assign  _seachx_data_in379 = map_value_arg379;
   assign  _seachx_data_in380 = map_value_arg380;
   assign  _seachx_data_in381 = map_value_arg381;
   assign  _seachx_data_in382 = map_value_arg382;
   assign  _seachx_data_in385 = map_value_arg385;
   assign  _seachx_data_in386 = map_value_arg386;
   assign  _seachx_data_in387 = map_value_arg387;
   assign  _seachx_data_in388 = map_value_arg388;
   assign  _seachx_data_in389 = map_value_arg389;
   assign  _seachx_data_in390 = map_value_arg390;
   assign  _seachx_data_in391 = map_value_arg391;
   assign  _seachx_data_in392 = map_value_arg392;
   assign  _seachx_data_in393 = map_value_arg393;
   assign  _seachx_data_in394 = map_value_arg394;
   assign  _seachx_data_in395 = map_value_arg395;
   assign  _seachx_data_in396 = map_value_arg396;
   assign  _seachx_data_in397 = map_value_arg397;
   assign  _seachx_data_in398 = map_value_arg398;
   assign  _seachx_data_in399 = map_value_arg399;
   assign  _seachx_data_in400 = map_value_arg400;
   assign  _seachx_data_in401 = map_value_arg401;
   assign  _seachx_data_in402 = map_value_arg402;
   assign  _seachx_data_in403 = map_value_arg403;
   assign  _seachx_data_in404 = map_value_arg404;
   assign  _seachx_data_in405 = map_value_arg405;
   assign  _seachx_data_in406 = map_value_arg406;
   assign  _seachx_data_in407 = map_value_arg407;
   assign  _seachx_data_in408 = map_value_arg408;
   assign  _seachx_data_in409 = map_value_arg409;
   assign  _seachx_data_in410 = map_value_arg410;
   assign  _seachx_data_in411 = map_value_arg411;
   assign  _seachx_data_in412 = map_value_arg412;
   assign  _seachx_data_in413 = map_value_arg413;
   assign  _seachx_data_in414 = map_value_arg414;
   assign  _seachx_data_in417 = map_value_arg417;
   assign  _seachx_data_in418 = map_value_arg418;
   assign  _seachx_data_in419 = map_value_arg419;
   assign  _seachx_data_in420 = map_value_arg420;
   assign  _seachx_data_in421 = map_value_arg421;
   assign  _seachx_data_in422 = map_value_arg422;
   assign  _seachx_data_in423 = map_value_arg423;
   assign  _seachx_data_in424 = map_value_arg424;
   assign  _seachx_data_in425 = map_value_arg425;
   assign  _seachx_data_in426 = map_value_arg426;
   assign  _seachx_data_in427 = map_value_arg427;
   assign  _seachx_data_in428 = map_value_arg428;
   assign  _seachx_data_in429 = map_value_arg429;
   assign  _seachx_data_in430 = map_value_arg430;
   assign  _seachx_data_in431 = map_value_arg431;
   assign  _seachx_data_in432 = map_value_arg432;
   assign  _seachx_data_in433 = map_value_arg433;
   assign  _seachx_data_in434 = map_value_arg434;
   assign  _seachx_data_in435 = map_value_arg435;
   assign  _seachx_data_in436 = map_value_arg436;
   assign  _seachx_data_in437 = map_value_arg437;
   assign  _seachx_data_in438 = map_value_arg438;
   assign  _seachx_data_in439 = map_value_arg439;
   assign  _seachx_data_in440 = map_value_arg440;
   assign  _seachx_data_in441 = map_value_arg441;
   assign  _seachx_data_in442 = map_value_arg442;
   assign  _seachx_data_in443 = map_value_arg443;
   assign  _seachx_data_in444 = map_value_arg444;
   assign  _seachx_data_in445 = map_value_arg445;
   assign  _seachx_data_in446 = map_value_arg446;
   assign  _seachx_data_in449 = map_value_arg449;
   assign  _seachx_data_in450 = map_value_arg450;
   assign  _seachx_data_in451 = map_value_arg451;
   assign  _seachx_data_in452 = map_value_arg452;
   assign  _seachx_data_in453 = map_value_arg453;
   assign  _seachx_data_in454 = map_value_arg454;
   assign  _seachx_data_in455 = map_value_arg455;
   assign  _seachx_data_in456 = map_value_arg456;
   assign  _seachx_data_in457 = map_value_arg457;
   assign  _seachx_data_in458 = map_value_arg458;
   assign  _seachx_data_in459 = map_value_arg459;
   assign  _seachx_data_in460 = map_value_arg460;
   assign  _seachx_data_in461 = map_value_arg461;
   assign  _seachx_data_in462 = map_value_arg462;
   assign  _seachx_data_in463 = map_value_arg463;
   assign  _seachx_data_in464 = map_value_arg464;
   assign  _seachx_data_in465 = map_value_arg465;
   assign  _seachx_data_in466 = map_value_arg466;
   assign  _seachx_data_in467 = map_value_arg467;
   assign  _seachx_data_in468 = map_value_arg468;
   assign  _seachx_data_in469 = map_value_arg469;
   assign  _seachx_data_in470 = map_value_arg470;
   assign  _seachx_data_in471 = map_value_arg471;
   assign  _seachx_data_in472 = map_value_arg472;
   assign  _seachx_data_in473 = map_value_arg473;
   assign  _seachx_data_in474 = map_value_arg474;
   assign  _seachx_data_in475 = map_value_arg475;
   assign  _seachx_data_in476 = map_value_arg476;
   assign  _seachx_data_in477 = map_value_arg477;
   assign  _seachx_data_in478 = map_value_arg478;
   assign  _seachx_in_do = _net_1;
   assign  _seachx_p_reset = p_reset;
   assign  _seachx_m_clock = m_clock;
   assign  _kanwa_x_data_in33 = _seachx_data_out33;
   assign  _kanwa_x_data_in34 = _seachx_data_out34;
   assign  _kanwa_x_data_in35 = _seachx_data_out35;
   assign  _kanwa_x_data_in36 = _seachx_data_out36;
   assign  _kanwa_x_data_in37 = _seachx_data_out37;
   assign  _kanwa_x_data_in38 = _seachx_data_out38;
   assign  _kanwa_x_data_in39 = _seachx_data_out39;
   assign  _kanwa_x_data_in40 = _seachx_data_out40;
   assign  _kanwa_x_data_in41 = _seachx_data_out41;
   assign  _kanwa_x_data_in42 = _seachx_data_out42;
   assign  _kanwa_x_data_in43 = _seachx_data_out43;
   assign  _kanwa_x_data_in44 = _seachx_data_out44;
   assign  _kanwa_x_data_in45 = _seachx_data_out45;
   assign  _kanwa_x_data_in46 = _seachx_data_out46;
   assign  _kanwa_x_data_in47 = _seachx_data_out47;
   assign  _kanwa_x_data_in48 = _seachx_data_out48;
   assign  _kanwa_x_data_in49 = _seachx_data_out49;
   assign  _kanwa_x_data_in50 = _seachx_data_out50;
   assign  _kanwa_x_data_in51 = _seachx_data_out51;
   assign  _kanwa_x_data_in52 = _seachx_data_out52;
   assign  _kanwa_x_data_in53 = _seachx_data_out53;
   assign  _kanwa_x_data_in54 = _seachx_data_out54;
   assign  _kanwa_x_data_in55 = _seachx_data_out55;
   assign  _kanwa_x_data_in56 = _seachx_data_out56;
   assign  _kanwa_x_data_in57 = _seachx_data_out57;
   assign  _kanwa_x_data_in58 = _seachx_data_out58;
   assign  _kanwa_x_data_in59 = _seachx_data_out59;
   assign  _kanwa_x_data_in60 = _seachx_data_out60;
   assign  _kanwa_x_data_in61 = _seachx_data_out61;
   assign  _kanwa_x_data_in62 = _seachx_data_out62;
   assign  _kanwa_x_data_in65 = _seachx_data_out65;
   assign  _kanwa_x_data_in66 = _seachx_data_out66;
   assign  _kanwa_x_data_in67 = _seachx_data_out67;
   assign  _kanwa_x_data_in68 = _seachx_data_out68;
   assign  _kanwa_x_data_in69 = _seachx_data_out69;
   assign  _kanwa_x_data_in70 = _seachx_data_out70;
   assign  _kanwa_x_data_in71 = _seachx_data_out71;
   assign  _kanwa_x_data_in72 = _seachx_data_out72;
   assign  _kanwa_x_data_in73 = _seachx_data_out73;
   assign  _kanwa_x_data_in74 = _seachx_data_out74;
   assign  _kanwa_x_data_in75 = _seachx_data_out75;
   assign  _kanwa_x_data_in76 = _seachx_data_out76;
   assign  _kanwa_x_data_in77 = _seachx_data_out77;
   assign  _kanwa_x_data_in78 = _seachx_data_out78;
   assign  _kanwa_x_data_in79 = _seachx_data_out79;
   assign  _kanwa_x_data_in80 = _seachx_data_out80;
   assign  _kanwa_x_data_in81 = _seachx_data_out81;
   assign  _kanwa_x_data_in82 = _seachx_data_out82;
   assign  _kanwa_x_data_in83 = _seachx_data_out83;
   assign  _kanwa_x_data_in84 = _seachx_data_out84;
   assign  _kanwa_x_data_in85 = _seachx_data_out85;
   assign  _kanwa_x_data_in86 = _seachx_data_out86;
   assign  _kanwa_x_data_in87 = _seachx_data_out87;
   assign  _kanwa_x_data_in88 = _seachx_data_out88;
   assign  _kanwa_x_data_in89 = _seachx_data_out89;
   assign  _kanwa_x_data_in90 = _seachx_data_out90;
   assign  _kanwa_x_data_in91 = _seachx_data_out91;
   assign  _kanwa_x_data_in92 = _seachx_data_out92;
   assign  _kanwa_x_data_in93 = _seachx_data_out93;
   assign  _kanwa_x_data_in94 = _seachx_data_out94;
   assign  _kanwa_x_data_in97 = _seachx_data_out97;
   assign  _kanwa_x_data_in98 = _seachx_data_out98;
   assign  _kanwa_x_data_in99 = _seachx_data_out99;
   assign  _kanwa_x_data_in100 = _seachx_data_out100;
   assign  _kanwa_x_data_in101 = _seachx_data_out101;
   assign  _kanwa_x_data_in102 = _seachx_data_out102;
   assign  _kanwa_x_data_in103 = _seachx_data_out103;
   assign  _kanwa_x_data_in104 = _seachx_data_out104;
   assign  _kanwa_x_data_in105 = _seachx_data_out105;
   assign  _kanwa_x_data_in106 = _seachx_data_out106;
   assign  _kanwa_x_data_in107 = _seachx_data_out107;
   assign  _kanwa_x_data_in108 = _seachx_data_out108;
   assign  _kanwa_x_data_in109 = _seachx_data_out109;
   assign  _kanwa_x_data_in110 = _seachx_data_out110;
   assign  _kanwa_x_data_in111 = _seachx_data_out111;
   assign  _kanwa_x_data_in112 = _seachx_data_out112;
   assign  _kanwa_x_data_in113 = _seachx_data_out113;
   assign  _kanwa_x_data_in114 = _seachx_data_out114;
   assign  _kanwa_x_data_in115 = _seachx_data_out115;
   assign  _kanwa_x_data_in116 = _seachx_data_out116;
   assign  _kanwa_x_data_in117 = _seachx_data_out117;
   assign  _kanwa_x_data_in118 = _seachx_data_out118;
   assign  _kanwa_x_data_in119 = _seachx_data_out119;
   assign  _kanwa_x_data_in120 = _seachx_data_out120;
   assign  _kanwa_x_data_in121 = _seachx_data_out121;
   assign  _kanwa_x_data_in122 = _seachx_data_out122;
   assign  _kanwa_x_data_in123 = _seachx_data_out123;
   assign  _kanwa_x_data_in124 = _seachx_data_out124;
   assign  _kanwa_x_data_in125 = _seachx_data_out125;
   assign  _kanwa_x_data_in126 = _seachx_data_out126;
   assign  _kanwa_x_data_in129 = _seachx_data_out129;
   assign  _kanwa_x_data_in130 = _seachx_data_out130;
   assign  _kanwa_x_data_in131 = _seachx_data_out131;
   assign  _kanwa_x_data_in132 = _seachx_data_out132;
   assign  _kanwa_x_data_in133 = _seachx_data_out133;
   assign  _kanwa_x_data_in134 = _seachx_data_out134;
   assign  _kanwa_x_data_in135 = _seachx_data_out135;
   assign  _kanwa_x_data_in136 = _seachx_data_out136;
   assign  _kanwa_x_data_in137 = _seachx_data_out137;
   assign  _kanwa_x_data_in138 = _seachx_data_out138;
   assign  _kanwa_x_data_in139 = _seachx_data_out139;
   assign  _kanwa_x_data_in140 = _seachx_data_out140;
   assign  _kanwa_x_data_in141 = _seachx_data_out141;
   assign  _kanwa_x_data_in142 = _seachx_data_out142;
   assign  _kanwa_x_data_in143 = _seachx_data_out143;
   assign  _kanwa_x_data_in144 = _seachx_data_out144;
   assign  _kanwa_x_data_in145 = _seachx_data_out145;
   assign  _kanwa_x_data_in146 = _seachx_data_out146;
   assign  _kanwa_x_data_in147 = _seachx_data_out147;
   assign  _kanwa_x_data_in148 = _seachx_data_out148;
   assign  _kanwa_x_data_in149 = _seachx_data_out149;
   assign  _kanwa_x_data_in150 = _seachx_data_out150;
   assign  _kanwa_x_data_in151 = _seachx_data_out151;
   assign  _kanwa_x_data_in152 = _seachx_data_out152;
   assign  _kanwa_x_data_in153 = _seachx_data_out153;
   assign  _kanwa_x_data_in154 = _seachx_data_out154;
   assign  _kanwa_x_data_in155 = _seachx_data_out155;
   assign  _kanwa_x_data_in156 = _seachx_data_out156;
   assign  _kanwa_x_data_in157 = _seachx_data_out157;
   assign  _kanwa_x_data_in158 = _seachx_data_out158;
   assign  _kanwa_x_data_in161 = _seachx_data_out161;
   assign  _kanwa_x_data_in162 = _seachx_data_out162;
   assign  _kanwa_x_data_in163 = _seachx_data_out163;
   assign  _kanwa_x_data_in164 = _seachx_data_out164;
   assign  _kanwa_x_data_in165 = _seachx_data_out165;
   assign  _kanwa_x_data_in166 = _seachx_data_out166;
   assign  _kanwa_x_data_in167 = _seachx_data_out167;
   assign  _kanwa_x_data_in168 = _seachx_data_out168;
   assign  _kanwa_x_data_in169 = _seachx_data_out169;
   assign  _kanwa_x_data_in170 = _seachx_data_out170;
   assign  _kanwa_x_data_in171 = _seachx_data_out171;
   assign  _kanwa_x_data_in172 = _seachx_data_out172;
   assign  _kanwa_x_data_in173 = _seachx_data_out173;
   assign  _kanwa_x_data_in174 = _seachx_data_out174;
   assign  _kanwa_x_data_in175 = _seachx_data_out175;
   assign  _kanwa_x_data_in176 = _seachx_data_out176;
   assign  _kanwa_x_data_in177 = _seachx_data_out177;
   assign  _kanwa_x_data_in178 = _seachx_data_out178;
   assign  _kanwa_x_data_in179 = _seachx_data_out179;
   assign  _kanwa_x_data_in180 = _seachx_data_out180;
   assign  _kanwa_x_data_in181 = _seachx_data_out181;
   assign  _kanwa_x_data_in182 = _seachx_data_out182;
   assign  _kanwa_x_data_in183 = _seachx_data_out183;
   assign  _kanwa_x_data_in184 = _seachx_data_out184;
   assign  _kanwa_x_data_in185 = _seachx_data_out185;
   assign  _kanwa_x_data_in186 = _seachx_data_out186;
   assign  _kanwa_x_data_in187 = _seachx_data_out187;
   assign  _kanwa_x_data_in188 = _seachx_data_out188;
   assign  _kanwa_x_data_in189 = _seachx_data_out189;
   assign  _kanwa_x_data_in190 = _seachx_data_out190;
   assign  _kanwa_x_data_in193 = _seachx_data_out193;
   assign  _kanwa_x_data_in194 = _seachx_data_out194;
   assign  _kanwa_x_data_in195 = _seachx_data_out195;
   assign  _kanwa_x_data_in196 = _seachx_data_out196;
   assign  _kanwa_x_data_in197 = _seachx_data_out197;
   assign  _kanwa_x_data_in198 = _seachx_data_out198;
   assign  _kanwa_x_data_in199 = _seachx_data_out199;
   assign  _kanwa_x_data_in200 = _seachx_data_out200;
   assign  _kanwa_x_data_in201 = _seachx_data_out201;
   assign  _kanwa_x_data_in202 = _seachx_data_out202;
   assign  _kanwa_x_data_in203 = _seachx_data_out203;
   assign  _kanwa_x_data_in204 = _seachx_data_out204;
   assign  _kanwa_x_data_in205 = _seachx_data_out205;
   assign  _kanwa_x_data_in206 = _seachx_data_out206;
   assign  _kanwa_x_data_in207 = _seachx_data_out207;
   assign  _kanwa_x_data_in208 = _seachx_data_out208;
   assign  _kanwa_x_data_in209 = _seachx_data_out209;
   assign  _kanwa_x_data_in210 = _seachx_data_out210;
   assign  _kanwa_x_data_in211 = _seachx_data_out211;
   assign  _kanwa_x_data_in212 = _seachx_data_out212;
   assign  _kanwa_x_data_in213 = _seachx_data_out213;
   assign  _kanwa_x_data_in214 = _seachx_data_out214;
   assign  _kanwa_x_data_in215 = _seachx_data_out215;
   assign  _kanwa_x_data_in216 = _seachx_data_out216;
   assign  _kanwa_x_data_in217 = _seachx_data_out217;
   assign  _kanwa_x_data_in218 = _seachx_data_out218;
   assign  _kanwa_x_data_in219 = _seachx_data_out219;
   assign  _kanwa_x_data_in220 = _seachx_data_out220;
   assign  _kanwa_x_data_in221 = _seachx_data_out221;
   assign  _kanwa_x_data_in222 = _seachx_data_out222;
   assign  _kanwa_x_data_in225 = _seachx_data_out225;
   assign  _kanwa_x_data_in226 = _seachx_data_out226;
   assign  _kanwa_x_data_in227 = _seachx_data_out227;
   assign  _kanwa_x_data_in228 = _seachx_data_out228;
   assign  _kanwa_x_data_in229 = _seachx_data_out229;
   assign  _kanwa_x_data_in230 = _seachx_data_out230;
   assign  _kanwa_x_data_in231 = _seachx_data_out231;
   assign  _kanwa_x_data_in232 = _seachx_data_out232;
   assign  _kanwa_x_data_in233 = _seachx_data_out233;
   assign  _kanwa_x_data_in234 = _seachx_data_out234;
   assign  _kanwa_x_data_in235 = _seachx_data_out235;
   assign  _kanwa_x_data_in236 = _seachx_data_out236;
   assign  _kanwa_x_data_in237 = _seachx_data_out237;
   assign  _kanwa_x_data_in238 = _seachx_data_out238;
   assign  _kanwa_x_data_in239 = _seachx_data_out239;
   assign  _kanwa_x_data_in240 = _seachx_data_out240;
   assign  _kanwa_x_data_in241 = _seachx_data_out241;
   assign  _kanwa_x_data_in242 = _seachx_data_out242;
   assign  _kanwa_x_data_in243 = _seachx_data_out243;
   assign  _kanwa_x_data_in244 = _seachx_data_out244;
   assign  _kanwa_x_data_in245 = _seachx_data_out245;
   assign  _kanwa_x_data_in246 = _seachx_data_out246;
   assign  _kanwa_x_data_in247 = _seachx_data_out247;
   assign  _kanwa_x_data_in248 = _seachx_data_out248;
   assign  _kanwa_x_data_in249 = _seachx_data_out249;
   assign  _kanwa_x_data_in250 = _seachx_data_out250;
   assign  _kanwa_x_data_in251 = _seachx_data_out251;
   assign  _kanwa_x_data_in252 = _seachx_data_out252;
   assign  _kanwa_x_data_in253 = _seachx_data_out253;
   assign  _kanwa_x_data_in254 = _seachx_data_out254;
   assign  _kanwa_x_data_in257 = _seachx_data_out257;
   assign  _kanwa_x_data_in258 = _seachx_data_out258;
   assign  _kanwa_x_data_in259 = _seachx_data_out259;
   assign  _kanwa_x_data_in260 = _seachx_data_out260;
   assign  _kanwa_x_data_in261 = _seachx_data_out261;
   assign  _kanwa_x_data_in262 = _seachx_data_out262;
   assign  _kanwa_x_data_in263 = _seachx_data_out263;
   assign  _kanwa_x_data_in264 = _seachx_data_out264;
   assign  _kanwa_x_data_in265 = _seachx_data_out265;
   assign  _kanwa_x_data_in266 = _seachx_data_out266;
   assign  _kanwa_x_data_in267 = _seachx_data_out267;
   assign  _kanwa_x_data_in268 = _seachx_data_out268;
   assign  _kanwa_x_data_in269 = _seachx_data_out269;
   assign  _kanwa_x_data_in270 = _seachx_data_out270;
   assign  _kanwa_x_data_in271 = _seachx_data_out271;
   assign  _kanwa_x_data_in272 = _seachx_data_out272;
   assign  _kanwa_x_data_in273 = _seachx_data_out273;
   assign  _kanwa_x_data_in274 = _seachx_data_out274;
   assign  _kanwa_x_data_in275 = _seachx_data_out275;
   assign  _kanwa_x_data_in276 = _seachx_data_out276;
   assign  _kanwa_x_data_in277 = _seachx_data_out277;
   assign  _kanwa_x_data_in278 = _seachx_data_out278;
   assign  _kanwa_x_data_in279 = _seachx_data_out279;
   assign  _kanwa_x_data_in280 = _seachx_data_out280;
   assign  _kanwa_x_data_in281 = _seachx_data_out281;
   assign  _kanwa_x_data_in282 = _seachx_data_out282;
   assign  _kanwa_x_data_in283 = _seachx_data_out283;
   assign  _kanwa_x_data_in284 = _seachx_data_out284;
   assign  _kanwa_x_data_in285 = _seachx_data_out285;
   assign  _kanwa_x_data_in286 = _seachx_data_out286;
   assign  _kanwa_x_data_in289 = _seachx_data_out289;
   assign  _kanwa_x_data_in290 = _seachx_data_out290;
   assign  _kanwa_x_data_in291 = _seachx_data_out291;
   assign  _kanwa_x_data_in292 = _seachx_data_out292;
   assign  _kanwa_x_data_in293 = _seachx_data_out293;
   assign  _kanwa_x_data_in294 = _seachx_data_out294;
   assign  _kanwa_x_data_in295 = _seachx_data_out295;
   assign  _kanwa_x_data_in296 = _seachx_data_out296;
   assign  _kanwa_x_data_in297 = _seachx_data_out297;
   assign  _kanwa_x_data_in298 = _seachx_data_out298;
   assign  _kanwa_x_data_in299 = _seachx_data_out299;
   assign  _kanwa_x_data_in300 = _seachx_data_out300;
   assign  _kanwa_x_data_in301 = _seachx_data_out301;
   assign  _kanwa_x_data_in302 = _seachx_data_out302;
   assign  _kanwa_x_data_in303 = _seachx_data_out303;
   assign  _kanwa_x_data_in304 = _seachx_data_out304;
   assign  _kanwa_x_data_in305 = _seachx_data_out305;
   assign  _kanwa_x_data_in306 = _seachx_data_out306;
   assign  _kanwa_x_data_in307 = _seachx_data_out307;
   assign  _kanwa_x_data_in308 = _seachx_data_out308;
   assign  _kanwa_x_data_in309 = _seachx_data_out309;
   assign  _kanwa_x_data_in310 = _seachx_data_out310;
   assign  _kanwa_x_data_in311 = _seachx_data_out311;
   assign  _kanwa_x_data_in312 = _seachx_data_out312;
   assign  _kanwa_x_data_in313 = _seachx_data_out313;
   assign  _kanwa_x_data_in314 = _seachx_data_out314;
   assign  _kanwa_x_data_in315 = _seachx_data_out315;
   assign  _kanwa_x_data_in316 = _seachx_data_out316;
   assign  _kanwa_x_data_in317 = _seachx_data_out317;
   assign  _kanwa_x_data_in318 = _seachx_data_out318;
   assign  _kanwa_x_data_in321 = _seachx_data_out321;
   assign  _kanwa_x_data_in322 = _seachx_data_out322;
   assign  _kanwa_x_data_in323 = _seachx_data_out323;
   assign  _kanwa_x_data_in324 = _seachx_data_out324;
   assign  _kanwa_x_data_in325 = _seachx_data_out325;
   assign  _kanwa_x_data_in326 = _seachx_data_out326;
   assign  _kanwa_x_data_in327 = _seachx_data_out327;
   assign  _kanwa_x_data_in328 = _seachx_data_out328;
   assign  _kanwa_x_data_in329 = _seachx_data_out329;
   assign  _kanwa_x_data_in330 = _seachx_data_out330;
   assign  _kanwa_x_data_in331 = _seachx_data_out331;
   assign  _kanwa_x_data_in332 = _seachx_data_out332;
   assign  _kanwa_x_data_in333 = _seachx_data_out333;
   assign  _kanwa_x_data_in334 = _seachx_data_out334;
   assign  _kanwa_x_data_in335 = _seachx_data_out335;
   assign  _kanwa_x_data_in336 = _seachx_data_out336;
   assign  _kanwa_x_data_in337 = _seachx_data_out337;
   assign  _kanwa_x_data_in338 = _seachx_data_out338;
   assign  _kanwa_x_data_in339 = _seachx_data_out339;
   assign  _kanwa_x_data_in340 = _seachx_data_out340;
   assign  _kanwa_x_data_in341 = _seachx_data_out341;
   assign  _kanwa_x_data_in342 = _seachx_data_out342;
   assign  _kanwa_x_data_in343 = _seachx_data_out343;
   assign  _kanwa_x_data_in344 = _seachx_data_out344;
   assign  _kanwa_x_data_in345 = _seachx_data_out345;
   assign  _kanwa_x_data_in346 = _seachx_data_out346;
   assign  _kanwa_x_data_in347 = _seachx_data_out347;
   assign  _kanwa_x_data_in348 = _seachx_data_out348;
   assign  _kanwa_x_data_in349 = _seachx_data_out349;
   assign  _kanwa_x_data_in350 = _seachx_data_out350;
   assign  _kanwa_x_data_in353 = _seachx_data_out353;
   assign  _kanwa_x_data_in354 = _seachx_data_out354;
   assign  _kanwa_x_data_in355 = _seachx_data_out355;
   assign  _kanwa_x_data_in356 = _seachx_data_out356;
   assign  _kanwa_x_data_in357 = _seachx_data_out357;
   assign  _kanwa_x_data_in358 = _seachx_data_out358;
   assign  _kanwa_x_data_in359 = _seachx_data_out359;
   assign  _kanwa_x_data_in360 = _seachx_data_out360;
   assign  _kanwa_x_data_in361 = _seachx_data_out361;
   assign  _kanwa_x_data_in362 = _seachx_data_out362;
   assign  _kanwa_x_data_in363 = _seachx_data_out363;
   assign  _kanwa_x_data_in364 = _seachx_data_out364;
   assign  _kanwa_x_data_in365 = _seachx_data_out365;
   assign  _kanwa_x_data_in366 = _seachx_data_out366;
   assign  _kanwa_x_data_in367 = _seachx_data_out367;
   assign  _kanwa_x_data_in368 = _seachx_data_out368;
   assign  _kanwa_x_data_in369 = _seachx_data_out369;
   assign  _kanwa_x_data_in370 = _seachx_data_out370;
   assign  _kanwa_x_data_in371 = _seachx_data_out371;
   assign  _kanwa_x_data_in372 = _seachx_data_out372;
   assign  _kanwa_x_data_in373 = _seachx_data_out373;
   assign  _kanwa_x_data_in374 = _seachx_data_out374;
   assign  _kanwa_x_data_in375 = _seachx_data_out375;
   assign  _kanwa_x_data_in376 = _seachx_data_out376;
   assign  _kanwa_x_data_in377 = _seachx_data_out377;
   assign  _kanwa_x_data_in378 = _seachx_data_out378;
   assign  _kanwa_x_data_in379 = _seachx_data_out379;
   assign  _kanwa_x_data_in380 = _seachx_data_out380;
   assign  _kanwa_x_data_in381 = _seachx_data_out381;
   assign  _kanwa_x_data_in382 = _seachx_data_out382;
   assign  _kanwa_x_data_in385 = _seachx_data_out385;
   assign  _kanwa_x_data_in386 = _seachx_data_out386;
   assign  _kanwa_x_data_in387 = _seachx_data_out387;
   assign  _kanwa_x_data_in388 = _seachx_data_out388;
   assign  _kanwa_x_data_in389 = _seachx_data_out389;
   assign  _kanwa_x_data_in390 = _seachx_data_out390;
   assign  _kanwa_x_data_in391 = _seachx_data_out391;
   assign  _kanwa_x_data_in392 = _seachx_data_out392;
   assign  _kanwa_x_data_in393 = _seachx_data_out393;
   assign  _kanwa_x_data_in394 = _seachx_data_out394;
   assign  _kanwa_x_data_in395 = _seachx_data_out395;
   assign  _kanwa_x_data_in396 = _seachx_data_out396;
   assign  _kanwa_x_data_in397 = _seachx_data_out397;
   assign  _kanwa_x_data_in398 = _seachx_data_out398;
   assign  _kanwa_x_data_in399 = _seachx_data_out399;
   assign  _kanwa_x_data_in400 = _seachx_data_out400;
   assign  _kanwa_x_data_in401 = _seachx_data_out401;
   assign  _kanwa_x_data_in402 = _seachx_data_out402;
   assign  _kanwa_x_data_in403 = _seachx_data_out403;
   assign  _kanwa_x_data_in404 = _seachx_data_out404;
   assign  _kanwa_x_data_in405 = _seachx_data_out405;
   assign  _kanwa_x_data_in406 = _seachx_data_out406;
   assign  _kanwa_x_data_in407 = _seachx_data_out407;
   assign  _kanwa_x_data_in408 = _seachx_data_out408;
   assign  _kanwa_x_data_in409 = _seachx_data_out409;
   assign  _kanwa_x_data_in410 = _seachx_data_out410;
   assign  _kanwa_x_data_in411 = _seachx_data_out411;
   assign  _kanwa_x_data_in412 = _seachx_data_out412;
   assign  _kanwa_x_data_in413 = _seachx_data_out413;
   assign  _kanwa_x_data_in414 = _seachx_data_out414;
   assign  _kanwa_x_data_in417 = _seachx_data_out417;
   assign  _kanwa_x_data_in418 = _seachx_data_out418;
   assign  _kanwa_x_data_in419 = _seachx_data_out419;
   assign  _kanwa_x_data_in420 = _seachx_data_out420;
   assign  _kanwa_x_data_in421 = _seachx_data_out421;
   assign  _kanwa_x_data_in422 = _seachx_data_out422;
   assign  _kanwa_x_data_in423 = _seachx_data_out423;
   assign  _kanwa_x_data_in424 = _seachx_data_out424;
   assign  _kanwa_x_data_in425 = _seachx_data_out425;
   assign  _kanwa_x_data_in426 = _seachx_data_out426;
   assign  _kanwa_x_data_in427 = _seachx_data_out427;
   assign  _kanwa_x_data_in428 = _seachx_data_out428;
   assign  _kanwa_x_data_in429 = _seachx_data_out429;
   assign  _kanwa_x_data_in430 = _seachx_data_out430;
   assign  _kanwa_x_data_in431 = _seachx_data_out431;
   assign  _kanwa_x_data_in432 = _seachx_data_out432;
   assign  _kanwa_x_data_in433 = _seachx_data_out433;
   assign  _kanwa_x_data_in434 = _seachx_data_out434;
   assign  _kanwa_x_data_in435 = _seachx_data_out435;
   assign  _kanwa_x_data_in436 = _seachx_data_out436;
   assign  _kanwa_x_data_in437 = _seachx_data_out437;
   assign  _kanwa_x_data_in438 = _seachx_data_out438;
   assign  _kanwa_x_data_in439 = _seachx_data_out439;
   assign  _kanwa_x_data_in440 = _seachx_data_out440;
   assign  _kanwa_x_data_in441 = _seachx_data_out441;
   assign  _kanwa_x_data_in442 = _seachx_data_out442;
   assign  _kanwa_x_data_in443 = _seachx_data_out443;
   assign  _kanwa_x_data_in444 = _seachx_data_out444;
   assign  _kanwa_x_data_in445 = _seachx_data_out445;
   assign  _kanwa_x_data_in446 = _seachx_data_out446;
   assign  _kanwa_x_data_in449 = _seachx_data_out449;
   assign  _kanwa_x_data_in450 = _seachx_data_out450;
   assign  _kanwa_x_data_in451 = _seachx_data_out451;
   assign  _kanwa_x_data_in452 = _seachx_data_out452;
   assign  _kanwa_x_data_in453 = _seachx_data_out453;
   assign  _kanwa_x_data_in454 = _seachx_data_out454;
   assign  _kanwa_x_data_in455 = _seachx_data_out455;
   assign  _kanwa_x_data_in456 = _seachx_data_out456;
   assign  _kanwa_x_data_in457 = _seachx_data_out457;
   assign  _kanwa_x_data_in458 = _seachx_data_out458;
   assign  _kanwa_x_data_in459 = _seachx_data_out459;
   assign  _kanwa_x_data_in460 = _seachx_data_out460;
   assign  _kanwa_x_data_in461 = _seachx_data_out461;
   assign  _kanwa_x_data_in462 = _seachx_data_out462;
   assign  _kanwa_x_data_in463 = _seachx_data_out463;
   assign  _kanwa_x_data_in464 = _seachx_data_out464;
   assign  _kanwa_x_data_in465 = _seachx_data_out465;
   assign  _kanwa_x_data_in466 = _seachx_data_out466;
   assign  _kanwa_x_data_in467 = _seachx_data_out467;
   assign  _kanwa_x_data_in468 = _seachx_data_out468;
   assign  _kanwa_x_data_in469 = _seachx_data_out469;
   assign  _kanwa_x_data_in470 = _seachx_data_out470;
   assign  _kanwa_x_data_in471 = _seachx_data_out471;
   assign  _kanwa_x_data_in472 = _seachx_data_out472;
   assign  _kanwa_x_data_in473 = _seachx_data_out473;
   assign  _kanwa_x_data_in474 = _seachx_data_out474;
   assign  _kanwa_x_data_in475 = _seachx_data_out475;
   assign  _kanwa_x_data_in476 = _seachx_data_out476;
   assign  _kanwa_x_data_in477 = _seachx_data_out477;
   assign  _kanwa_x_data_in478 = _seachx_data_out478;
   assign  _kanwa_x_start = _seachx_startplot;
   assign  _kanwa_x_goal = _seachx_goalplot;
   assign  _kanwa_x_in_do = _seachx_out_do;
   assign  _kanwa_x_p_reset = p_reset;
   assign  _kanwa_x_m_clock = m_clock;
   assign  _kouka_x_data_in33 = _kanwa_x_data_out33;
   assign  _kouka_x_data_in34 = _kanwa_x_data_out34;
   assign  _kouka_x_data_in35 = _kanwa_x_data_out35;
   assign  _kouka_x_data_in36 = _kanwa_x_data_out36;
   assign  _kouka_x_data_in37 = _kanwa_x_data_out37;
   assign  _kouka_x_data_in38 = _kanwa_x_data_out38;
   assign  _kouka_x_data_in39 = _kanwa_x_data_out39;
   assign  _kouka_x_data_in40 = _kanwa_x_data_out40;
   assign  _kouka_x_data_in41 = _kanwa_x_data_out41;
   assign  _kouka_x_data_in42 = _kanwa_x_data_out42;
   assign  _kouka_x_data_in43 = _kanwa_x_data_out43;
   assign  _kouka_x_data_in44 = _kanwa_x_data_out44;
   assign  _kouka_x_data_in45 = _kanwa_x_data_out45;
   assign  _kouka_x_data_in46 = _kanwa_x_data_out46;
   assign  _kouka_x_data_in47 = _kanwa_x_data_out47;
   assign  _kouka_x_data_in48 = _kanwa_x_data_out48;
   assign  _kouka_x_data_in49 = _kanwa_x_data_out49;
   assign  _kouka_x_data_in50 = _kanwa_x_data_out50;
   assign  _kouka_x_data_in51 = _kanwa_x_data_out51;
   assign  _kouka_x_data_in52 = _kanwa_x_data_out52;
   assign  _kouka_x_data_in53 = _kanwa_x_data_out53;
   assign  _kouka_x_data_in54 = _kanwa_x_data_out54;
   assign  _kouka_x_data_in55 = _kanwa_x_data_out55;
   assign  _kouka_x_data_in56 = _kanwa_x_data_out56;
   assign  _kouka_x_data_in57 = _kanwa_x_data_out57;
   assign  _kouka_x_data_in58 = _kanwa_x_data_out58;
   assign  _kouka_x_data_in59 = _kanwa_x_data_out59;
   assign  _kouka_x_data_in60 = _kanwa_x_data_out60;
   assign  _kouka_x_data_in61 = _kanwa_x_data_out61;
   assign  _kouka_x_data_in62 = _kanwa_x_data_out62;
   assign  _kouka_x_data_in65 = _kanwa_x_data_out65;
   assign  _kouka_x_data_in66 = _kanwa_x_data_out66;
   assign  _kouka_x_data_in67 = _kanwa_x_data_out67;
   assign  _kouka_x_data_in68 = _kanwa_x_data_out68;
   assign  _kouka_x_data_in69 = _kanwa_x_data_out69;
   assign  _kouka_x_data_in70 = _kanwa_x_data_out70;
   assign  _kouka_x_data_in71 = _kanwa_x_data_out71;
   assign  _kouka_x_data_in72 = _kanwa_x_data_out72;
   assign  _kouka_x_data_in73 = _kanwa_x_data_out73;
   assign  _kouka_x_data_in74 = _kanwa_x_data_out74;
   assign  _kouka_x_data_in75 = _kanwa_x_data_out75;
   assign  _kouka_x_data_in76 = _kanwa_x_data_out76;
   assign  _kouka_x_data_in77 = _kanwa_x_data_out77;
   assign  _kouka_x_data_in78 = _kanwa_x_data_out78;
   assign  _kouka_x_data_in79 = _kanwa_x_data_out79;
   assign  _kouka_x_data_in80 = _kanwa_x_data_out80;
   assign  _kouka_x_data_in81 = _kanwa_x_data_out81;
   assign  _kouka_x_data_in82 = _kanwa_x_data_out82;
   assign  _kouka_x_data_in83 = _kanwa_x_data_out83;
   assign  _kouka_x_data_in84 = _kanwa_x_data_out84;
   assign  _kouka_x_data_in85 = _kanwa_x_data_out85;
   assign  _kouka_x_data_in86 = _kanwa_x_data_out86;
   assign  _kouka_x_data_in87 = _kanwa_x_data_out87;
   assign  _kouka_x_data_in88 = _kanwa_x_data_out88;
   assign  _kouka_x_data_in89 = _kanwa_x_data_out89;
   assign  _kouka_x_data_in90 = _kanwa_x_data_out90;
   assign  _kouka_x_data_in91 = _kanwa_x_data_out91;
   assign  _kouka_x_data_in92 = _kanwa_x_data_out92;
   assign  _kouka_x_data_in93 = _kanwa_x_data_out93;
   assign  _kouka_x_data_in94 = _kanwa_x_data_out94;
   assign  _kouka_x_data_in97 = _kanwa_x_data_out97;
   assign  _kouka_x_data_in98 = _kanwa_x_data_out98;
   assign  _kouka_x_data_in99 = _kanwa_x_data_out99;
   assign  _kouka_x_data_in100 = _kanwa_x_data_out100;
   assign  _kouka_x_data_in101 = _kanwa_x_data_out101;
   assign  _kouka_x_data_in102 = _kanwa_x_data_out102;
   assign  _kouka_x_data_in103 = _kanwa_x_data_out103;
   assign  _kouka_x_data_in104 = _kanwa_x_data_out104;
   assign  _kouka_x_data_in105 = _kanwa_x_data_out105;
   assign  _kouka_x_data_in106 = _kanwa_x_data_out106;
   assign  _kouka_x_data_in107 = _kanwa_x_data_out107;
   assign  _kouka_x_data_in108 = _kanwa_x_data_out108;
   assign  _kouka_x_data_in109 = _kanwa_x_data_out109;
   assign  _kouka_x_data_in110 = _kanwa_x_data_out110;
   assign  _kouka_x_data_in111 = _kanwa_x_data_out111;
   assign  _kouka_x_data_in112 = _kanwa_x_data_out112;
   assign  _kouka_x_data_in113 = _kanwa_x_data_out113;
   assign  _kouka_x_data_in114 = _kanwa_x_data_out114;
   assign  _kouka_x_data_in115 = _kanwa_x_data_out115;
   assign  _kouka_x_data_in116 = _kanwa_x_data_out116;
   assign  _kouka_x_data_in117 = _kanwa_x_data_out117;
   assign  _kouka_x_data_in118 = _kanwa_x_data_out118;
   assign  _kouka_x_data_in119 = _kanwa_x_data_out119;
   assign  _kouka_x_data_in120 = _kanwa_x_data_out120;
   assign  _kouka_x_data_in121 = _kanwa_x_data_out121;
   assign  _kouka_x_data_in122 = _kanwa_x_data_out122;
   assign  _kouka_x_data_in123 = _kanwa_x_data_out123;
   assign  _kouka_x_data_in124 = _kanwa_x_data_out124;
   assign  _kouka_x_data_in125 = _kanwa_x_data_out125;
   assign  _kouka_x_data_in126 = _kanwa_x_data_out126;
   assign  _kouka_x_data_in129 = _kanwa_x_data_out129;
   assign  _kouka_x_data_in130 = _kanwa_x_data_out130;
   assign  _kouka_x_data_in131 = _kanwa_x_data_out131;
   assign  _kouka_x_data_in132 = _kanwa_x_data_out132;
   assign  _kouka_x_data_in133 = _kanwa_x_data_out133;
   assign  _kouka_x_data_in134 = _kanwa_x_data_out134;
   assign  _kouka_x_data_in135 = _kanwa_x_data_out135;
   assign  _kouka_x_data_in136 = _kanwa_x_data_out136;
   assign  _kouka_x_data_in137 = _kanwa_x_data_out137;
   assign  _kouka_x_data_in138 = _kanwa_x_data_out138;
   assign  _kouka_x_data_in139 = _kanwa_x_data_out139;
   assign  _kouka_x_data_in140 = _kanwa_x_data_out140;
   assign  _kouka_x_data_in141 = _kanwa_x_data_out141;
   assign  _kouka_x_data_in142 = _kanwa_x_data_out142;
   assign  _kouka_x_data_in143 = _kanwa_x_data_out143;
   assign  _kouka_x_data_in144 = _kanwa_x_data_out144;
   assign  _kouka_x_data_in145 = _kanwa_x_data_out145;
   assign  _kouka_x_data_in146 = _kanwa_x_data_out146;
   assign  _kouka_x_data_in147 = _kanwa_x_data_out147;
   assign  _kouka_x_data_in148 = _kanwa_x_data_out148;
   assign  _kouka_x_data_in149 = _kanwa_x_data_out149;
   assign  _kouka_x_data_in150 = _kanwa_x_data_out150;
   assign  _kouka_x_data_in151 = _kanwa_x_data_out151;
   assign  _kouka_x_data_in152 = _kanwa_x_data_out152;
   assign  _kouka_x_data_in153 = _kanwa_x_data_out153;
   assign  _kouka_x_data_in154 = _kanwa_x_data_out154;
   assign  _kouka_x_data_in155 = _kanwa_x_data_out155;
   assign  _kouka_x_data_in156 = _kanwa_x_data_out156;
   assign  _kouka_x_data_in157 = _kanwa_x_data_out157;
   assign  _kouka_x_data_in158 = _kanwa_x_data_out158;
   assign  _kouka_x_data_in161 = _kanwa_x_data_out161;
   assign  _kouka_x_data_in162 = _kanwa_x_data_out162;
   assign  _kouka_x_data_in163 = _kanwa_x_data_out163;
   assign  _kouka_x_data_in164 = _kanwa_x_data_out164;
   assign  _kouka_x_data_in165 = _kanwa_x_data_out165;
   assign  _kouka_x_data_in166 = _kanwa_x_data_out166;
   assign  _kouka_x_data_in167 = _kanwa_x_data_out167;
   assign  _kouka_x_data_in168 = _kanwa_x_data_out168;
   assign  _kouka_x_data_in169 = _kanwa_x_data_out169;
   assign  _kouka_x_data_in170 = _kanwa_x_data_out170;
   assign  _kouka_x_data_in171 = _kanwa_x_data_out171;
   assign  _kouka_x_data_in172 = _kanwa_x_data_out172;
   assign  _kouka_x_data_in173 = _kanwa_x_data_out173;
   assign  _kouka_x_data_in174 = _kanwa_x_data_out174;
   assign  _kouka_x_data_in175 = _kanwa_x_data_out175;
   assign  _kouka_x_data_in176 = _kanwa_x_data_out176;
   assign  _kouka_x_data_in177 = _kanwa_x_data_out177;
   assign  _kouka_x_data_in178 = _kanwa_x_data_out178;
   assign  _kouka_x_data_in179 = _kanwa_x_data_out179;
   assign  _kouka_x_data_in180 = _kanwa_x_data_out180;
   assign  _kouka_x_data_in181 = _kanwa_x_data_out181;
   assign  _kouka_x_data_in182 = _kanwa_x_data_out182;
   assign  _kouka_x_data_in183 = _kanwa_x_data_out183;
   assign  _kouka_x_data_in184 = _kanwa_x_data_out184;
   assign  _kouka_x_data_in185 = _kanwa_x_data_out185;
   assign  _kouka_x_data_in186 = _kanwa_x_data_out186;
   assign  _kouka_x_data_in187 = _kanwa_x_data_out187;
   assign  _kouka_x_data_in188 = _kanwa_x_data_out188;
   assign  _kouka_x_data_in189 = _kanwa_x_data_out189;
   assign  _kouka_x_data_in190 = _kanwa_x_data_out190;
   assign  _kouka_x_data_in193 = _kanwa_x_data_out193;
   assign  _kouka_x_data_in194 = _kanwa_x_data_out194;
   assign  _kouka_x_data_in195 = _kanwa_x_data_out195;
   assign  _kouka_x_data_in196 = _kanwa_x_data_out196;
   assign  _kouka_x_data_in197 = _kanwa_x_data_out197;
   assign  _kouka_x_data_in198 = _kanwa_x_data_out198;
   assign  _kouka_x_data_in199 = _kanwa_x_data_out199;
   assign  _kouka_x_data_in200 = _kanwa_x_data_out200;
   assign  _kouka_x_data_in201 = _kanwa_x_data_out201;
   assign  _kouka_x_data_in202 = _kanwa_x_data_out202;
   assign  _kouka_x_data_in203 = _kanwa_x_data_out203;
   assign  _kouka_x_data_in204 = _kanwa_x_data_out204;
   assign  _kouka_x_data_in205 = _kanwa_x_data_out205;
   assign  _kouka_x_data_in206 = _kanwa_x_data_out206;
   assign  _kouka_x_data_in207 = _kanwa_x_data_out207;
   assign  _kouka_x_data_in208 = _kanwa_x_data_out208;
   assign  _kouka_x_data_in209 = _kanwa_x_data_out209;
   assign  _kouka_x_data_in210 = _kanwa_x_data_out210;
   assign  _kouka_x_data_in211 = _kanwa_x_data_out211;
   assign  _kouka_x_data_in212 = _kanwa_x_data_out212;
   assign  _kouka_x_data_in213 = _kanwa_x_data_out213;
   assign  _kouka_x_data_in214 = _kanwa_x_data_out214;
   assign  _kouka_x_data_in215 = _kanwa_x_data_out215;
   assign  _kouka_x_data_in216 = _kanwa_x_data_out216;
   assign  _kouka_x_data_in217 = _kanwa_x_data_out217;
   assign  _kouka_x_data_in218 = _kanwa_x_data_out218;
   assign  _kouka_x_data_in219 = _kanwa_x_data_out219;
   assign  _kouka_x_data_in220 = _kanwa_x_data_out220;
   assign  _kouka_x_data_in221 = _kanwa_x_data_out221;
   assign  _kouka_x_data_in222 = _kanwa_x_data_out222;
   assign  _kouka_x_data_in225 = _kanwa_x_data_out225;
   assign  _kouka_x_data_in226 = _kanwa_x_data_out226;
   assign  _kouka_x_data_in227 = _kanwa_x_data_out227;
   assign  _kouka_x_data_in228 = _kanwa_x_data_out228;
   assign  _kouka_x_data_in229 = _kanwa_x_data_out229;
   assign  _kouka_x_data_in230 = _kanwa_x_data_out230;
   assign  _kouka_x_data_in231 = _kanwa_x_data_out231;
   assign  _kouka_x_data_in232 = _kanwa_x_data_out232;
   assign  _kouka_x_data_in233 = _kanwa_x_data_out233;
   assign  _kouka_x_data_in234 = _kanwa_x_data_out234;
   assign  _kouka_x_data_in235 = _kanwa_x_data_out235;
   assign  _kouka_x_data_in236 = _kanwa_x_data_out236;
   assign  _kouka_x_data_in237 = _kanwa_x_data_out237;
   assign  _kouka_x_data_in238 = _kanwa_x_data_out238;
   assign  _kouka_x_data_in239 = _kanwa_x_data_out239;
   assign  _kouka_x_data_in240 = _kanwa_x_data_out240;
   assign  _kouka_x_data_in241 = _kanwa_x_data_out241;
   assign  _kouka_x_data_in242 = _kanwa_x_data_out242;
   assign  _kouka_x_data_in243 = _kanwa_x_data_out243;
   assign  _kouka_x_data_in244 = _kanwa_x_data_out244;
   assign  _kouka_x_data_in245 = _kanwa_x_data_out245;
   assign  _kouka_x_data_in246 = _kanwa_x_data_out246;
   assign  _kouka_x_data_in247 = _kanwa_x_data_out247;
   assign  _kouka_x_data_in248 = _kanwa_x_data_out248;
   assign  _kouka_x_data_in249 = _kanwa_x_data_out249;
   assign  _kouka_x_data_in250 = _kanwa_x_data_out250;
   assign  _kouka_x_data_in251 = _kanwa_x_data_out251;
   assign  _kouka_x_data_in252 = _kanwa_x_data_out252;
   assign  _kouka_x_data_in253 = _kanwa_x_data_out253;
   assign  _kouka_x_data_in254 = _kanwa_x_data_out254;
   assign  _kouka_x_data_in257 = _kanwa_x_data_out257;
   assign  _kouka_x_data_in258 = _kanwa_x_data_out258;
   assign  _kouka_x_data_in259 = _kanwa_x_data_out259;
   assign  _kouka_x_data_in260 = _kanwa_x_data_out260;
   assign  _kouka_x_data_in261 = _kanwa_x_data_out261;
   assign  _kouka_x_data_in262 = _kanwa_x_data_out262;
   assign  _kouka_x_data_in263 = _kanwa_x_data_out263;
   assign  _kouka_x_data_in264 = _kanwa_x_data_out264;
   assign  _kouka_x_data_in265 = _kanwa_x_data_out265;
   assign  _kouka_x_data_in266 = _kanwa_x_data_out266;
   assign  _kouka_x_data_in267 = _kanwa_x_data_out267;
   assign  _kouka_x_data_in268 = _kanwa_x_data_out268;
   assign  _kouka_x_data_in269 = _kanwa_x_data_out269;
   assign  _kouka_x_data_in270 = _kanwa_x_data_out270;
   assign  _kouka_x_data_in271 = _kanwa_x_data_out271;
   assign  _kouka_x_data_in272 = _kanwa_x_data_out272;
   assign  _kouka_x_data_in273 = _kanwa_x_data_out273;
   assign  _kouka_x_data_in274 = _kanwa_x_data_out274;
   assign  _kouka_x_data_in275 = _kanwa_x_data_out275;
   assign  _kouka_x_data_in276 = _kanwa_x_data_out276;
   assign  _kouka_x_data_in277 = _kanwa_x_data_out277;
   assign  _kouka_x_data_in278 = _kanwa_x_data_out278;
   assign  _kouka_x_data_in279 = _kanwa_x_data_out279;
   assign  _kouka_x_data_in280 = _kanwa_x_data_out280;
   assign  _kouka_x_data_in281 = _kanwa_x_data_out281;
   assign  _kouka_x_data_in282 = _kanwa_x_data_out282;
   assign  _kouka_x_data_in283 = _kanwa_x_data_out283;
   assign  _kouka_x_data_in284 = _kanwa_x_data_out284;
   assign  _kouka_x_data_in285 = _kanwa_x_data_out285;
   assign  _kouka_x_data_in286 = _kanwa_x_data_out286;
   assign  _kouka_x_data_in289 = _kanwa_x_data_out289;
   assign  _kouka_x_data_in290 = _kanwa_x_data_out290;
   assign  _kouka_x_data_in291 = _kanwa_x_data_out291;
   assign  _kouka_x_data_in292 = _kanwa_x_data_out292;
   assign  _kouka_x_data_in293 = _kanwa_x_data_out293;
   assign  _kouka_x_data_in294 = _kanwa_x_data_out294;
   assign  _kouka_x_data_in295 = _kanwa_x_data_out295;
   assign  _kouka_x_data_in296 = _kanwa_x_data_out296;
   assign  _kouka_x_data_in297 = _kanwa_x_data_out297;
   assign  _kouka_x_data_in298 = _kanwa_x_data_out298;
   assign  _kouka_x_data_in299 = _kanwa_x_data_out299;
   assign  _kouka_x_data_in300 = _kanwa_x_data_out300;
   assign  _kouka_x_data_in301 = _kanwa_x_data_out301;
   assign  _kouka_x_data_in302 = _kanwa_x_data_out302;
   assign  _kouka_x_data_in303 = _kanwa_x_data_out303;
   assign  _kouka_x_data_in304 = _kanwa_x_data_out304;
   assign  _kouka_x_data_in305 = _kanwa_x_data_out305;
   assign  _kouka_x_data_in306 = _kanwa_x_data_out306;
   assign  _kouka_x_data_in307 = _kanwa_x_data_out307;
   assign  _kouka_x_data_in308 = _kanwa_x_data_out308;
   assign  _kouka_x_data_in309 = _kanwa_x_data_out309;
   assign  _kouka_x_data_in310 = _kanwa_x_data_out310;
   assign  _kouka_x_data_in311 = _kanwa_x_data_out311;
   assign  _kouka_x_data_in312 = _kanwa_x_data_out312;
   assign  _kouka_x_data_in313 = _kanwa_x_data_out313;
   assign  _kouka_x_data_in314 = _kanwa_x_data_out314;
   assign  _kouka_x_data_in315 = _kanwa_x_data_out315;
   assign  _kouka_x_data_in316 = _kanwa_x_data_out316;
   assign  _kouka_x_data_in317 = _kanwa_x_data_out317;
   assign  _kouka_x_data_in318 = _kanwa_x_data_out318;
   assign  _kouka_x_data_in321 = _kanwa_x_data_out321;
   assign  _kouka_x_data_in322 = _kanwa_x_data_out322;
   assign  _kouka_x_data_in323 = _kanwa_x_data_out323;
   assign  _kouka_x_data_in324 = _kanwa_x_data_out324;
   assign  _kouka_x_data_in325 = _kanwa_x_data_out325;
   assign  _kouka_x_data_in326 = _kanwa_x_data_out326;
   assign  _kouka_x_data_in327 = _kanwa_x_data_out327;
   assign  _kouka_x_data_in328 = _kanwa_x_data_out328;
   assign  _kouka_x_data_in329 = _kanwa_x_data_out329;
   assign  _kouka_x_data_in330 = _kanwa_x_data_out330;
   assign  _kouka_x_data_in331 = _kanwa_x_data_out331;
   assign  _kouka_x_data_in332 = _kanwa_x_data_out332;
   assign  _kouka_x_data_in333 = _kanwa_x_data_out333;
   assign  _kouka_x_data_in334 = _kanwa_x_data_out334;
   assign  _kouka_x_data_in335 = _kanwa_x_data_out335;
   assign  _kouka_x_data_in336 = _kanwa_x_data_out336;
   assign  _kouka_x_data_in337 = _kanwa_x_data_out337;
   assign  _kouka_x_data_in338 = _kanwa_x_data_out338;
   assign  _kouka_x_data_in339 = _kanwa_x_data_out339;
   assign  _kouka_x_data_in340 = _kanwa_x_data_out340;
   assign  _kouka_x_data_in341 = _kanwa_x_data_out341;
   assign  _kouka_x_data_in342 = _kanwa_x_data_out342;
   assign  _kouka_x_data_in343 = _kanwa_x_data_out343;
   assign  _kouka_x_data_in344 = _kanwa_x_data_out344;
   assign  _kouka_x_data_in345 = _kanwa_x_data_out345;
   assign  _kouka_x_data_in346 = _kanwa_x_data_out346;
   assign  _kouka_x_data_in347 = _kanwa_x_data_out347;
   assign  _kouka_x_data_in348 = _kanwa_x_data_out348;
   assign  _kouka_x_data_in349 = _kanwa_x_data_out349;
   assign  _kouka_x_data_in350 = _kanwa_x_data_out350;
   assign  _kouka_x_data_in353 = _kanwa_x_data_out353;
   assign  _kouka_x_data_in354 = _kanwa_x_data_out354;
   assign  _kouka_x_data_in355 = _kanwa_x_data_out355;
   assign  _kouka_x_data_in356 = _kanwa_x_data_out356;
   assign  _kouka_x_data_in357 = _kanwa_x_data_out357;
   assign  _kouka_x_data_in358 = _kanwa_x_data_out358;
   assign  _kouka_x_data_in359 = _kanwa_x_data_out359;
   assign  _kouka_x_data_in360 = _kanwa_x_data_out360;
   assign  _kouka_x_data_in361 = _kanwa_x_data_out361;
   assign  _kouka_x_data_in362 = _kanwa_x_data_out362;
   assign  _kouka_x_data_in363 = _kanwa_x_data_out363;
   assign  _kouka_x_data_in364 = _kanwa_x_data_out364;
   assign  _kouka_x_data_in365 = _kanwa_x_data_out365;
   assign  _kouka_x_data_in366 = _kanwa_x_data_out366;
   assign  _kouka_x_data_in367 = _kanwa_x_data_out367;
   assign  _kouka_x_data_in368 = _kanwa_x_data_out368;
   assign  _kouka_x_data_in369 = _kanwa_x_data_out369;
   assign  _kouka_x_data_in370 = _kanwa_x_data_out370;
   assign  _kouka_x_data_in371 = _kanwa_x_data_out371;
   assign  _kouka_x_data_in372 = _kanwa_x_data_out372;
   assign  _kouka_x_data_in373 = _kanwa_x_data_out373;
   assign  _kouka_x_data_in374 = _kanwa_x_data_out374;
   assign  _kouka_x_data_in375 = _kanwa_x_data_out375;
   assign  _kouka_x_data_in376 = _kanwa_x_data_out376;
   assign  _kouka_x_data_in377 = _kanwa_x_data_out377;
   assign  _kouka_x_data_in378 = _kanwa_x_data_out378;
   assign  _kouka_x_data_in379 = _kanwa_x_data_out379;
   assign  _kouka_x_data_in380 = _kanwa_x_data_out380;
   assign  _kouka_x_data_in381 = _kanwa_x_data_out381;
   assign  _kouka_x_data_in382 = _kanwa_x_data_out382;
   assign  _kouka_x_data_in385 = _kanwa_x_data_out385;
   assign  _kouka_x_data_in386 = _kanwa_x_data_out386;
   assign  _kouka_x_data_in387 = _kanwa_x_data_out387;
   assign  _kouka_x_data_in388 = _kanwa_x_data_out388;
   assign  _kouka_x_data_in389 = _kanwa_x_data_out389;
   assign  _kouka_x_data_in390 = _kanwa_x_data_out390;
   assign  _kouka_x_data_in391 = _kanwa_x_data_out391;
   assign  _kouka_x_data_in392 = _kanwa_x_data_out392;
   assign  _kouka_x_data_in393 = _kanwa_x_data_out393;
   assign  _kouka_x_data_in394 = _kanwa_x_data_out394;
   assign  _kouka_x_data_in395 = _kanwa_x_data_out395;
   assign  _kouka_x_data_in396 = _kanwa_x_data_out396;
   assign  _kouka_x_data_in397 = _kanwa_x_data_out397;
   assign  _kouka_x_data_in398 = _kanwa_x_data_out398;
   assign  _kouka_x_data_in399 = _kanwa_x_data_out399;
   assign  _kouka_x_data_in400 = _kanwa_x_data_out400;
   assign  _kouka_x_data_in401 = _kanwa_x_data_out401;
   assign  _kouka_x_data_in402 = _kanwa_x_data_out402;
   assign  _kouka_x_data_in403 = _kanwa_x_data_out403;
   assign  _kouka_x_data_in404 = _kanwa_x_data_out404;
   assign  _kouka_x_data_in405 = _kanwa_x_data_out405;
   assign  _kouka_x_data_in406 = _kanwa_x_data_out406;
   assign  _kouka_x_data_in407 = _kanwa_x_data_out407;
   assign  _kouka_x_data_in408 = _kanwa_x_data_out408;
   assign  _kouka_x_data_in409 = _kanwa_x_data_out409;
   assign  _kouka_x_data_in410 = _kanwa_x_data_out410;
   assign  _kouka_x_data_in411 = _kanwa_x_data_out411;
   assign  _kouka_x_data_in412 = _kanwa_x_data_out412;
   assign  _kouka_x_data_in413 = _kanwa_x_data_out413;
   assign  _kouka_x_data_in414 = _kanwa_x_data_out414;
   assign  _kouka_x_data_in417 = _kanwa_x_data_out417;
   assign  _kouka_x_data_in418 = _kanwa_x_data_out418;
   assign  _kouka_x_data_in419 = _kanwa_x_data_out419;
   assign  _kouka_x_data_in420 = _kanwa_x_data_out420;
   assign  _kouka_x_data_in421 = _kanwa_x_data_out421;
   assign  _kouka_x_data_in422 = _kanwa_x_data_out422;
   assign  _kouka_x_data_in423 = _kanwa_x_data_out423;
   assign  _kouka_x_data_in424 = _kanwa_x_data_out424;
   assign  _kouka_x_data_in425 = _kanwa_x_data_out425;
   assign  _kouka_x_data_in426 = _kanwa_x_data_out426;
   assign  _kouka_x_data_in427 = _kanwa_x_data_out427;
   assign  _kouka_x_data_in428 = _kanwa_x_data_out428;
   assign  _kouka_x_data_in429 = _kanwa_x_data_out429;
   assign  _kouka_x_data_in430 = _kanwa_x_data_out430;
   assign  _kouka_x_data_in431 = _kanwa_x_data_out431;
   assign  _kouka_x_data_in432 = _kanwa_x_data_out432;
   assign  _kouka_x_data_in433 = _kanwa_x_data_out433;
   assign  _kouka_x_data_in434 = _kanwa_x_data_out434;
   assign  _kouka_x_data_in435 = _kanwa_x_data_out435;
   assign  _kouka_x_data_in436 = _kanwa_x_data_out436;
   assign  _kouka_x_data_in437 = _kanwa_x_data_out437;
   assign  _kouka_x_data_in438 = _kanwa_x_data_out438;
   assign  _kouka_x_data_in439 = _kanwa_x_data_out439;
   assign  _kouka_x_data_in440 = _kanwa_x_data_out440;
   assign  _kouka_x_data_in441 = _kanwa_x_data_out441;
   assign  _kouka_x_data_in442 = _kanwa_x_data_out442;
   assign  _kouka_x_data_in443 = _kanwa_x_data_out443;
   assign  _kouka_x_data_in444 = _kanwa_x_data_out444;
   assign  _kouka_x_data_in445 = _kanwa_x_data_out445;
   assign  _kouka_x_data_in446 = _kanwa_x_data_out446;
   assign  _kouka_x_data_in449 = _kanwa_x_data_out449;
   assign  _kouka_x_data_in450 = _kanwa_x_data_out450;
   assign  _kouka_x_data_in451 = _kanwa_x_data_out451;
   assign  _kouka_x_data_in452 = _kanwa_x_data_out452;
   assign  _kouka_x_data_in453 = _kanwa_x_data_out453;
   assign  _kouka_x_data_in454 = _kanwa_x_data_out454;
   assign  _kouka_x_data_in455 = _kanwa_x_data_out455;
   assign  _kouka_x_data_in456 = _kanwa_x_data_out456;
   assign  _kouka_x_data_in457 = _kanwa_x_data_out457;
   assign  _kouka_x_data_in458 = _kanwa_x_data_out458;
   assign  _kouka_x_data_in459 = _kanwa_x_data_out459;
   assign  _kouka_x_data_in460 = _kanwa_x_data_out460;
   assign  _kouka_x_data_in461 = _kanwa_x_data_out461;
   assign  _kouka_x_data_in462 = _kanwa_x_data_out462;
   assign  _kouka_x_data_in463 = _kanwa_x_data_out463;
   assign  _kouka_x_data_in464 = _kanwa_x_data_out464;
   assign  _kouka_x_data_in465 = _kanwa_x_data_out465;
   assign  _kouka_x_data_in466 = _kanwa_x_data_out466;
   assign  _kouka_x_data_in467 = _kanwa_x_data_out467;
   assign  _kouka_x_data_in468 = _kanwa_x_data_out468;
   assign  _kouka_x_data_in469 = _kanwa_x_data_out469;
   assign  _kouka_x_data_in470 = _kanwa_x_data_out470;
   assign  _kouka_x_data_in471 = _kanwa_x_data_out471;
   assign  _kouka_x_data_in472 = _kanwa_x_data_out472;
   assign  _kouka_x_data_in473 = _kanwa_x_data_out473;
   assign  _kouka_x_data_in474 = _kanwa_x_data_out474;
   assign  _kouka_x_data_in475 = _kanwa_x_data_out475;
   assign  _kouka_x_data_in476 = _kanwa_x_data_out476;
   assign  _kouka_x_data_in477 = _kanwa_x_data_out477;
   assign  _kouka_x_data_in478 = _kanwa_x_data_out478;
   assign  _kouka_x_start = _seachx_startplot;
   assign  _kouka_x_goal = _seachx_goalplot;
   assign  _kouka_x_in_do = _kanwa_x_out_do;
   assign  _kouka_x_p_reset = p_reset;
   assign  _kouka_x_m_clock = m_clock;
   assign  _net_1 = (in_do|_reg_0);
   assign  _net_2 = (in_do|_reg_0);
   assign  _net_3 = (in_do|_reg_0);
   assign  _net_4 = (in_do|_reg_0);
   assign  _net_5 = (in_do|_reg_0);
   assign  _net_6 = (in_do|_reg_0);
   assign  _net_7 = (in_do|_reg_0);
   assign  _net_8 = (in_do|_reg_0);
   assign  _net_9 = (in_do|_reg_0);
   assign  _net_10 = (in_do|_reg_0);
   assign  _net_11 = (in_do|_reg_0);
   assign  _net_12 = (in_do|_reg_0);
   assign  _net_13 = (in_do|_reg_0);
   assign  _net_14 = (in_do|_reg_0);
   assign  _net_15 = (in_do|_reg_0);
   assign  _net_16 = (in_do|_reg_0);
   assign  _net_17 = (in_do|_reg_0);
   assign  _net_18 = (in_do|_reg_0);
   assign  _net_19 = (in_do|_reg_0);
   assign  _net_20 = (in_do|_reg_0);
   assign  _net_21 = (in_do|_reg_0);
   assign  _net_22 = (in_do|_reg_0);
   assign  _net_23 = (in_do|_reg_0);
   assign  _net_24 = (in_do|_reg_0);
   assign  _net_25 = (in_do|_reg_0);
   assign  _net_26 = (in_do|_reg_0);
   assign  _net_27 = (in_do|_reg_0);
   assign  _net_28 = (in_do|_reg_0);
   assign  _net_29 = (in_do|_reg_0);
   assign  _net_30 = (in_do|_reg_0);
   assign  _net_31 = (in_do|_reg_0);
   assign  _net_32 = (in_do|_reg_0);
   assign  _net_33 = (in_do|_reg_0);
   assign  _net_34 = (in_do|_reg_0);
   assign  _net_35 = (in_do|_reg_0);
   assign  _net_36 = (in_do|_reg_0);
   assign  _net_37 = (in_do|_reg_0);
   assign  _net_38 = (in_do|_reg_0);
   assign  _net_39 = (in_do|_reg_0);
   assign  _net_40 = (in_do|_reg_0);
   assign  _net_41 = (in_do|_reg_0);
   assign  _net_42 = (in_do|_reg_0);
   assign  _net_43 = (in_do|_reg_0);
   assign  _net_44 = (in_do|_reg_0);
   assign  _net_45 = (in_do|_reg_0);
   assign  _net_46 = (in_do|_reg_0);
   assign  _net_47 = (in_do|_reg_0);
   assign  _net_48 = (in_do|_reg_0);
   assign  _net_49 = (in_do|_reg_0);
   assign  _net_50 = (in_do|_reg_0);
   assign  _net_51 = (in_do|_reg_0);
   assign  _net_52 = (in_do|_reg_0);
   assign  _net_53 = (in_do|_reg_0);
   assign  _net_54 = (in_do|_reg_0);
   assign  _net_55 = (in_do|_reg_0);
   assign  _net_56 = (in_do|_reg_0);
   assign  _net_57 = (in_do|_reg_0);
   assign  _net_58 = (in_do|_reg_0);
   assign  _net_59 = (in_do|_reg_0);
   assign  _net_60 = (in_do|_reg_0);
   assign  _net_61 = (in_do|_reg_0);
   assign  _net_62 = (in_do|_reg_0);
   assign  _net_63 = (in_do|_reg_0);
   assign  _net_64 = (in_do|_reg_0);
   assign  _net_65 = (in_do|_reg_0);
   assign  _net_66 = (in_do|_reg_0);
   assign  _net_67 = (in_do|_reg_0);
   assign  _net_68 = (in_do|_reg_0);
   assign  _net_69 = (in_do|_reg_0);
   assign  _net_70 = (in_do|_reg_0);
   assign  _net_71 = (in_do|_reg_0);
   assign  _net_72 = (in_do|_reg_0);
   assign  _net_73 = (in_do|_reg_0);
   assign  _net_74 = (in_do|_reg_0);
   assign  _net_75 = (in_do|_reg_0);
   assign  _net_76 = (in_do|_reg_0);
   assign  _net_77 = (in_do|_reg_0);
   assign  _net_78 = (in_do|_reg_0);
   assign  _net_79 = (in_do|_reg_0);
   assign  _net_80 = (in_do|_reg_0);
   assign  _net_81 = (in_do|_reg_0);
   assign  _net_82 = (in_do|_reg_0);
   assign  _net_83 = (in_do|_reg_0);
   assign  _net_84 = (in_do|_reg_0);
   assign  _net_85 = (in_do|_reg_0);
   assign  _net_86 = (in_do|_reg_0);
   assign  _net_87 = (in_do|_reg_0);
   assign  _net_88 = (in_do|_reg_0);
   assign  _net_89 = (in_do|_reg_0);
   assign  _net_90 = (in_do|_reg_0);
   assign  _net_91 = (in_do|_reg_0);
   assign  _net_92 = (in_do|_reg_0);
   assign  _net_93 = (in_do|_reg_0);
   assign  _net_94 = (in_do|_reg_0);
   assign  _net_95 = (in_do|_reg_0);
   assign  _net_96 = (in_do|_reg_0);
   assign  _net_97 = (in_do|_reg_0);
   assign  _net_98 = (in_do|_reg_0);
   assign  _net_99 = (in_do|_reg_0);
   assign  _net_100 = (in_do|_reg_0);
   assign  _net_101 = (in_do|_reg_0);
   assign  _net_102 = (in_do|_reg_0);
   assign  _net_103 = (in_do|_reg_0);
   assign  _net_104 = (in_do|_reg_0);
   assign  _net_105 = (in_do|_reg_0);
   assign  _net_106 = (in_do|_reg_0);
   assign  _net_107 = (in_do|_reg_0);
   assign  _net_108 = (in_do|_reg_0);
   assign  _net_109 = (in_do|_reg_0);
   assign  _net_110 = (in_do|_reg_0);
   assign  _net_111 = (in_do|_reg_0);
   assign  _net_112 = (in_do|_reg_0);
   assign  _net_113 = (in_do|_reg_0);
   assign  _net_114 = (in_do|_reg_0);
   assign  _net_115 = (in_do|_reg_0);
   assign  _net_116 = (in_do|_reg_0);
   assign  _net_117 = (in_do|_reg_0);
   assign  _net_118 = (in_do|_reg_0);
   assign  _net_119 = (in_do|_reg_0);
   assign  _net_120 = (in_do|_reg_0);
   assign  _net_121 = (in_do|_reg_0);
   assign  _net_122 = (in_do|_reg_0);
   assign  _net_123 = (in_do|_reg_0);
   assign  _net_124 = (in_do|_reg_0);
   assign  _net_125 = (in_do|_reg_0);
   assign  _net_126 = (in_do|_reg_0);
   assign  _net_127 = (in_do|_reg_0);
   assign  _net_128 = (in_do|_reg_0);
   assign  _net_129 = (in_do|_reg_0);
   assign  _net_130 = (in_do|_reg_0);
   assign  _net_131 = (in_do|_reg_0);
   assign  _net_132 = (in_do|_reg_0);
   assign  _net_133 = (in_do|_reg_0);
   assign  _net_134 = (in_do|_reg_0);
   assign  _net_135 = (in_do|_reg_0);
   assign  _net_136 = (in_do|_reg_0);
   assign  _net_137 = (in_do|_reg_0);
   assign  _net_138 = (in_do|_reg_0);
   assign  _net_139 = (in_do|_reg_0);
   assign  _net_140 = (in_do|_reg_0);
   assign  _net_141 = (in_do|_reg_0);
   assign  _net_142 = (in_do|_reg_0);
   assign  _net_143 = (in_do|_reg_0);
   assign  _net_144 = (in_do|_reg_0);
   assign  _net_145 = (in_do|_reg_0);
   assign  _net_146 = (in_do|_reg_0);
   assign  _net_147 = (in_do|_reg_0);
   assign  _net_148 = (in_do|_reg_0);
   assign  _net_149 = (in_do|_reg_0);
   assign  _net_150 = (in_do|_reg_0);
   assign  _net_151 = (in_do|_reg_0);
   assign  _net_152 = (in_do|_reg_0);
   assign  _net_153 = (in_do|_reg_0);
   assign  _net_154 = (in_do|_reg_0);
   assign  _net_155 = (in_do|_reg_0);
   assign  _net_156 = (in_do|_reg_0);
   assign  _net_157 = (in_do|_reg_0);
   assign  _net_158 = (in_do|_reg_0);
   assign  _net_159 = (in_do|_reg_0);
   assign  _net_160 = (in_do|_reg_0);
   assign  _net_161 = (in_do|_reg_0);
   assign  _net_162 = (in_do|_reg_0);
   assign  _net_163 = (in_do|_reg_0);
   assign  _net_164 = (in_do|_reg_0);
   assign  _net_165 = (in_do|_reg_0);
   assign  _net_166 = (in_do|_reg_0);
   assign  _net_167 = (in_do|_reg_0);
   assign  _net_168 = (in_do|_reg_0);
   assign  _net_169 = (in_do|_reg_0);
   assign  _net_170 = (in_do|_reg_0);
   assign  _net_171 = (in_do|_reg_0);
   assign  _net_172 = (in_do|_reg_0);
   assign  _net_173 = (in_do|_reg_0);
   assign  _net_174 = (in_do|_reg_0);
   assign  _net_175 = (in_do|_reg_0);
   assign  _net_176 = (in_do|_reg_0);
   assign  _net_177 = (in_do|_reg_0);
   assign  _net_178 = (in_do|_reg_0);
   assign  _net_179 = (in_do|_reg_0);
   assign  _net_180 = (in_do|_reg_0);
   assign  _net_181 = (in_do|_reg_0);
   assign  _net_182 = (in_do|_reg_0);
   assign  _net_183 = (in_do|_reg_0);
   assign  _net_184 = (in_do|_reg_0);
   assign  _net_185 = (in_do|_reg_0);
   assign  _net_186 = (in_do|_reg_0);
   assign  _net_187 = (in_do|_reg_0);
   assign  _net_188 = (in_do|_reg_0);
   assign  _net_189 = (in_do|_reg_0);
   assign  _net_190 = (in_do|_reg_0);
   assign  _net_191 = (in_do|_reg_0);
   assign  _net_192 = (in_do|_reg_0);
   assign  _net_193 = (in_do|_reg_0);
   assign  _net_194 = (in_do|_reg_0);
   assign  _net_195 = (in_do|_reg_0);
   assign  _net_196 = (in_do|_reg_0);
   assign  _net_197 = (in_do|_reg_0);
   assign  _net_198 = (in_do|_reg_0);
   assign  _net_199 = (in_do|_reg_0);
   assign  _net_200 = (in_do|_reg_0);
   assign  _net_201 = (in_do|_reg_0);
   assign  _net_202 = (in_do|_reg_0);
   assign  _net_203 = (in_do|_reg_0);
   assign  _net_204 = (in_do|_reg_0);
   assign  _net_205 = (in_do|_reg_0);
   assign  _net_206 = (in_do|_reg_0);
   assign  _net_207 = (in_do|_reg_0);
   assign  _net_208 = (in_do|_reg_0);
   assign  _net_209 = (in_do|_reg_0);
   assign  _net_210 = (in_do|_reg_0);
   assign  _net_211 = (in_do|_reg_0);
   assign  _net_212 = (in_do|_reg_0);
   assign  _net_213 = (in_do|_reg_0);
   assign  _net_214 = (in_do|_reg_0);
   assign  _net_215 = (in_do|_reg_0);
   assign  _net_216 = (in_do|_reg_0);
   assign  _net_217 = (in_do|_reg_0);
   assign  _net_218 = (in_do|_reg_0);
   assign  _net_219 = (in_do|_reg_0);
   assign  _net_220 = (in_do|_reg_0);
   assign  _net_221 = (in_do|_reg_0);
   assign  _net_222 = (in_do|_reg_0);
   assign  _net_223 = (in_do|_reg_0);
   assign  _net_224 = (in_do|_reg_0);
   assign  _net_225 = (in_do|_reg_0);
   assign  _net_226 = (in_do|_reg_0);
   assign  _net_227 = (in_do|_reg_0);
   assign  _net_228 = (in_do|_reg_0);
   assign  _net_229 = (in_do|_reg_0);
   assign  _net_230 = (in_do|_reg_0);
   assign  _net_231 = (in_do|_reg_0);
   assign  _net_232 = (in_do|_reg_0);
   assign  _net_233 = (in_do|_reg_0);
   assign  _net_234 = (in_do|_reg_0);
   assign  _net_235 = (in_do|_reg_0);
   assign  _net_236 = (in_do|_reg_0);
   assign  _net_237 = (in_do|_reg_0);
   assign  _net_238 = (in_do|_reg_0);
   assign  _net_239 = (in_do|_reg_0);
   assign  _net_240 = (in_do|_reg_0);
   assign  _net_241 = (in_do|_reg_0);
   assign  _net_242 = (in_do|_reg_0);
   assign  _net_243 = (in_do|_reg_0);
   assign  _net_244 = (in_do|_reg_0);
   assign  _net_245 = (in_do|_reg_0);
   assign  _net_246 = (in_do|_reg_0);
   assign  _net_247 = (in_do|_reg_0);
   assign  _net_248 = (in_do|_reg_0);
   assign  _net_249 = (in_do|_reg_0);
   assign  _net_250 = (in_do|_reg_0);
   assign  _net_251 = (in_do|_reg_0);
   assign  _net_252 = (in_do|_reg_0);
   assign  _net_253 = (in_do|_reg_0);
   assign  _net_254 = (in_do|_reg_0);
   assign  _net_255 = (in_do|_reg_0);
   assign  _net_256 = (in_do|_reg_0);
   assign  _net_257 = (in_do|_reg_0);
   assign  _net_258 = (in_do|_reg_0);
   assign  _net_259 = (in_do|_reg_0);
   assign  _net_260 = (in_do|_reg_0);
   assign  _net_261 = (in_do|_reg_0);
   assign  _net_262 = (in_do|_reg_0);
   assign  _net_263 = (in_do|_reg_0);
   assign  _net_264 = (in_do|_reg_0);
   assign  _net_265 = (in_do|_reg_0);
   assign  _net_266 = (in_do|_reg_0);
   assign  _net_267 = (in_do|_reg_0);
   assign  _net_268 = (in_do|_reg_0);
   assign  _net_269 = (in_do|_reg_0);
   assign  _net_270 = (in_do|_reg_0);
   assign  _net_271 = (in_do|_reg_0);
   assign  _net_272 = (in_do|_reg_0);
   assign  _net_273 = (in_do|_reg_0);
   assign  _net_274 = (in_do|_reg_0);
   assign  _net_275 = (in_do|_reg_0);
   assign  _net_276 = (in_do|_reg_0);
   assign  _net_277 = (in_do|_reg_0);
   assign  _net_278 = (in_do|_reg_0);
   assign  _net_279 = (in_do|_reg_0);
   assign  _net_280 = (in_do|_reg_0);
   assign  _net_281 = (in_do|_reg_0);
   assign  _net_282 = (in_do|_reg_0);
   assign  _net_283 = (in_do|_reg_0);
   assign  _net_284 = (in_do|_reg_0);
   assign  _net_285 = (in_do|_reg_0);
   assign  _net_286 = (in_do|_reg_0);
   assign  _net_287 = (in_do|_reg_0);
   assign  _net_288 = (in_do|_reg_0);
   assign  _net_289 = (in_do|_reg_0);
   assign  _net_290 = (in_do|_reg_0);
   assign  _net_291 = (in_do|_reg_0);
   assign  _net_292 = (in_do|_reg_0);
   assign  _net_293 = (in_do|_reg_0);
   assign  _net_294 = (in_do|_reg_0);
   assign  _net_295 = (in_do|_reg_0);
   assign  _net_296 = (in_do|_reg_0);
   assign  _net_297 = (in_do|_reg_0);
   assign  _net_298 = (in_do|_reg_0);
   assign  _net_299 = (in_do|_reg_0);
   assign  _net_300 = (in_do|_reg_0);
   assign  _net_301 = (in_do|_reg_0);
   assign  _net_302 = (in_do|_reg_0);
   assign  _net_303 = (in_do|_reg_0);
   assign  _net_304 = (in_do|_reg_0);
   assign  _net_305 = (in_do|_reg_0);
   assign  _net_306 = (in_do|_reg_0);
   assign  _net_307 = (in_do|_reg_0);
   assign  _net_308 = (in_do|_reg_0);
   assign  _net_309 = (in_do|_reg_0);
   assign  _net_310 = (in_do|_reg_0);
   assign  _net_311 = (in_do|_reg_0);
   assign  _net_312 = (in_do|_reg_0);
   assign  _net_313 = (in_do|_reg_0);
   assign  _net_314 = (in_do|_reg_0);
   assign  _net_315 = (in_do|_reg_0);
   assign  _net_316 = (in_do|_reg_0);
   assign  _net_317 = (in_do|_reg_0);
   assign  _net_318 = (in_do|_reg_0);
   assign  _net_319 = (in_do|_reg_0);
   assign  _net_320 = (in_do|_reg_0);
   assign  _net_321 = (in_do|_reg_0);
   assign  _net_322 = (in_do|_reg_0);
   assign  _net_323 = (in_do|_reg_0);
   assign  _net_324 = (in_do|_reg_0);
   assign  _net_325 = (in_do|_reg_0);
   assign  _net_326 = (in_do|_reg_0);
   assign  _net_327 = (in_do|_reg_0);
   assign  _net_328 = (in_do|_reg_0);
   assign  _net_329 = (in_do|_reg_0);
   assign  _net_330 = (in_do|_reg_0);
   assign  _net_331 = (in_do|_reg_0);
   assign  _net_332 = (in_do|_reg_0);
   assign  _net_333 = (in_do|_reg_0);
   assign  _net_334 = (in_do|_reg_0);
   assign  _net_335 = (in_do|_reg_0);
   assign  _net_336 = (in_do|_reg_0);
   assign  _net_337 = (in_do|_reg_0);
   assign  _net_338 = (in_do|_reg_0);
   assign  _net_339 = (in_do|_reg_0);
   assign  _net_340 = (in_do|_reg_0);
   assign  _net_341 = (in_do|_reg_0);
   assign  _net_342 = (in_do|_reg_0);
   assign  _net_343 = (in_do|_reg_0);
   assign  _net_344 = (in_do|_reg_0);
   assign  _net_345 = (in_do|_reg_0);
   assign  _net_346 = (in_do|_reg_0);
   assign  _net_347 = (in_do|_reg_0);
   assign  _net_348 = (in_do|_reg_0);
   assign  _net_349 = (in_do|_reg_0);
   assign  _net_350 = (in_do|_reg_0);
   assign  _net_351 = (in_do|_reg_0);
   assign  _net_352 = (in_do|_reg_0);
   assign  _net_353 = (in_do|_reg_0);
   assign  _net_354 = (in_do|_reg_0);
   assign  _net_355 = (in_do|_reg_0);
   assign  _net_356 = (in_do|_reg_0);
   assign  _net_357 = (in_do|_reg_0);
   assign  _net_358 = (in_do|_reg_0);
   assign  _net_359 = (in_do|_reg_0);
   assign  _net_360 = (in_do|_reg_0);
   assign  _net_361 = (in_do|_reg_0);
   assign  _net_362 = (in_do|_reg_0);
   assign  _net_363 = (in_do|_reg_0);
   assign  _net_364 = (in_do|_reg_0);
   assign  _net_365 = (in_do|_reg_0);
   assign  _net_366 = (in_do|_reg_0);
   assign  _net_367 = (in_do|_reg_0);
   assign  _net_368 = (in_do|_reg_0);
   assign  _net_369 = (in_do|_reg_0);
   assign  _net_370 = (in_do|_reg_0);
   assign  _net_371 = (in_do|_reg_0);
   assign  _net_372 = (in_do|_reg_0);
   assign  _net_373 = (in_do|_reg_0);
   assign  _net_374 = (in_do|_reg_0);
   assign  _net_375 = (in_do|_reg_0);
   assign  _net_376 = (in_do|_reg_0);
   assign  _net_377 = (in_do|_reg_0);
   assign  _net_378 = (in_do|_reg_0);
   assign  _net_379 = (in_do|_reg_0);
   assign  _net_380 = (in_do|_reg_0);
   assign  _net_381 = (in_do|_reg_0);
   assign  _net_382 = (in_do|_reg_0);
   assign  _net_383 = (in_do|_reg_0);
   assign  _net_384 = (in_do|_reg_0);
   assign  _net_385 = (in_do|_reg_0);
   assign  _net_386 = (in_do|_reg_0);
   assign  _net_387 = (in_do|_reg_0);
   assign  _net_388 = (in_do|_reg_0);
   assign  _net_389 = (in_do|_reg_0);
   assign  _net_390 = (in_do|_reg_0);
   assign  _net_391 = (in_do|_reg_0);
   assign  _net_392 = (in_do|_reg_0);
   assign  _net_393 = (in_do|_reg_0);
   assign  _net_394 = (in_do|_reg_0);
   assign  _net_395 = (in_do|_reg_0);
   assign  _net_396 = (in_do|_reg_0);
   assign  _net_397 = (in_do|_reg_0);
   assign  _net_398 = (in_do|_reg_0);
   assign  _net_399 = (in_do|_reg_0);
   assign  _net_400 = (in_do|_reg_0);
   assign  _net_401 = (in_do|_reg_0);
   assign  _net_402 = (in_do|_reg_0);
   assign  _net_403 = (in_do|_reg_0);
   assign  _net_404 = (in_do|_reg_0);
   assign  _net_405 = (in_do|_reg_0);
   assign  _net_406 = (in_do|_reg_0);
   assign  _net_407 = (in_do|_reg_0);
   assign  _net_408 = (in_do|_reg_0);
   assign  _net_409 = (in_do|_reg_0);
   assign  _net_410 = (in_do|_reg_0);
   assign  _net_411 = (in_do|_reg_0);
   assign  _net_412 = (in_do|_reg_0);
   assign  _net_413 = (in_do|_reg_0);
   assign  _net_414 = (in_do|_reg_0);
   assign  _net_415 = (in_do|_reg_0);
   assign  _net_416 = (in_do|_reg_0);
   assign  _net_417 = (in_do|_reg_0);
   assign  _net_418 = (in_do|_reg_0);
   assign  _net_419 = (in_do|_reg_0);
   assign  _net_420 = (in_do|_reg_0);
   assign  _net_421 = (in_do|_reg_0);

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_seachx_out_do)
    begin
    $display("start %d goal %d",_seachx_startplot,_seachx_goalplot);
    end
  end

// synthesis translate_on
// synopsys translate_on

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
    if(_seachx_out_do)
    begin
    $display("out0=%d",_seachx_data_out33);
    end
  end

// synthesis translate_on
// synopsys translate_on
   assign  kekka_out0 = _kouka_x_loot_out0;
   assign  kekka_out1 = _kouka_x_loot_out1;
   assign  kekka_out2 = _kouka_x_loot_out2;
   assign  kekka_out3 = _kouka_x_loot_out3;
   assign  kekka_out4 = _kouka_x_loot_out4;
   assign  kekka_out5 = _kouka_x_loot_out5;
   assign  kekka_out6 = _kouka_x_loot_out6;
   assign  kekka_out7 = _kouka_x_loot_out7;
   assign  kekka_out8 = _kouka_x_loot_out8;
   assign  kekka_out9 = _kouka_x_loot_out9;
   assign  kekka_out10 = _kouka_x_loot_out10;
   assign  kekka_out11 = _kouka_x_loot_out11;
   assign  kekka_out12 = _kouka_x_loot_out12;
   assign  kekka_out13 = _kouka_x_loot_out13;
   assign  kekka_out14 = _kouka_x_loot_out14;
   assign  kekka_out15 = _kouka_x_loot_out15;
   assign  kekka_out16 = _kouka_x_loot_out16;
   assign  kekka_out17 = _kouka_x_loot_out17;
   assign  kekka_out18 = _kouka_x_loot_out18;
   assign  kekka_out19 = _kouka_x_loot_out19;
   assign  kekka_out20 = _kouka_x_loot_out20;
   assign  kekka_out21 = _kouka_x_loot_out21;
   assign  kekka_out22 = _kouka_x_loot_out22;
   assign  kekka_out23 = _kouka_x_loot_out23;
   assign  kekka_out24 = _kouka_x_loot_out24;
   assign  kekka_out25 = _kouka_x_loot_out25;
   assign  kekka_out26 = _kouka_x_loot_out26;
   assign  kekka_out27 = _kouka_x_loot_out27;
   assign  kekka_out28 = _kouka_x_loot_out28;
   assign  kekka_out29 = _kouka_x_loot_out29;
   assign  kekka_out30 = _kouka_x_loot_out30;
   assign  kekka_out31 = _kouka_x_loot_out31;
   assign  kekka_out32 = _kouka_x_loot_out32;
   assign  kekka_out33 = _kouka_x_loot_out33;
   assign  kekka_out34 = _kouka_x_loot_out34;
   assign  kekka_out35 = _kouka_x_loot_out35;
   assign  kekka_out36 = _kouka_x_loot_out36;
   assign  kekka_out37 = _kouka_x_loot_out37;
   assign  kekka_out38 = _kouka_x_loot_out38;
   assign  kekka_out39 = _kouka_x_loot_out39;
   assign  kekka_out40 = _kouka_x_loot_out40;
   assign  kekka_out41 = _kouka_x_loot_out41;
   assign  kekka_out42 = _kouka_x_loot_out42;
   assign  kekka_out43 = _kouka_x_loot_out43;
   assign  kekka_out44 = _kouka_x_loot_out44;
   assign  kekka_out45 = _kouka_x_loot_out45;
   assign  kekka_out46 = _kouka_x_loot_out46;
   assign  kekka_out47 = _kouka_x_loot_out47;
   assign  kekka_out48 = _kouka_x_loot_out48;
   assign  kekka_out49 = _kouka_x_loot_out49;
   assign  kekka_out50 = _kouka_x_loot_out50;
   assign  kekka_out51 = _kouka_x_loot_out51;
   assign  kekka_out52 = _kouka_x_loot_out52;
   assign  kekka_out53 = _kouka_x_loot_out53;
   assign  kekka_out54 = _kouka_x_loot_out54;
   assign  kekka_out55 = _kouka_x_loot_out55;
   assign  kekka_out56 = _kouka_x_loot_out56;
   assign  kekka_out57 = _kouka_x_loot_out57;
   assign  kekka_out58 = _kouka_x_loot_out58;
   assign  kekka_out59 = _kouka_x_loot_out59;
   assign  kekka_out60 = _kouka_x_loot_out60;
   assign  kekka_out61 = _kouka_x_loot_out61;
   assign  kekka_out62 = _kouka_x_loot_out62;
   assign  kekka_out63 = _kouka_x_loot_out63;
   assign  kekka_out64 = _kouka_x_loot_out64;
   assign  kekka_out65 = _kouka_x_loot_out65;
   assign  kekka_out66 = _kouka_x_loot_out66;
   assign  kekka_out67 = _kouka_x_loot_out67;
   assign  kekka_out68 = _kouka_x_loot_out68;
   assign  kekka_out69 = _kouka_x_loot_out69;
   assign  kekka_out70 = _kouka_x_loot_out70;
   assign  kekka_out71 = _kouka_x_loot_out71;
   assign  kekka_out72 = _kouka_x_loot_out72;
   assign  kekka_out73 = _kouka_x_loot_out73;
   assign  kekka_out74 = _kouka_x_loot_out74;
   assign  kekka_out75 = _kouka_x_loot_out75;
   assign  kekka_out76 = _kouka_x_loot_out76;
   assign  kekka_out77 = _kouka_x_loot_out77;
   assign  kekka_out78 = _kouka_x_loot_out78;
   assign  kekka_out79 = _kouka_x_loot_out79;
   assign  kekka_out80 = _kouka_x_loot_out80;
   assign  kekka_out81 = _kouka_x_loot_out81;
   assign  kekka_out82 = _kouka_x_loot_out82;
   assign  kekka_out83 = _kouka_x_loot_out83;
   assign  kekka_out84 = _kouka_x_loot_out84;
   assign  kekka_out85 = _kouka_x_loot_out85;
   assign  kekka_out86 = _kouka_x_loot_out86;
   assign  kekka_out87 = _kouka_x_loot_out87;
   assign  kekka_out88 = _kouka_x_loot_out88;
   assign  kekka_out89 = _kouka_x_loot_out89;
   assign  kekka_out90 = _kouka_x_loot_out90;
   assign  kekka_out91 = _kouka_x_loot_out91;
   assign  kekka_out92 = _kouka_x_loot_out92;
   assign  kekka_out93 = _kouka_x_loot_out93;
   assign  kekka_out94 = _kouka_x_loot_out94;
   assign  kekka_out95 = _kouka_x_loot_out95;
   assign  kekka_out96 = _kouka_x_loot_out96;
   assign  kekka_out97 = _kouka_x_loot_out97;
   assign  kekka_out98 = _kouka_x_loot_out98;
   assign  kekka_out99 = _kouka_x_loot_out99;
   assign  kekka_out100 = _kouka_x_loot_out100;
   assign  kekka_out101 = _kouka_x_loot_out101;
   assign  kekka_out102 = _kouka_x_loot_out102;
   assign  kekka_out103 = _kouka_x_loot_out103;
   assign  kekka_out104 = _kouka_x_loot_out104;
   assign  kekka_out105 = _kouka_x_loot_out105;
   assign  kekka_out106 = _kouka_x_loot_out106;
   assign  kekka_out107 = _kouka_x_loot_out107;
   assign  kekka_out108 = _kouka_x_loot_out108;
   assign  kekka_out109 = _kouka_x_loot_out109;
   assign  kekka_out110 = _kouka_x_loot_out110;
   assign  kekka_out111 = _kouka_x_loot_out111;
   assign  kekka_out112 = _kouka_x_loot_out112;
   assign  kekka_out113 = _kouka_x_loot_out113;
   assign  kekka_out114 = _kouka_x_loot_out114;
   assign  kekka_out115 = _kouka_x_loot_out115;
   assign  kekka_out116 = _kouka_x_loot_out116;
   assign  kekka_out117 = _kouka_x_loot_out117;
   assign  kekka_out118 = _kouka_x_loot_out118;
   assign  kekka_out119 = _kouka_x_loot_out119;
   assign  kekka_out120 = _kouka_x_loot_out120;
   assign  kekka_out121 = _kouka_x_loot_out121;
   assign  kekka_out122 = _kouka_x_loot_out122;
   assign  kekka_out123 = _kouka_x_loot_out123;
   assign  kekka_out124 = _kouka_x_loot_out124;
   assign  kekka_out125 = _kouka_x_loot_out125;
   assign  kekka_out126 = _kouka_x_loot_out126;
   assign  kekka_out127 = _kouka_x_loot_out127;
   assign  kekka_out128 = _kouka_x_loot_out128;
   assign  kekka_out129 = _kouka_x_loot_out129;
   assign  kekka_out130 = _kouka_x_loot_out130;
   assign  kekka_out131 = _kouka_x_loot_out131;
   assign  kekka_out132 = _kouka_x_loot_out132;
   assign  kekka_out133 = _kouka_x_loot_out133;
   assign  kekka_out134 = _kouka_x_loot_out134;
   assign  kekka_out135 = _kouka_x_loot_out135;
   assign  kekka_out136 = _kouka_x_loot_out136;
   assign  kekka_out137 = _kouka_x_loot_out137;
   assign  kekka_out138 = _kouka_x_loot_out138;
   assign  kekka_out139 = _kouka_x_loot_out139;
   assign  kekka_out140 = _kouka_x_loot_out140;
   assign  kekka_out141 = _kouka_x_loot_out141;
   assign  kekka_out142 = _kouka_x_loot_out142;
   assign  kekka_out143 = _kouka_x_loot_out143;
   assign  kekka_out144 = _kouka_x_loot_out144;
   assign  kekka_out145 = _kouka_x_loot_out145;
   assign  kekka_out146 = _kouka_x_loot_out146;
   assign  kekka_out147 = _kouka_x_loot_out147;
   assign  kekka_out148 = _kouka_x_loot_out148;
   assign  kekka_out149 = _kouka_x_loot_out149;
   assign  kekka_out150 = _kouka_x_loot_out150;
   assign  kekka_out151 = _kouka_x_loot_out151;
   assign  kekka_out152 = _kouka_x_loot_out152;
   assign  kekka_out153 = _kouka_x_loot_out153;
   assign  kekka_out154 = _kouka_x_loot_out154;
   assign  kekka_out155 = _kouka_x_loot_out155;
   assign  kekka_out156 = _kouka_x_loot_out156;
   assign  kekka_out157 = _kouka_x_loot_out157;
   assign  kekka_out158 = _kouka_x_loot_out158;
   assign  kekka_out159 = _kouka_x_loot_out159;
   assign  kekka_out160 = _kouka_x_loot_out160;
   assign  kekka_out161 = _kouka_x_loot_out161;
   assign  kekka_out162 = _kouka_x_loot_out162;
   assign  kekka_out163 = _kouka_x_loot_out163;
   assign  kekka_out164 = _kouka_x_loot_out164;
   assign  kekka_out165 = _kouka_x_loot_out165;
   assign  kekka_out166 = _kouka_x_loot_out166;
   assign  kekka_out167 = _kouka_x_loot_out167;
   assign  kekka_out168 = _kouka_x_loot_out168;
   assign  kekka_out169 = _kouka_x_loot_out169;
   assign  kekka_out170 = _kouka_x_loot_out170;
   assign  kekka_out171 = _kouka_x_loot_out171;
   assign  kekka_out172 = _kouka_x_loot_out172;
   assign  kekka_out173 = _kouka_x_loot_out173;
   assign  kekka_out174 = _kouka_x_loot_out174;
   assign  kekka_out175 = _kouka_x_loot_out175;
   assign  kekka_out176 = _kouka_x_loot_out176;
   assign  kekka_out177 = _kouka_x_loot_out177;
   assign  kekka_out178 = _kouka_x_loot_out178;
   assign  kekka_out179 = _kouka_x_loot_out179;
   assign  kekka_out180 = _kouka_x_loot_out180;
   assign  kekka_out181 = _kouka_x_loot_out181;
   assign  kekka_out182 = _kouka_x_loot_out182;
   assign  kekka_out183 = _kouka_x_loot_out183;
   assign  kekka_out184 = _kouka_x_loot_out184;
   assign  kekka_out185 = _kouka_x_loot_out185;
   assign  kekka_out186 = _kouka_x_loot_out186;
   assign  kekka_out187 = _kouka_x_loot_out187;
   assign  kekka_out188 = _kouka_x_loot_out188;
   assign  kekka_out189 = _kouka_x_loot_out189;
   assign  kekka_out190 = _kouka_x_loot_out190;
   assign  kekka_out191 = _kouka_x_loot_out191;
   assign  kekka_out192 = _kouka_x_loot_out192;
   assign  kekka_out193 = _kouka_x_loot_out193;
   assign  kekka_out194 = _kouka_x_loot_out194;
   assign  kekka_out195 = _kouka_x_loot_out195;
   assign  kekka_out196 = _kouka_x_loot_out196;
   assign  kekka_out197 = _kouka_x_loot_out197;
   assign  kekka_out198 = _kouka_x_loot_out198;
   assign  kekka_out199 = _kouka_x_loot_out199;
   assign  kekka_out200 = _kouka_x_loot_out200;
   assign  kekka_out201 = _kouka_x_loot_out201;
   assign  kekka_out202 = _kouka_x_loot_out202;
   assign  kekka_out203 = _kouka_x_loot_out203;
   assign  kekka_out204 = _kouka_x_loot_out204;
   assign  kekka_out205 = _kouka_x_loot_out205;
   assign  kekka_out206 = _kouka_x_loot_out206;
   assign  kekka_out207 = _kouka_x_loot_out207;
   assign  kekka_out208 = _kouka_x_loot_out208;
   assign  kekka_out209 = _kouka_x_loot_out209;
   assign  kekka_out210 = _kouka_x_loot_out210;
   assign  kekka_out211 = _kouka_x_loot_out211;
   assign  kekka_out212 = _kouka_x_loot_out212;
   assign  kekka_out213 = _kouka_x_loot_out213;
   assign  kekka_out214 = _kouka_x_loot_out214;
   assign  kekka_out215 = _kouka_x_loot_out215;
   assign  kekka_out216 = _kouka_x_loot_out216;
   assign  kekka_out217 = _kouka_x_loot_out217;
   assign  kekka_out218 = _kouka_x_loot_out218;
   assign  kekka_out219 = _kouka_x_loot_out219;
   assign  kekka_out220 = _kouka_x_loot_out220;
   assign  kekka_out221 = _kouka_x_loot_out221;
   assign  kekka_out222 = _kouka_x_loot_out222;
   assign  end_meiro = _kouka_x_out_do;
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     count <= 10'b0000000000;
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_0 <= 1'b0;
else if ((_reg_0)) 
      _reg_0 <= 1'b0;
end
endmodule

/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 14:47:40 2023
 Licensed to :EVALUATION USER*/
