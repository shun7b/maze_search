
/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 14:47:42 2023
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module add_all ( p_reset , m_clock , sig , start , goal , dig_w , data_in33 , data_in34 , data_in35 , data_in36 , data_in37 , data_in38 , data_in39 , data_in40 , data_in41 , data_in42 , data_in43 , data_in44 , data_in45 , data_in46 , data_in47 , data_in48 , data_in49 , data_in50 , data_in51 , data_in52 , data_in53 , data_in54 , data_in55 , data_in56 , data_in57 , data_in58 , data_in59 , data_in60 , data_in61 , data_in62 , data_in65 , data_in66 , data_in67 , data_in68 , data_in69 , data_in70 , data_in71 , data_in72 , data_in73 , data_in74 , data_in75 , data_in76 , data_in77 , data_in78 , data_in79 , data_in80 , data_in81 , data_in82 , data_in83 , data_in84 , data_in85 , data_in86 , data_in87 , data_in88 , data_in89 , data_in90 , data_in91 , data_in92 , data_in93 , data_in94 , data_in97 , data_in98 , data_in99 , data_in100 , data_in101 , data_in102 , data_in103 , data_in104 , data_in105 , data_in106 , data_in107 , data_in108 , data_in109 , data_in110 , data_in111 , data_in112 , data_in113 , data_in114 , data_in115 , data_in116 , data_in117 , data_in118 , data_in119 , data_in120 , data_in121 , data_in122 , data_in123 , data_in124 , data_in125 , data_in126 , data_in129 , data_in130 , data_in131 , data_in132 , data_in133 , data_in134 , data_in135 , data_in136 , data_in137 , data_in138 , data_in139 , data_in140 , data_in141 , data_in142 , data_in143 , data_in144 , data_in145 , data_in146 , data_in147 , data_in148 , data_in149 , data_in150 , data_in151 , data_in152 , data_in153 , data_in154 , data_in155 , data_in156 , data_in157 , data_in158 , data_in161 , data_in162 , data_in163 , data_in164 , data_in165 , data_in166 , data_in167 , data_in168 , data_in169 , data_in170 , data_in171 , data_in172 , data_in173 , data_in174 , data_in175 , data_in176 , data_in177 , data_in178 , data_in179 , data_in180 , data_in181 , data_in182 , data_in183 , data_in184 , data_in185 , data_in186 , data_in187 , data_in188 , data_in189 , data_in190 , data_in193 , data_in194 , data_in195 , data_in196 , data_in197 , data_in198 , data_in199 , data_in200 , data_in201 , data_in202 , data_in203 , data_in204 , data_in205 , data_in206 , data_in207 , data_in208 , data_in209 , data_in210 , data_in211 , data_in212 , data_in213 , data_in214 , data_in215 , data_in216 , data_in217 , data_in218 , data_in219 , data_in220 , data_in221 , data_in222 , data_in225 , data_in226 , data_in227 , data_in228 , data_in229 , data_in230 , data_in231 , data_in232 , data_in233 , data_in234 , data_in235 , data_in236 , data_in237 , data_in238 , data_in239 , data_in240 , data_in241 , data_in242 , data_in243 , data_in244 , data_in245 , data_in246 , data_in247 , data_in248 , data_in249 , data_in250 , data_in251 , data_in252 , data_in253 , data_in254 , data_in257 , data_in258 , data_in259 , data_in260 , data_in261 , data_in262 , data_in263 , data_in264 , data_in265 , data_in266 , data_in267 , data_in268 , data_in269 , data_in270 , data_in271 , data_in272 , data_in273 , data_in274 , data_in275 , data_in276 , data_in277 , data_in278 , data_in279 , data_in280 , data_in281 , data_in282 , data_in283 , data_in284 , data_in285 , data_in286 , data_in289 , data_in290 , data_in291 , data_in292 , data_in293 , data_in294 , data_in295 , data_in296 , data_in297 , data_in298 , data_in299 , data_in300 , data_in301 , data_in302 , data_in303 , data_in304 , data_in305 , data_in306 , data_in307 , data_in308 , data_in309 , data_in310 , data_in311 , data_in312 , data_in313 , data_in314 , data_in315 , data_in316 , data_in317 , data_in318 , data_in321 , data_in322 , data_in323 , data_in324 , data_in325 , data_in326 , data_in327 , data_in328 , data_in329 , data_in330 , data_in331 , data_in332 , data_in333 , data_in334 , data_in335 , data_in336 , data_in337 , data_in338 , data_in339 , data_in340 , data_in341 , data_in342 , data_in343 , data_in344 , data_in345 , data_in346 , data_in347 , data_in348 , data_in349 , data_in350 , data_in353 , data_in354 , data_in355 , data_in356 , data_in357 , data_in358 , data_in359 , data_in360 , data_in361 , data_in362 , data_in363 , data_in364 , data_in365 , data_in366 , data_in367 , data_in368 , data_in369 , data_in370 , data_in371 , data_in372 , data_in373 , data_in374 , data_in375 , data_in376 , data_in377 , data_in378 , data_in379 , data_in380 , data_in381 , data_in382 , data_in385 , data_in386 , data_in387 , data_in388 , data_in389 , data_in390 , data_in391 , data_in392 , data_in393 , data_in394 , data_in395 , data_in396 , data_in397 , data_in398 , data_in399 , data_in400 , data_in401 , data_in402 , data_in403 , data_in404 , data_in405 , data_in406 , data_in407 , data_in408 , data_in409 , data_in410 , data_in411 , data_in412 , data_in413 , data_in414 , data_in417 , data_in418 , data_in419 , data_in420 , data_in421 , data_in422 , data_in423 , data_in424 , data_in425 , data_in426 , data_in427 , data_in428 , data_in429 , data_in430 , data_in431 , data_in432 , data_in433 , data_in434 , data_in435 , data_in436 , data_in437 , data_in438 , data_in439 , data_in440 , data_in441 , data_in442 , data_in443 , data_in444 , data_in445 , data_in446 , data_in449 , data_in450 , data_in451 , data_in452 , data_in453 , data_in454 , data_in455 , data_in456 , data_in457 , data_in458 , data_in459 , data_in460 , data_in461 , data_in462 , data_in463 , data_in464 , data_in465 , data_in466 , data_in467 , data_in468 , data_in469 , data_in470 , data_in471 , data_in472 , data_in473 , data_in474 , data_in475 , data_in476 , data_in477 , data_in478 , data_out_org33 , data_out_org34 , data_out_org35 , data_out_org36 , data_out_org37 , data_out_org38 , data_out_org39 , data_out_org40 , data_out_org41 , data_out_org42 , data_out_org43 , data_out_org44 , data_out_org45 , data_out_org46 , data_out_org47 , data_out_org48 , data_out_org49 , data_out_org50 , data_out_org51 , data_out_org52 , data_out_org53 , data_out_org54 , data_out_org55 , data_out_org56 , data_out_org57 , data_out_org58 , data_out_org59 , data_out_org60 , data_out_org61 , data_out_org62 , data_out_org65 , data_out_org66 , data_out_org67 , data_out_org68 , data_out_org69 , data_out_org70 , data_out_org71 , data_out_org72 , data_out_org73 , data_out_org74 , data_out_org75 , data_out_org76 , data_out_org77 , data_out_org78 , data_out_org79 , data_out_org80 , data_out_org81 , data_out_org82 , data_out_org83 , data_out_org84 , data_out_org85 , data_out_org86 , data_out_org87 , data_out_org88 , data_out_org89 , data_out_org90 , data_out_org91 , data_out_org92 , data_out_org93 , data_out_org94 , data_out_org97 , data_out_org98 , data_out_org99 , data_out_org100 , data_out_org101 , data_out_org102 , data_out_org103 , data_out_org104 , data_out_org105 , data_out_org106 , data_out_org107 , data_out_org108 , data_out_org109 , data_out_org110 , data_out_org111 , data_out_org112 , data_out_org113 , data_out_org114 , data_out_org115 , data_out_org116 , data_out_org117 , data_out_org118 , data_out_org119 , data_out_org120 , data_out_org121 , data_out_org122 , data_out_org123 , data_out_org124 , data_out_org125 , data_out_org126 , data_out_org129 , data_out_org130 , data_out_org131 , data_out_org132 , data_out_org133 , data_out_org134 , data_out_org135 , data_out_org136 , data_out_org137 , data_out_org138 , data_out_org139 , data_out_org140 , data_out_org141 , data_out_org142 , data_out_org143 , data_out_org144 , data_out_org145 , data_out_org146 , data_out_org147 , data_out_org148 , data_out_org149 , data_out_org150 , data_out_org151 , data_out_org152 , data_out_org153 , data_out_org154 , data_out_org155 , data_out_org156 , data_out_org157 , data_out_org158 , data_out_org161 , data_out_org162 , data_out_org163 , data_out_org164 , data_out_org165 , data_out_org166 , data_out_org167 , data_out_org168 , data_out_org169 , data_out_org170 , data_out_org171 , data_out_org172 , data_out_org173 , data_out_org174 , data_out_org175 , data_out_org176 , data_out_org177 , data_out_org178 , data_out_org179 , data_out_org180 , data_out_org181 , data_out_org182 , data_out_org183 , data_out_org184 , data_out_org185 , data_out_org186 , data_out_org187 , data_out_org188 , data_out_org189 , data_out_org190 , data_out_org193 , data_out_org194 , data_out_org195 , data_out_org196 , data_out_org197 , data_out_org198 , data_out_org199 , data_out_org200 , data_out_org201 , data_out_org202 , data_out_org203 , data_out_org204 , data_out_org205 , data_out_org206 , data_out_org207 , data_out_org208 , data_out_org209 , data_out_org210 , data_out_org211 , data_out_org212 , data_out_org213 , data_out_org214 , data_out_org215 , data_out_org216 , data_out_org217 , data_out_org218 , data_out_org219 , data_out_org220 , data_out_org221 , data_out_org222 , data_out_org225 , data_out_org226 , data_out_org227 , data_out_org228 , data_out_org229 , data_out_org230 , data_out_org231 , data_out_org232 , data_out_org233 , data_out_org234 , data_out_org235 , data_out_org236 , data_out_org237 , data_out_org238 , data_out_org239 , data_out_org240 , data_out_org241 , data_out_org242 , data_out_org243 , data_out_org244 , data_out_org245 , data_out_org246 , data_out_org247 , data_out_org248 , data_out_org249 , data_out_org250 , data_out_org251 , data_out_org252 , data_out_org253 , data_out_org254 , data_out_org257 , data_out_org258 , data_out_org259 , data_out_org260 , data_out_org261 , data_out_org262 , data_out_org263 , data_out_org264 , data_out_org265 , data_out_org266 , data_out_org267 , data_out_org268 , data_out_org269 , data_out_org270 , data_out_org271 , data_out_org272 , data_out_org273 , data_out_org274 , data_out_org275 , data_out_org276 , data_out_org277 , data_out_org278 , data_out_org279 , data_out_org280 , data_out_org281 , data_out_org282 , data_out_org283 , data_out_org284 , data_out_org285 , data_out_org286 , data_out_org289 , data_out_org290 , data_out_org291 , data_out_org292 , data_out_org293 , data_out_org294 , data_out_org295 , data_out_org296 , data_out_org297 , data_out_org298 , data_out_org299 , data_out_org300 , data_out_org301 , data_out_org302 , data_out_org303 , data_out_org304 , data_out_org305 , data_out_org306 , data_out_org307 , data_out_org308 , data_out_org309 , data_out_org310 , data_out_org311 , data_out_org312 , data_out_org313 , data_out_org314 , data_out_org315 , data_out_org316 , data_out_org317 , data_out_org318 , data_out_org321 , data_out_org322 , data_out_org323 , data_out_org324 , data_out_org325 , data_out_org326 , data_out_org327 , data_out_org328 , data_out_org329 , data_out_org330 , data_out_org331 , data_out_org332 , data_out_org333 , data_out_org334 , data_out_org335 , data_out_org336 , data_out_org337 , data_out_org338 , data_out_org339 , data_out_org340 , data_out_org341 , data_out_org342 , data_out_org343 , data_out_org344 , data_out_org345 , data_out_org346 , data_out_org347 , data_out_org348 , data_out_org349 , data_out_org350 , data_out_org353 , data_out_org354 , data_out_org355 , data_out_org356 , data_out_org357 , data_out_org358 , data_out_org359 , data_out_org360 , data_out_org361 , data_out_org362 , data_out_org363 , data_out_org364 , data_out_org365 , data_out_org366 , data_out_org367 , data_out_org368 , data_out_org369 , data_out_org370 , data_out_org371 , data_out_org372 , data_out_org373 , data_out_org374 , data_out_org375 , data_out_org376 , data_out_org377 , data_out_org378 , data_out_org379 , data_out_org380 , data_out_org381 , data_out_org382 , data_out_org385 , data_out_org386 , data_out_org387 , data_out_org388 , data_out_org389 , data_out_org390 , data_out_org391 , data_out_org392 , data_out_org393 , data_out_org394 , data_out_org395 , data_out_org396 , data_out_org397 , data_out_org398 , data_out_org399 , data_out_org400 , data_out_org401 , data_out_org402 , data_out_org403 , data_out_org404 , data_out_org405 , data_out_org406 , data_out_org407 , data_out_org408 , data_out_org409 , data_out_org410 , data_out_org411 , data_out_org412 , data_out_org413 , data_out_org414 , data_out_org417 , data_out_org418 , data_out_org419 , data_out_org420 , data_out_org421 , data_out_org422 , data_out_org423 , data_out_org424 , data_out_org425 , data_out_org426 , data_out_org427 , data_out_org428 , data_out_org429 , data_out_org430 , data_out_org431 , data_out_org432 , data_out_org433 , data_out_org434 , data_out_org435 , data_out_org436 , data_out_org437 , data_out_org438 , data_out_org439 , data_out_org440 , data_out_org441 , data_out_org442 , data_out_org443 , data_out_org444 , data_out_org445 , data_out_org446 , data_out_org449 , data_out_org450 , data_out_org451 , data_out_org452 , data_out_org453 , data_out_org454 , data_out_org455 , data_out_org456 , data_out_org457 , data_out_org458 , data_out_org459 , data_out_org460 , data_out_org461 , data_out_org462 , data_out_org463 , data_out_org464 , data_out_org465 , data_out_org466 , data_out_org467 , data_out_org468 , data_out_org469 , data_out_org470 , data_out_org471 , data_out_org472 , data_out_org473 , data_out_org474 , data_out_org475 , data_out_org476 , data_out_org477 , data_out_org478 , data_in_org33 , data_in_org34 , data_in_org35 , data_in_org36 , data_in_org37 , data_in_org38 , data_in_org39 , data_in_org40 , data_in_org41 , data_in_org42 , data_in_org43 , data_in_org44 , data_in_org45 , data_in_org46 , data_in_org47 , data_in_org48 , data_in_org49 , data_in_org50 , data_in_org51 , data_in_org52 , data_in_org53 , data_in_org54 , data_in_org55 , data_in_org56 , data_in_org57 , data_in_org58 , data_in_org59 , data_in_org60 , data_in_org61 , data_in_org62 , data_in_org65 , data_in_org66 , data_in_org67 , data_in_org68 , data_in_org69 , data_in_org70 , data_in_org71 , data_in_org72 , data_in_org73 , data_in_org74 , data_in_org75 , data_in_org76 , data_in_org77 , data_in_org78 , data_in_org79 , data_in_org80 , data_in_org81 , data_in_org82 , data_in_org83 , data_in_org84 , data_in_org85 , data_in_org86 , data_in_org87 , data_in_org88 , data_in_org89 , data_in_org90 , data_in_org91 , data_in_org92 , data_in_org93 , data_in_org94 , data_in_org97 , data_in_org98 , data_in_org99 , data_in_org100 , data_in_org101 , data_in_org102 , data_in_org103 , data_in_org104 , data_in_org105 , data_in_org106 , data_in_org107 , data_in_org108 , data_in_org109 , data_in_org110 , data_in_org111 , data_in_org112 , data_in_org113 , data_in_org114 , data_in_org115 , data_in_org116 , data_in_org117 , data_in_org118 , data_in_org119 , data_in_org120 , data_in_org121 , data_in_org122 , data_in_org123 , data_in_org124 , data_in_org125 , data_in_org126 , data_in_org129 , data_in_org130 , data_in_org131 , data_in_org132 , data_in_org133 , data_in_org134 , data_in_org135 , data_in_org136 , data_in_org137 , data_in_org138 , data_in_org139 , data_in_org140 , data_in_org141 , data_in_org142 , data_in_org143 , data_in_org144 , data_in_org145 , data_in_org146 , data_in_org147 , data_in_org148 , data_in_org149 , data_in_org150 , data_in_org151 , data_in_org152 , data_in_org153 , data_in_org154 , data_in_org155 , data_in_org156 , data_in_org157 , data_in_org158 , data_in_org161 , data_in_org162 , data_in_org163 , data_in_org164 , data_in_org165 , data_in_org166 , data_in_org167 , data_in_org168 , data_in_org169 , data_in_org170 , data_in_org171 , data_in_org172 , data_in_org173 , data_in_org174 , data_in_org175 , data_in_org176 , data_in_org177 , data_in_org178 , data_in_org179 , data_in_org180 , data_in_org181 , data_in_org182 , data_in_org183 , data_in_org184 , data_in_org185 , data_in_org186 , data_in_org187 , data_in_org188 , data_in_org189 , data_in_org190 , data_in_org193 , data_in_org194 , data_in_org195 , data_in_org196 , data_in_org197 , data_in_org198 , data_in_org199 , data_in_org200 , data_in_org201 , data_in_org202 , data_in_org203 , data_in_org204 , data_in_org205 , data_in_org206 , data_in_org207 , data_in_org208 , data_in_org209 , data_in_org210 , data_in_org211 , data_in_org212 , data_in_org213 , data_in_org214 , data_in_org215 , data_in_org216 , data_in_org217 , data_in_org218 , data_in_org219 , data_in_org220 , data_in_org221 , data_in_org222 , data_in_org225 , data_in_org226 , data_in_org227 , data_in_org228 , data_in_org229 , data_in_org230 , data_in_org231 , data_in_org232 , data_in_org233 , data_in_org234 , data_in_org235 , data_in_org236 , data_in_org237 , data_in_org238 , data_in_org239 , data_in_org240 , data_in_org241 , data_in_org242 , data_in_org243 , data_in_org244 , data_in_org245 , data_in_org246 , data_in_org247 , data_in_org248 , data_in_org249 , data_in_org250 , data_in_org251 , data_in_org252 , data_in_org253 , data_in_org254 , data_in_org257 , data_in_org258 , data_in_org259 , data_in_org260 , data_in_org261 , data_in_org262 , data_in_org263 , data_in_org264 , data_in_org265 , data_in_org266 , data_in_org267 , data_in_org268 , data_in_org269 , data_in_org270 , data_in_org271 , data_in_org272 , data_in_org273 , data_in_org274 , data_in_org275 , data_in_org276 , data_in_org277 , data_in_org278 , data_in_org279 , data_in_org280 , data_in_org281 , data_in_org282 , data_in_org283 , data_in_org284 , data_in_org285 , data_in_org286 , data_in_org289 , data_in_org290 , data_in_org291 , data_in_org292 , data_in_org293 , data_in_org294 , data_in_org295 , data_in_org296 , data_in_org297 , data_in_org298 , data_in_org299 , data_in_org300 , data_in_org301 , data_in_org302 , data_in_org303 , data_in_org304 , data_in_org305 , data_in_org306 , data_in_org307 , data_in_org308 , data_in_org309 , data_in_org310 , data_in_org311 , data_in_org312 , data_in_org313 , data_in_org314 , data_in_org315 , data_in_org316 , data_in_org317 , data_in_org318 , data_in_org321 , data_in_org322 , data_in_org323 , data_in_org324 , data_in_org325 , data_in_org326 , data_in_org327 , data_in_org328 , data_in_org329 , data_in_org330 , data_in_org331 , data_in_org332 , data_in_org333 , data_in_org334 , data_in_org335 , data_in_org336 , data_in_org337 , data_in_org338 , data_in_org339 , data_in_org340 , data_in_org341 , data_in_org342 , data_in_org343 , data_in_org344 , data_in_org345 , data_in_org346 , data_in_org347 , data_in_org348 , data_in_org349 , data_in_org350 , data_in_org353 , data_in_org354 , data_in_org355 , data_in_org356 , data_in_org357 , data_in_org358 , data_in_org359 , data_in_org360 , data_in_org361 , data_in_org362 , data_in_org363 , data_in_org364 , data_in_org365 , data_in_org366 , data_in_org367 , data_in_org368 , data_in_org369 , data_in_org370 , data_in_org371 , data_in_org372 , data_in_org373 , data_in_org374 , data_in_org375 , data_in_org376 , data_in_org377 , data_in_org378 , data_in_org379 , data_in_org380 , data_in_org381 , data_in_org382 , data_in_org385 , data_in_org386 , data_in_org387 , data_in_org388 , data_in_org389 , data_in_org390 , data_in_org391 , data_in_org392 , data_in_org393 , data_in_org394 , data_in_org395 , data_in_org396 , data_in_org397 , data_in_org398 , data_in_org399 , data_in_org400 , data_in_org401 , data_in_org402 , data_in_org403 , data_in_org404 , data_in_org405 , data_in_org406 , data_in_org407 , data_in_org408 , data_in_org409 , data_in_org410 , data_in_org411 , data_in_org412 , data_in_org413 , data_in_org414 , data_in_org417 , data_in_org418 , data_in_org419 , data_in_org420 , data_in_org421 , data_in_org422 , data_in_org423 , data_in_org424 , data_in_org425 , data_in_org426 , data_in_org427 , data_in_org428 , data_in_org429 , data_in_org430 , data_in_org431 , data_in_org432 , data_in_org433 , data_in_org434 , data_in_org435 , data_in_org436 , data_in_org437 , data_in_org438 , data_in_org439 , data_in_org440 , data_in_org441 , data_in_org442 , data_in_org443 , data_in_org444 , data_in_org445 , data_in_org446 , data_in_org449 , data_in_org450 , data_in_org451 , data_in_org452 , data_in_org453 , data_in_org454 , data_in_org455 , data_in_org456 , data_in_org457 , data_in_org458 , data_in_org459 , data_in_org460 , data_in_org461 , data_in_org462 , data_in_org463 , data_in_org464 , data_in_org465 , data_in_org466 , data_in_org467 , data_in_org468 , data_in_org469 , data_in_org470 , data_in_org471 , data_in_org472 , data_in_org473 , data_in_org474 , data_in_org475 , data_in_org476 , data_in_org477 , data_in_org478 , data_out33 , data_out34 , data_out35 , data_out36 , data_out37 , data_out38 , data_out39 , data_out40 , data_out41 , data_out42 , data_out43 , data_out44 , data_out45 , data_out46 , data_out47 , data_out48 , data_out49 , data_out50 , data_out51 , data_out52 , data_out53 , data_out54 , data_out55 , data_out56 , data_out57 , data_out58 , data_out59 , data_out60 , data_out61 , data_out62 , data_out65 , data_out66 , data_out67 , data_out68 , data_out69 , data_out70 , data_out71 , data_out72 , data_out73 , data_out74 , data_out75 , data_out76 , data_out77 , data_out78 , data_out79 , data_out80 , data_out81 , data_out82 , data_out83 , data_out84 , data_out85 , data_out86 , data_out87 , data_out88 , data_out89 , data_out90 , data_out91 , data_out92 , data_out93 , data_out94 , data_out97 , data_out98 , data_out99 , data_out100 , data_out101 , data_out102 , data_out103 , data_out104 , data_out105 , data_out106 , data_out107 , data_out108 , data_out109 , data_out110 , data_out111 , data_out112 , data_out113 , data_out114 , data_out115 , data_out116 , data_out117 , data_out118 , data_out119 , data_out120 , data_out121 , data_out122 , data_out123 , data_out124 , data_out125 , data_out126 , data_out129 , data_out130 , data_out131 , data_out132 , data_out133 , data_out134 , data_out135 , data_out136 , data_out137 , data_out138 , data_out139 , data_out140 , data_out141 , data_out142 , data_out143 , data_out144 , data_out145 , data_out146 , data_out147 , data_out148 , data_out149 , data_out150 , data_out151 , data_out152 , data_out153 , data_out154 , data_out155 , data_out156 , data_out157 , data_out158 , data_out161 , data_out162 , data_out163 , data_out164 , data_out165 , data_out166 , data_out167 , data_out168 , data_out169 , data_out170 , data_out171 , data_out172 , data_out173 , data_out174 , data_out175 , data_out176 , data_out177 , data_out178 , data_out179 , data_out180 , data_out181 , data_out182 , data_out183 , data_out184 , data_out185 , data_out186 , data_out187 , data_out188 , data_out189 , data_out190 , data_out193 , data_out194 , data_out195 , data_out196 , data_out197 , data_out198 , data_out199 , data_out200 , data_out201 , data_out202 , data_out203 , data_out204 , data_out205 , data_out206 , data_out207 , data_out208 , data_out209 , data_out210 , data_out211 , data_out212 , data_out213 , data_out214 , data_out215 , data_out216 , data_out217 , data_out218 , data_out219 , data_out220 , data_out221 , data_out222 , data_out225 , data_out226 , data_out227 , data_out228 , data_out229 , data_out230 , data_out231 , data_out232 , data_out233 , data_out234 , data_out235 , data_out236 , data_out237 , data_out238 , data_out239 , data_out240 , data_out241 , data_out242 , data_out243 , data_out244 , data_out245 , data_out246 , data_out247 , data_out248 , data_out249 , data_out250 , data_out251 , data_out252 , data_out253 , data_out254 , data_out257 , data_out258 , data_out259 , data_out260 , data_out261 , data_out262 , data_out263 , data_out264 , data_out265 , data_out266 , data_out267 , data_out268 , data_out269 , data_out270 , data_out271 , data_out272 , data_out273 , data_out274 , data_out275 , data_out276 , data_out277 , data_out278 , data_out279 , data_out280 , data_out281 , data_out282 , data_out283 , data_out284 , data_out285 , data_out286 , data_out289 , data_out290 , data_out291 , data_out292 , data_out293 , data_out294 , data_out295 , data_out296 , data_out297 , data_out298 , data_out299 , data_out300 , data_out301 , data_out302 , data_out303 , data_out304 , data_out305 , data_out306 , data_out307 , data_out308 , data_out309 , data_out310 , data_out311 , data_out312 , data_out313 , data_out314 , data_out315 , data_out316 , data_out317 , data_out318 , data_out321 , data_out322 , data_out323 , data_out324 , data_out325 , data_out326 , data_out327 , data_out328 , data_out329 , data_out330 , data_out331 , data_out332 , data_out333 , data_out334 , data_out335 , data_out336 , data_out337 , data_out338 , data_out339 , data_out340 , data_out341 , data_out342 , data_out343 , data_out344 , data_out345 , data_out346 , data_out347 , data_out348 , data_out349 , data_out350 , data_out353 , data_out354 , data_out355 , data_out356 , data_out357 , data_out358 , data_out359 , data_out360 , data_out361 , data_out362 , data_out363 , data_out364 , data_out365 , data_out366 , data_out367 , data_out368 , data_out369 , data_out370 , data_out371 , data_out372 , data_out373 , data_out374 , data_out375 , data_out376 , data_out377 , data_out378 , data_out379 , data_out380 , data_out381 , data_out382 , data_out385 , data_out386 , data_out387 , data_out388 , data_out389 , data_out390 , data_out391 , data_out392 , data_out393 , data_out394 , data_out395 , data_out396 , data_out397 , data_out398 , data_out399 , data_out400 , data_out401 , data_out402 , data_out403 , data_out404 , data_out405 , data_out406 , data_out407 , data_out408 , data_out409 , data_out410 , data_out411 , data_out412 , data_out413 , data_out414 , data_out417 , data_out418 , data_out419 , data_out420 , data_out421 , data_out422 , data_out423 , data_out424 , data_out425 , data_out426 , data_out427 , data_out428 , data_out429 , data_out430 , data_out431 , data_out432 , data_out433 , data_out434 , data_out435 , data_out436 , data_out437 , data_out438 , data_out439 , data_out440 , data_out441 , data_out442 , data_out443 , data_out444 , data_out445 , data_out446 , data_out449 , data_out450 , data_out451 , data_out452 , data_out453 , data_out454 , data_out455 , data_out456 , data_out457 , data_out458 , data_out459 , data_out460 , data_out461 , data_out462 , data_out463 , data_out464 , data_out465 , data_out466 , data_out467 , data_out468 , data_out469 , data_out470 , data_out471 , data_out472 , data_out473 , data_out474 , data_out475 , data_out476 , data_out477 , data_out478 , data_out_index33 , data_out_index34 , data_out_index35 , data_out_index36 , data_out_index37 , data_out_index38 , data_out_index39 , data_out_index40 , data_out_index41 , data_out_index42 , data_out_index43 , data_out_index44 , data_out_index45 , data_out_index46 , data_out_index47 , data_out_index48 , data_out_index49 , data_out_index50 , data_out_index51 , data_out_index52 , data_out_index53 , data_out_index54 , data_out_index55 , data_out_index56 , data_out_index57 , data_out_index58 , data_out_index59 , data_out_index60 , data_out_index61 , data_out_index62 , data_out_index65 , data_out_index66 , data_out_index67 , data_out_index68 , data_out_index69 , data_out_index70 , data_out_index71 , data_out_index72 , data_out_index73 , data_out_index74 , data_out_index75 , data_out_index76 , data_out_index77 , data_out_index78 , data_out_index79 , data_out_index80 , data_out_index81 , data_out_index82 , data_out_index83 , data_out_index84 , data_out_index85 , data_out_index86 , data_out_index87 , data_out_index88 , data_out_index89 , data_out_index90 , data_out_index91 , data_out_index92 , data_out_index93 , data_out_index94 , data_out_index97 , data_out_index98 , data_out_index99 , data_out_index100 , data_out_index101 , data_out_index102 , data_out_index103 , data_out_index104 , data_out_index105 , data_out_index106 , data_out_index107 , data_out_index108 , data_out_index109 , data_out_index110 , data_out_index111 , data_out_index112 , data_out_index113 , data_out_index114 , data_out_index115 , data_out_index116 , data_out_index117 , data_out_index118 , data_out_index119 , data_out_index120 , data_out_index121 , data_out_index122 , data_out_index123 , data_out_index124 , data_out_index125 , data_out_index126 , data_out_index129 , data_out_index130 , data_out_index131 , data_out_index132 , data_out_index133 , data_out_index134 , data_out_index135 , data_out_index136 , data_out_index137 , data_out_index138 , data_out_index139 , data_out_index140 , data_out_index141 , data_out_index142 , data_out_index143 , data_out_index144 , data_out_index145 , data_out_index146 , data_out_index147 , data_out_index148 , data_out_index149 , data_out_index150 , data_out_index151 , data_out_index152 , data_out_index153 , data_out_index154 , data_out_index155 , data_out_index156 , data_out_index157 , data_out_index158 , data_out_index161 , data_out_index162 , data_out_index163 , data_out_index164 , data_out_index165 , data_out_index166 , data_out_index167 , data_out_index168 , data_out_index169 , data_out_index170 , data_out_index171 , data_out_index172 , data_out_index173 , data_out_index174 , data_out_index175 , data_out_index176 , data_out_index177 , data_out_index178 , data_out_index179 , data_out_index180 , data_out_index181 , data_out_index182 , data_out_index183 , data_out_index184 , data_out_index185 , data_out_index186 , data_out_index187 , data_out_index188 , data_out_index189 , data_out_index190 , data_out_index193 , data_out_index194 , data_out_index195 , data_out_index196 , data_out_index197 , data_out_index198 , data_out_index199 , data_out_index200 , data_out_index201 , data_out_index202 , data_out_index203 , data_out_index204 , data_out_index205 , data_out_index206 , data_out_index207 , data_out_index208 , data_out_index209 , data_out_index210 , data_out_index211 , data_out_index212 , data_out_index213 , data_out_index214 , data_out_index215 , data_out_index216 , data_out_index217 , data_out_index218 , data_out_index219 , data_out_index220 , data_out_index221 , data_out_index222 , data_out_index225 , data_out_index226 , data_out_index227 , data_out_index228 , data_out_index229 , data_out_index230 , data_out_index231 , data_out_index232 , data_out_index233 , data_out_index234 , data_out_index235 , data_out_index236 , data_out_index237 , data_out_index238 , data_out_index239 , data_out_index240 , data_out_index241 , data_out_index242 , data_out_index243 , data_out_index244 , data_out_index245 , data_out_index246 , data_out_index247 , data_out_index248 , data_out_index249 , data_out_index250 , data_out_index251 , data_out_index252 , data_out_index253 , data_out_index254 , data_out_index257 , data_out_index258 , data_out_index259 , data_out_index260 , data_out_index261 , data_out_index262 , data_out_index263 , data_out_index264 , data_out_index265 , data_out_index266 , data_out_index267 , data_out_index268 , data_out_index269 , data_out_index270 , data_out_index271 , data_out_index272 , data_out_index273 , data_out_index274 , data_out_index275 , data_out_index276 , data_out_index277 , data_out_index278 , data_out_index279 , data_out_index280 , data_out_index281 , data_out_index282 , data_out_index283 , data_out_index284 , data_out_index285 , data_out_index286 , data_out_index289 , data_out_index290 , data_out_index291 , data_out_index292 , data_out_index293 , data_out_index294 , data_out_index295 , data_out_index296 , data_out_index297 , data_out_index298 , data_out_index299 , data_out_index300 , data_out_index301 , data_out_index302 , data_out_index303 , data_out_index304 , data_out_index305 , data_out_index306 , data_out_index307 , data_out_index308 , data_out_index309 , data_out_index310 , data_out_index311 , data_out_index312 , data_out_index313 , data_out_index314 , data_out_index315 , data_out_index316 , data_out_index317 , data_out_index318 , data_out_index321 , data_out_index322 , data_out_index323 , data_out_index324 , data_out_index325 , data_out_index326 , data_out_index327 , data_out_index328 , data_out_index329 , data_out_index330 , data_out_index331 , data_out_index332 , data_out_index333 , data_out_index334 , data_out_index335 , data_out_index336 , data_out_index337 , data_out_index338 , data_out_index339 , data_out_index340 , data_out_index341 , data_out_index342 , data_out_index343 , data_out_index344 , data_out_index345 , data_out_index346 , data_out_index347 , data_out_index348 , data_out_index349 , data_out_index350 , data_out_index353 , data_out_index354 , data_out_index355 , data_out_index356 , data_out_index357 , data_out_index358 , data_out_index359 , data_out_index360 , data_out_index361 , data_out_index362 , data_out_index363 , data_out_index364 , data_out_index365 , data_out_index366 , data_out_index367 , data_out_index368 , data_out_index369 , data_out_index370 , data_out_index371 , data_out_index372 , data_out_index373 , data_out_index374 , data_out_index375 , data_out_index376 , data_out_index377 , data_out_index378 , data_out_index379 , data_out_index380 , data_out_index381 , data_out_index382 , data_out_index385 , data_out_index386 , data_out_index387 , data_out_index388 , data_out_index389 , data_out_index390 , data_out_index391 , data_out_index392 , data_out_index393 , data_out_index394 , data_out_index395 , data_out_index396 , data_out_index397 , data_out_index398 , data_out_index399 , data_out_index400 , data_out_index401 , data_out_index402 , data_out_index403 , data_out_index404 , data_out_index405 , data_out_index406 , data_out_index407 , data_out_index408 , data_out_index409 , data_out_index410 , data_out_index411 , data_out_index412 , data_out_index413 , data_out_index414 , data_out_index417 , data_out_index418 , data_out_index419 , data_out_index420 , data_out_index421 , data_out_index422 , data_out_index423 , data_out_index424 , data_out_index425 , data_out_index426 , data_out_index427 , data_out_index428 , data_out_index429 , data_out_index430 , data_out_index431 , data_out_index432 , data_out_index433 , data_out_index434 , data_out_index435 , data_out_index436 , data_out_index437 , data_out_index438 , data_out_index439 , data_out_index440 , data_out_index441 , data_out_index442 , data_out_index443 , data_out_index444 , data_out_index445 , data_out_index446 , data_out_index449 , data_out_index450 , data_out_index451 , data_out_index452 , data_out_index453 , data_out_index454 , data_out_index455 , data_out_index456 , data_out_index457 , data_out_index458 , data_out_index459 , data_out_index460 , data_out_index461 , data_out_index462 , data_out_index463 , data_out_index464 , data_out_index465 , data_out_index466 , data_out_index467 , data_out_index468 , data_out_index469 , data_out_index470 , data_out_index471 , data_out_index472 , data_out_index473 , data_out_index474 , data_out_index475 , data_out_index476 , data_out_index477 , data_out_index478 , sg_in33 , sg_in34 , sg_in35 , sg_in36 , sg_in37 , sg_in38 , sg_in39 , sg_in40 , sg_in41 , sg_in42 , sg_in43 , sg_in44 , sg_in45 , sg_in46 , sg_in47 , sg_in48 , sg_in49 , sg_in50 , sg_in51 , sg_in52 , sg_in53 , sg_in54 , sg_in55 , sg_in56 , sg_in57 , sg_in58 , sg_in59 , sg_in60 , sg_in61 , sg_in62 , sg_in65 , sg_in66 , sg_in67 , sg_in68 , sg_in69 , sg_in70 , sg_in71 , sg_in72 , sg_in73 , sg_in74 , sg_in75 , sg_in76 , sg_in77 , sg_in78 , sg_in79 , sg_in80 , sg_in81 , sg_in82 , sg_in83 , sg_in84 , sg_in85 , sg_in86 , sg_in87 , sg_in88 , sg_in89 , sg_in90 , sg_in91 , sg_in92 , sg_in93 , sg_in94 , sg_in97 , sg_in98 , sg_in99 , sg_in100 , sg_in101 , sg_in102 , sg_in103 , sg_in104 , sg_in105 , sg_in106 , sg_in107 , sg_in108 , sg_in109 , sg_in110 , sg_in111 , sg_in112 , sg_in113 , sg_in114 , sg_in115 , sg_in116 , sg_in117 , sg_in118 , sg_in119 , sg_in120 , sg_in121 , sg_in122 , sg_in123 , sg_in124 , sg_in125 , sg_in126 , sg_in129 , sg_in130 , sg_in131 , sg_in132 , sg_in133 , sg_in134 , sg_in135 , sg_in136 , sg_in137 , sg_in138 , sg_in139 , sg_in140 , sg_in141 , sg_in142 , sg_in143 , sg_in144 , sg_in145 , sg_in146 , sg_in147 , sg_in148 , sg_in149 , sg_in150 , sg_in151 , sg_in152 , sg_in153 , sg_in154 , sg_in155 , sg_in156 , sg_in157 , sg_in158 , sg_in161 , sg_in162 , sg_in163 , sg_in164 , sg_in165 , sg_in166 , sg_in167 , sg_in168 , sg_in169 , sg_in170 , sg_in171 , sg_in172 , sg_in173 , sg_in174 , sg_in175 , sg_in176 , sg_in177 , sg_in178 , sg_in179 , sg_in180 , sg_in181 , sg_in182 , sg_in183 , sg_in184 , sg_in185 , sg_in186 , sg_in187 , sg_in188 , sg_in189 , sg_in190 , sg_in193 , sg_in194 , sg_in195 , sg_in196 , sg_in197 , sg_in198 , sg_in199 , sg_in200 , sg_in201 , sg_in202 , sg_in203 , sg_in204 , sg_in205 , sg_in206 , sg_in207 , sg_in208 , sg_in209 , sg_in210 , sg_in211 , sg_in212 , sg_in213 , sg_in214 , sg_in215 , sg_in216 , sg_in217 , sg_in218 , sg_in219 , sg_in220 , sg_in221 , sg_in222 , sg_in225 , sg_in226 , sg_in227 , sg_in228 , sg_in229 , sg_in230 , sg_in231 , sg_in232 , sg_in233 , sg_in234 , sg_in235 , sg_in236 , sg_in237 , sg_in238 , sg_in239 , sg_in240 , sg_in241 , sg_in242 , sg_in243 , sg_in244 , sg_in245 , sg_in246 , sg_in247 , sg_in248 , sg_in249 , sg_in250 , sg_in251 , sg_in252 , sg_in253 , sg_in254 , sg_in257 , sg_in258 , sg_in259 , sg_in260 , sg_in261 , sg_in262 , sg_in263 , sg_in264 , sg_in265 , sg_in266 , sg_in267 , sg_in268 , sg_in269 , sg_in270 , sg_in271 , sg_in272 , sg_in273 , sg_in274 , sg_in275 , sg_in276 , sg_in277 , sg_in278 , sg_in279 , sg_in280 , sg_in281 , sg_in282 , sg_in283 , sg_in284 , sg_in285 , sg_in286 , sg_in289 , sg_in290 , sg_in291 , sg_in292 , sg_in293 , sg_in294 , sg_in295 , sg_in296 , sg_in297 , sg_in298 , sg_in299 , sg_in300 , sg_in301 , sg_in302 , sg_in303 , sg_in304 , sg_in305 , sg_in306 , sg_in307 , sg_in308 , sg_in309 , sg_in310 , sg_in311 , sg_in312 , sg_in313 , sg_in314 , sg_in315 , sg_in316 , sg_in317 , sg_in318 , sg_in321 , sg_in322 , sg_in323 , sg_in324 , sg_in325 , sg_in326 , sg_in327 , sg_in328 , sg_in329 , sg_in330 , sg_in331 , sg_in332 , sg_in333 , sg_in334 , sg_in335 , sg_in336 , sg_in337 , sg_in338 , sg_in339 , sg_in340 , sg_in341 , sg_in342 , sg_in343 , sg_in344 , sg_in345 , sg_in346 , sg_in347 , sg_in348 , sg_in349 , sg_in350 , sg_in353 , sg_in354 , sg_in355 , sg_in356 , sg_in357 , sg_in358 , sg_in359 , sg_in360 , sg_in361 , sg_in362 , sg_in363 , sg_in364 , sg_in365 , sg_in366 , sg_in367 , sg_in368 , sg_in369 , sg_in370 , sg_in371 , sg_in372 , sg_in373 , sg_in374 , sg_in375 , sg_in376 , sg_in377 , sg_in378 , sg_in379 , sg_in380 , sg_in381 , sg_in382 , sg_in385 , sg_in386 , sg_in387 , sg_in388 , sg_in389 , sg_in390 , sg_in391 , sg_in392 , sg_in393 , sg_in394 , sg_in395 , sg_in396 , sg_in397 , sg_in398 , sg_in399 , sg_in400 , sg_in401 , sg_in402 , sg_in403 , sg_in404 , sg_in405 , sg_in406 , sg_in407 , sg_in408 , sg_in409 , sg_in410 , sg_in411 , sg_in412 , sg_in413 , sg_in414 , sg_in417 , sg_in418 , sg_in419 , sg_in420 , sg_in421 , sg_in422 , sg_in423 , sg_in424 , sg_in425 , sg_in426 , sg_in427 , sg_in428 , sg_in429 , sg_in430 , sg_in431 , sg_in432 , sg_in433 , sg_in434 , sg_in435 , sg_in436 , sg_in437 , sg_in438 , sg_in439 , sg_in440 , sg_in441 , sg_in442 , sg_in443 , sg_in444 , sg_in445 , sg_in446 , sg_in449 , sg_in450 , sg_in451 , sg_in452 , sg_in453 , sg_in454 , sg_in455 , sg_in456 , sg_in457 , sg_in458 , sg_in459 , sg_in460 , sg_in461 , sg_in462 , sg_in463 , sg_in464 , sg_in465 , sg_in466 , sg_in467 , sg_in468 , sg_in469 , sg_in470 , sg_in471 , sg_in472 , sg_in473 , sg_in474 , sg_in475 , sg_in476 , sg_in477 , sg_in478 , sg_out33 , sg_out34 , sg_out35 , sg_out36 , sg_out37 , sg_out38 , sg_out39 , sg_out40 , sg_out41 , sg_out42 , sg_out43 , sg_out44 , sg_out45 , sg_out46 , sg_out47 , sg_out48 , sg_out49 , sg_out50 , sg_out51 , sg_out52 , sg_out53 , sg_out54 , sg_out55 , sg_out56 , sg_out57 , sg_out58 , sg_out59 , sg_out60 , sg_out61 , sg_out62 , sg_out65 , sg_out66 , sg_out67 , sg_out68 , sg_out69 , sg_out70 , sg_out71 , sg_out72 , sg_out73 , sg_out74 , sg_out75 , sg_out76 , sg_out77 , sg_out78 , sg_out79 , sg_out80 , sg_out81 , sg_out82 , sg_out83 , sg_out84 , sg_out85 , sg_out86 , sg_out87 , sg_out88 , sg_out89 , sg_out90 , sg_out91 , sg_out92 , sg_out93 , sg_out94 , sg_out97 , sg_out98 , sg_out99 , sg_out100 , sg_out101 , sg_out102 , sg_out103 , sg_out104 , sg_out105 , sg_out106 , sg_out107 , sg_out108 , sg_out109 , sg_out110 , sg_out111 , sg_out112 , sg_out113 , sg_out114 , sg_out115 , sg_out116 , sg_out117 , sg_out118 , sg_out119 , sg_out120 , sg_out121 , sg_out122 , sg_out123 , sg_out124 , sg_out125 , sg_out126 , sg_out129 , sg_out130 , sg_out131 , sg_out132 , sg_out133 , sg_out134 , sg_out135 , sg_out136 , sg_out137 , sg_out138 , sg_out139 , sg_out140 , sg_out141 , sg_out142 , sg_out143 , sg_out144 , sg_out145 , sg_out146 , sg_out147 , sg_out148 , sg_out149 , sg_out150 , sg_out151 , sg_out152 , sg_out153 , sg_out154 , sg_out155 , sg_out156 , sg_out157 , sg_out158 , sg_out161 , sg_out162 , sg_out163 , sg_out164 , sg_out165 , sg_out166 , sg_out167 , sg_out168 , sg_out169 , sg_out170 , sg_out171 , sg_out172 , sg_out173 , sg_out174 , sg_out175 , sg_out176 , sg_out177 , sg_out178 , sg_out179 , sg_out180 , sg_out181 , sg_out182 , sg_out183 , sg_out184 , sg_out185 , sg_out186 , sg_out187 , sg_out188 , sg_out189 , sg_out190 , sg_out193 , sg_out194 , sg_out195 , sg_out196 , sg_out197 , sg_out198 , sg_out199 , sg_out200 , sg_out201 , sg_out202 , sg_out203 , sg_out204 , sg_out205 , sg_out206 , sg_out207 , sg_out208 , sg_out209 , sg_out210 , sg_out211 , sg_out212 , sg_out213 , sg_out214 , sg_out215 , sg_out216 , sg_out217 , sg_out218 , sg_out219 , sg_out220 , sg_out221 , sg_out222 , sg_out225 , sg_out226 , sg_out227 , sg_out228 , sg_out229 , sg_out230 , sg_out231 , sg_out232 , sg_out233 , sg_out234 , sg_out235 , sg_out236 , sg_out237 , sg_out238 , sg_out239 , sg_out240 , sg_out241 , sg_out242 , sg_out243 , sg_out244 , sg_out245 , sg_out246 , sg_out247 , sg_out248 , sg_out249 , sg_out250 , sg_out251 , sg_out252 , sg_out253 , sg_out254 , sg_out257 , sg_out258 , sg_out259 , sg_out260 , sg_out261 , sg_out262 , sg_out263 , sg_out264 , sg_out265 , sg_out266 , sg_out267 , sg_out268 , sg_out269 , sg_out270 , sg_out271 , sg_out272 , sg_out273 , sg_out274 , sg_out275 , sg_out276 , sg_out277 , sg_out278 , sg_out279 , sg_out280 , sg_out281 , sg_out282 , sg_out283 , sg_out284 , sg_out285 , sg_out286 , sg_out289 , sg_out290 , sg_out291 , sg_out292 , sg_out293 , sg_out294 , sg_out295 , sg_out296 , sg_out297 , sg_out298 , sg_out299 , sg_out300 , sg_out301 , sg_out302 , sg_out303 , sg_out304 , sg_out305 , sg_out306 , sg_out307 , sg_out308 , sg_out309 , sg_out310 , sg_out311 , sg_out312 , sg_out313 , sg_out314 , sg_out315 , sg_out316 , sg_out317 , sg_out318 , sg_out321 , sg_out322 , sg_out323 , sg_out324 , sg_out325 , sg_out326 , sg_out327 , sg_out328 , sg_out329 , sg_out330 , sg_out331 , sg_out332 , sg_out333 , sg_out334 , sg_out335 , sg_out336 , sg_out337 , sg_out338 , sg_out339 , sg_out340 , sg_out341 , sg_out342 , sg_out343 , sg_out344 , sg_out345 , sg_out346 , sg_out347 , sg_out348 , sg_out349 , sg_out350 , sg_out353 , sg_out354 , sg_out355 , sg_out356 , sg_out357 , sg_out358 , sg_out359 , sg_out360 , sg_out361 , sg_out362 , sg_out363 , sg_out364 , sg_out365 , sg_out366 , sg_out367 , sg_out368 , sg_out369 , sg_out370 , sg_out371 , sg_out372 , sg_out373 , sg_out374 , sg_out375 , sg_out376 , sg_out377 , sg_out378 , sg_out379 , sg_out380 , sg_out381 , sg_out382 , sg_out385 , sg_out386 , sg_out387 , sg_out388 , sg_out389 , sg_out390 , sg_out391 , sg_out392 , sg_out393 , sg_out394 , sg_out395 , sg_out396 , sg_out397 , sg_out398 , sg_out399 , sg_out400 , sg_out401 , sg_out402 , sg_out403 , sg_out404 , sg_out405 , sg_out406 , sg_out407 , sg_out408 , sg_out409 , sg_out410 , sg_out411 , sg_out412 , sg_out413 , sg_out414 , sg_out417 , sg_out418 , sg_out419 , sg_out420 , sg_out421 , sg_out422 , sg_out423 , sg_out424 , sg_out425 , sg_out426 , sg_out427 , sg_out428 , sg_out429 , sg_out430 , sg_out431 , sg_out432 , sg_out433 , sg_out434 , sg_out435 , sg_out436 , sg_out437 , sg_out438 , sg_out439 , sg_out440 , sg_out441 , sg_out442 , sg_out443 , sg_out444 , sg_out445 , sg_out446 , sg_out449 , sg_out450 , sg_out451 , sg_out452 , sg_out453 , sg_out454 , sg_out455 , sg_out456 , sg_out457 , sg_out458 , sg_out459 , sg_out460 , sg_out461 , sg_out462 , sg_out463 , sg_out464 , sg_out465 , sg_out466 , sg_out467 , sg_out468 , sg_out469 , sg_out470 , sg_out471 , sg_out472 , sg_out473 , sg_out474 , sg_out475 , sg_out476 , sg_out477 , sg_out478 , dig_t0 , dig_t1 , dig_t2 , dig_t3 , dig_t4 , dig_t5 , dig_t6 , dig_t7 , dig_t8 , dig_t9 , dig_t10 , dig_t11 , dig_t12 , dig_t13 , dig_t14 , dig_t15 , dig_t16 , dig_t17 , dig_t18 , dig_t19 , dig_t20 , dig_t21 , dig_t22 , dig_t23 , dig_t24 , dig_t25 , dig_t26 , dig_t27 , dig_t28 , dig_t29 , dig_t30 , dig_t31 , dig_t32 , dig_t33 , dig_t34 , dig_t35 , dig_t36 , dig_t37 , dig_t38 , dig_t39 , dig_t40 , dig_t41 , dig_t42 , dig_t43 , dig_t44 , dig_t45 , dig_t46 , dig_t47 , dig_t48 , dig_t49 , dig_t50 , dig_t51 , dig_t52 , dig_t53 , dig_t54 , dig_t55 , dig_t56 , dig_t57 , dig_t58 , dig_t59 , dig_t60 , dig_t61 , dig_t62 , dig_t63 , dig_t64 , dig_t65 , dig_t66 , dig_t67 , dig_t68 , dig_t69 , dig_t70 , dig_t71 , dig_t72 , dig_t73 , dig_t74 , dig_t75 , dig_t76 , dig_t77 , dig_t78 , dig_t79 , dig_t80 , dig_t81 , dig_t82 , dig_t83 , dig_t84 , dig_t85 , dig_t86 , dig_t87 , dig_t88 , dig_t89 , dig_t90 , dig_t91 , dig_t92 , dig_t93 , dig_t94 , dig_t95 , dig_t96 , dig_t97 , dig_t98 , dig_t99 , dig_t100 , dig_t101 , dig_t102 , dig_t103 , dig_t104 , dig_t105 , dig_t106 , dig_t107 , dig_t108 , dig_t109 , dig_t110 , dig_t111 , dig_t112 , dig_t113 , dig_t114 , dig_t115 , dig_t116 , dig_t117 , dig_t118 , dig_t119 , dig_t120 , dig_t121 , dig_t122 , dig_t123 , dig_t124 , dig_t125 , dig_t126 , dig_t127 , dig_t128 , dig_t129 , dig_t130 , dig_t131 , dig_t132 , dig_t133 , dig_t134 , dig_t135 , dig_t136 , dig_t137 , dig_t138 , dig_t139 , dig_t140 , dig_t141 , dig_t142 , dig_t143 , dig_t144 , dig_t145 , dig_t146 , dig_t147 , dig_t148 , dig_t149 , dig_t150 , dig_t151 , dig_t152 , dig_t153 , dig_t154 , dig_t155 , dig_t156 , dig_t157 , dig_t158 , dig_t159 , dig_t160 , dig_t161 , dig_t162 , dig_t163 , dig_t164 , dig_t165 , dig_t166 , dig_t167 , dig_t168 , dig_t169 , dig_t170 , dig_t171 , dig_t172 , dig_t173 , dig_t174 , dig_t175 , dig_t176 , dig_t177 , dig_t178 , dig_t179 , dig_t180 , dig_t181 , dig_t182 , dig_t183 , dig_t184 , dig_t185 , dig_t186 , dig_t187 , dig_t188 , dig_t189 , dig_t190 , dig_t191 , dig_t192 , dig_t193 , dig_t194 , dig_t195 , dig_t196 , dig_t197 , dig_t198 , dig_t199 , dig_t200 , dig_t201 , dig_t202 , dig_t203 , dig_t204 , dig_t205 , dig_t206 , dig_t207 , dig_t208 , dig_t209 , in_do , out_do , out_data );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input sig;
  wire sig;
  input [9:0] start;
  wire [9:0] start;
  input [9:0] goal;
  wire [9:0] goal;
  input dig_w;
  wire dig_w;
  input [9:0] data_in33;
  wire [9:0] data_in33;
  input [9:0] data_in34;
  wire [9:0] data_in34;
  input [9:0] data_in35;
  wire [9:0] data_in35;
  input [9:0] data_in36;
  wire [9:0] data_in36;
  input [9:0] data_in37;
  wire [9:0] data_in37;
  input [9:0] data_in38;
  wire [9:0] data_in38;
  input [9:0] data_in39;
  wire [9:0] data_in39;
  input [9:0] data_in40;
  wire [9:0] data_in40;
  input [9:0] data_in41;
  wire [9:0] data_in41;
  input [9:0] data_in42;
  wire [9:0] data_in42;
  input [9:0] data_in43;
  wire [9:0] data_in43;
  input [9:0] data_in44;
  wire [9:0] data_in44;
  input [9:0] data_in45;
  wire [9:0] data_in45;
  input [9:0] data_in46;
  wire [9:0] data_in46;
  input [9:0] data_in47;
  wire [9:0] data_in47;
  input [9:0] data_in48;
  wire [9:0] data_in48;
  input [9:0] data_in49;
  wire [9:0] data_in49;
  input [9:0] data_in50;
  wire [9:0] data_in50;
  input [9:0] data_in51;
  wire [9:0] data_in51;
  input [9:0] data_in52;
  wire [9:0] data_in52;
  input [9:0] data_in53;
  wire [9:0] data_in53;
  input [9:0] data_in54;
  wire [9:0] data_in54;
  input [9:0] data_in55;
  wire [9:0] data_in55;
  input [9:0] data_in56;
  wire [9:0] data_in56;
  input [9:0] data_in57;
  wire [9:0] data_in57;
  input [9:0] data_in58;
  wire [9:0] data_in58;
  input [9:0] data_in59;
  wire [9:0] data_in59;
  input [9:0] data_in60;
  wire [9:0] data_in60;
  input [9:0] data_in61;
  wire [9:0] data_in61;
  input [9:0] data_in62;
  wire [9:0] data_in62;
  input [9:0] data_in65;
  wire [9:0] data_in65;
  input [9:0] data_in66;
  wire [9:0] data_in66;
  input [9:0] data_in67;
  wire [9:0] data_in67;
  input [9:0] data_in68;
  wire [9:0] data_in68;
  input [9:0] data_in69;
  wire [9:0] data_in69;
  input [9:0] data_in70;
  wire [9:0] data_in70;
  input [9:0] data_in71;
  wire [9:0] data_in71;
  input [9:0] data_in72;
  wire [9:0] data_in72;
  input [9:0] data_in73;
  wire [9:0] data_in73;
  input [9:0] data_in74;
  wire [9:0] data_in74;
  input [9:0] data_in75;
  wire [9:0] data_in75;
  input [9:0] data_in76;
  wire [9:0] data_in76;
  input [9:0] data_in77;
  wire [9:0] data_in77;
  input [9:0] data_in78;
  wire [9:0] data_in78;
  input [9:0] data_in79;
  wire [9:0] data_in79;
  input [9:0] data_in80;
  wire [9:0] data_in80;
  input [9:0] data_in81;
  wire [9:0] data_in81;
  input [9:0] data_in82;
  wire [9:0] data_in82;
  input [9:0] data_in83;
  wire [9:0] data_in83;
  input [9:0] data_in84;
  wire [9:0] data_in84;
  input [9:0] data_in85;
  wire [9:0] data_in85;
  input [9:0] data_in86;
  wire [9:0] data_in86;
  input [9:0] data_in87;
  wire [9:0] data_in87;
  input [9:0] data_in88;
  wire [9:0] data_in88;
  input [9:0] data_in89;
  wire [9:0] data_in89;
  input [9:0] data_in90;
  wire [9:0] data_in90;
  input [9:0] data_in91;
  wire [9:0] data_in91;
  input [9:0] data_in92;
  wire [9:0] data_in92;
  input [9:0] data_in93;
  wire [9:0] data_in93;
  input [9:0] data_in94;
  wire [9:0] data_in94;
  input [9:0] data_in97;
  wire [9:0] data_in97;
  input [9:0] data_in98;
  wire [9:0] data_in98;
  input [9:0] data_in99;
  wire [9:0] data_in99;
  input [9:0] data_in100;
  wire [9:0] data_in100;
  input [9:0] data_in101;
  wire [9:0] data_in101;
  input [9:0] data_in102;
  wire [9:0] data_in102;
  input [9:0] data_in103;
  wire [9:0] data_in103;
  input [9:0] data_in104;
  wire [9:0] data_in104;
  input [9:0] data_in105;
  wire [9:0] data_in105;
  input [9:0] data_in106;
  wire [9:0] data_in106;
  input [9:0] data_in107;
  wire [9:0] data_in107;
  input [9:0] data_in108;
  wire [9:0] data_in108;
  input [9:0] data_in109;
  wire [9:0] data_in109;
  input [9:0] data_in110;
  wire [9:0] data_in110;
  input [9:0] data_in111;
  wire [9:0] data_in111;
  input [9:0] data_in112;
  wire [9:0] data_in112;
  input [9:0] data_in113;
  wire [9:0] data_in113;
  input [9:0] data_in114;
  wire [9:0] data_in114;
  input [9:0] data_in115;
  wire [9:0] data_in115;
  input [9:0] data_in116;
  wire [9:0] data_in116;
  input [9:0] data_in117;
  wire [9:0] data_in117;
  input [9:0] data_in118;
  wire [9:0] data_in118;
  input [9:0] data_in119;
  wire [9:0] data_in119;
  input [9:0] data_in120;
  wire [9:0] data_in120;
  input [9:0] data_in121;
  wire [9:0] data_in121;
  input [9:0] data_in122;
  wire [9:0] data_in122;
  input [9:0] data_in123;
  wire [9:0] data_in123;
  input [9:0] data_in124;
  wire [9:0] data_in124;
  input [9:0] data_in125;
  wire [9:0] data_in125;
  input [9:0] data_in126;
  wire [9:0] data_in126;
  input [9:0] data_in129;
  wire [9:0] data_in129;
  input [9:0] data_in130;
  wire [9:0] data_in130;
  input [9:0] data_in131;
  wire [9:0] data_in131;
  input [9:0] data_in132;
  wire [9:0] data_in132;
  input [9:0] data_in133;
  wire [9:0] data_in133;
  input [9:0] data_in134;
  wire [9:0] data_in134;
  input [9:0] data_in135;
  wire [9:0] data_in135;
  input [9:0] data_in136;
  wire [9:0] data_in136;
  input [9:0] data_in137;
  wire [9:0] data_in137;
  input [9:0] data_in138;
  wire [9:0] data_in138;
  input [9:0] data_in139;
  wire [9:0] data_in139;
  input [9:0] data_in140;
  wire [9:0] data_in140;
  input [9:0] data_in141;
  wire [9:0] data_in141;
  input [9:0] data_in142;
  wire [9:0] data_in142;
  input [9:0] data_in143;
  wire [9:0] data_in143;
  input [9:0] data_in144;
  wire [9:0] data_in144;
  input [9:0] data_in145;
  wire [9:0] data_in145;
  input [9:0] data_in146;
  wire [9:0] data_in146;
  input [9:0] data_in147;
  wire [9:0] data_in147;
  input [9:0] data_in148;
  wire [9:0] data_in148;
  input [9:0] data_in149;
  wire [9:0] data_in149;
  input [9:0] data_in150;
  wire [9:0] data_in150;
  input [9:0] data_in151;
  wire [9:0] data_in151;
  input [9:0] data_in152;
  wire [9:0] data_in152;
  input [9:0] data_in153;
  wire [9:0] data_in153;
  input [9:0] data_in154;
  wire [9:0] data_in154;
  input [9:0] data_in155;
  wire [9:0] data_in155;
  input [9:0] data_in156;
  wire [9:0] data_in156;
  input [9:0] data_in157;
  wire [9:0] data_in157;
  input [9:0] data_in158;
  wire [9:0] data_in158;
  input [9:0] data_in161;
  wire [9:0] data_in161;
  input [9:0] data_in162;
  wire [9:0] data_in162;
  input [9:0] data_in163;
  wire [9:0] data_in163;
  input [9:0] data_in164;
  wire [9:0] data_in164;
  input [9:0] data_in165;
  wire [9:0] data_in165;
  input [9:0] data_in166;
  wire [9:0] data_in166;
  input [9:0] data_in167;
  wire [9:0] data_in167;
  input [9:0] data_in168;
  wire [9:0] data_in168;
  input [9:0] data_in169;
  wire [9:0] data_in169;
  input [9:0] data_in170;
  wire [9:0] data_in170;
  input [9:0] data_in171;
  wire [9:0] data_in171;
  input [9:0] data_in172;
  wire [9:0] data_in172;
  input [9:0] data_in173;
  wire [9:0] data_in173;
  input [9:0] data_in174;
  wire [9:0] data_in174;
  input [9:0] data_in175;
  wire [9:0] data_in175;
  input [9:0] data_in176;
  wire [9:0] data_in176;
  input [9:0] data_in177;
  wire [9:0] data_in177;
  input [9:0] data_in178;
  wire [9:0] data_in178;
  input [9:0] data_in179;
  wire [9:0] data_in179;
  input [9:0] data_in180;
  wire [9:0] data_in180;
  input [9:0] data_in181;
  wire [9:0] data_in181;
  input [9:0] data_in182;
  wire [9:0] data_in182;
  input [9:0] data_in183;
  wire [9:0] data_in183;
  input [9:0] data_in184;
  wire [9:0] data_in184;
  input [9:0] data_in185;
  wire [9:0] data_in185;
  input [9:0] data_in186;
  wire [9:0] data_in186;
  input [9:0] data_in187;
  wire [9:0] data_in187;
  input [9:0] data_in188;
  wire [9:0] data_in188;
  input [9:0] data_in189;
  wire [9:0] data_in189;
  input [9:0] data_in190;
  wire [9:0] data_in190;
  input [9:0] data_in193;
  wire [9:0] data_in193;
  input [9:0] data_in194;
  wire [9:0] data_in194;
  input [9:0] data_in195;
  wire [9:0] data_in195;
  input [9:0] data_in196;
  wire [9:0] data_in196;
  input [9:0] data_in197;
  wire [9:0] data_in197;
  input [9:0] data_in198;
  wire [9:0] data_in198;
  input [9:0] data_in199;
  wire [9:0] data_in199;
  input [9:0] data_in200;
  wire [9:0] data_in200;
  input [9:0] data_in201;
  wire [9:0] data_in201;
  input [9:0] data_in202;
  wire [9:0] data_in202;
  input [9:0] data_in203;
  wire [9:0] data_in203;
  input [9:0] data_in204;
  wire [9:0] data_in204;
  input [9:0] data_in205;
  wire [9:0] data_in205;
  input [9:0] data_in206;
  wire [9:0] data_in206;
  input [9:0] data_in207;
  wire [9:0] data_in207;
  input [9:0] data_in208;
  wire [9:0] data_in208;
  input [9:0] data_in209;
  wire [9:0] data_in209;
  input [9:0] data_in210;
  wire [9:0] data_in210;
  input [9:0] data_in211;
  wire [9:0] data_in211;
  input [9:0] data_in212;
  wire [9:0] data_in212;
  input [9:0] data_in213;
  wire [9:0] data_in213;
  input [9:0] data_in214;
  wire [9:0] data_in214;
  input [9:0] data_in215;
  wire [9:0] data_in215;
  input [9:0] data_in216;
  wire [9:0] data_in216;
  input [9:0] data_in217;
  wire [9:0] data_in217;
  input [9:0] data_in218;
  wire [9:0] data_in218;
  input [9:0] data_in219;
  wire [9:0] data_in219;
  input [9:0] data_in220;
  wire [9:0] data_in220;
  input [9:0] data_in221;
  wire [9:0] data_in221;
  input [9:0] data_in222;
  wire [9:0] data_in222;
  input [9:0] data_in225;
  wire [9:0] data_in225;
  input [9:0] data_in226;
  wire [9:0] data_in226;
  input [9:0] data_in227;
  wire [9:0] data_in227;
  input [9:0] data_in228;
  wire [9:0] data_in228;
  input [9:0] data_in229;
  wire [9:0] data_in229;
  input [9:0] data_in230;
  wire [9:0] data_in230;
  input [9:0] data_in231;
  wire [9:0] data_in231;
  input [9:0] data_in232;
  wire [9:0] data_in232;
  input [9:0] data_in233;
  wire [9:0] data_in233;
  input [9:0] data_in234;
  wire [9:0] data_in234;
  input [9:0] data_in235;
  wire [9:0] data_in235;
  input [9:0] data_in236;
  wire [9:0] data_in236;
  input [9:0] data_in237;
  wire [9:0] data_in237;
  input [9:0] data_in238;
  wire [9:0] data_in238;
  input [9:0] data_in239;
  wire [9:0] data_in239;
  input [9:0] data_in240;
  wire [9:0] data_in240;
  input [9:0] data_in241;
  wire [9:0] data_in241;
  input [9:0] data_in242;
  wire [9:0] data_in242;
  input [9:0] data_in243;
  wire [9:0] data_in243;
  input [9:0] data_in244;
  wire [9:0] data_in244;
  input [9:0] data_in245;
  wire [9:0] data_in245;
  input [9:0] data_in246;
  wire [9:0] data_in246;
  input [9:0] data_in247;
  wire [9:0] data_in247;
  input [9:0] data_in248;
  wire [9:0] data_in248;
  input [9:0] data_in249;
  wire [9:0] data_in249;
  input [9:0] data_in250;
  wire [9:0] data_in250;
  input [9:0] data_in251;
  wire [9:0] data_in251;
  input [9:0] data_in252;
  wire [9:0] data_in252;
  input [9:0] data_in253;
  wire [9:0] data_in253;
  input [9:0] data_in254;
  wire [9:0] data_in254;
  input [9:0] data_in257;
  wire [9:0] data_in257;
  input [9:0] data_in258;
  wire [9:0] data_in258;
  input [9:0] data_in259;
  wire [9:0] data_in259;
  input [9:0] data_in260;
  wire [9:0] data_in260;
  input [9:0] data_in261;
  wire [9:0] data_in261;
  input [9:0] data_in262;
  wire [9:0] data_in262;
  input [9:0] data_in263;
  wire [9:0] data_in263;
  input [9:0] data_in264;
  wire [9:0] data_in264;
  input [9:0] data_in265;
  wire [9:0] data_in265;
  input [9:0] data_in266;
  wire [9:0] data_in266;
  input [9:0] data_in267;
  wire [9:0] data_in267;
  input [9:0] data_in268;
  wire [9:0] data_in268;
  input [9:0] data_in269;
  wire [9:0] data_in269;
  input [9:0] data_in270;
  wire [9:0] data_in270;
  input [9:0] data_in271;
  wire [9:0] data_in271;
  input [9:0] data_in272;
  wire [9:0] data_in272;
  input [9:0] data_in273;
  wire [9:0] data_in273;
  input [9:0] data_in274;
  wire [9:0] data_in274;
  input [9:0] data_in275;
  wire [9:0] data_in275;
  input [9:0] data_in276;
  wire [9:0] data_in276;
  input [9:0] data_in277;
  wire [9:0] data_in277;
  input [9:0] data_in278;
  wire [9:0] data_in278;
  input [9:0] data_in279;
  wire [9:0] data_in279;
  input [9:0] data_in280;
  wire [9:0] data_in280;
  input [9:0] data_in281;
  wire [9:0] data_in281;
  input [9:0] data_in282;
  wire [9:0] data_in282;
  input [9:0] data_in283;
  wire [9:0] data_in283;
  input [9:0] data_in284;
  wire [9:0] data_in284;
  input [9:0] data_in285;
  wire [9:0] data_in285;
  input [9:0] data_in286;
  wire [9:0] data_in286;
  input [9:0] data_in289;
  wire [9:0] data_in289;
  input [9:0] data_in290;
  wire [9:0] data_in290;
  input [9:0] data_in291;
  wire [9:0] data_in291;
  input [9:0] data_in292;
  wire [9:0] data_in292;
  input [9:0] data_in293;
  wire [9:0] data_in293;
  input [9:0] data_in294;
  wire [9:0] data_in294;
  input [9:0] data_in295;
  wire [9:0] data_in295;
  input [9:0] data_in296;
  wire [9:0] data_in296;
  input [9:0] data_in297;
  wire [9:0] data_in297;
  input [9:0] data_in298;
  wire [9:0] data_in298;
  input [9:0] data_in299;
  wire [9:0] data_in299;
  input [9:0] data_in300;
  wire [9:0] data_in300;
  input [9:0] data_in301;
  wire [9:0] data_in301;
  input [9:0] data_in302;
  wire [9:0] data_in302;
  input [9:0] data_in303;
  wire [9:0] data_in303;
  input [9:0] data_in304;
  wire [9:0] data_in304;
  input [9:0] data_in305;
  wire [9:0] data_in305;
  input [9:0] data_in306;
  wire [9:0] data_in306;
  input [9:0] data_in307;
  wire [9:0] data_in307;
  input [9:0] data_in308;
  wire [9:0] data_in308;
  input [9:0] data_in309;
  wire [9:0] data_in309;
  input [9:0] data_in310;
  wire [9:0] data_in310;
  input [9:0] data_in311;
  wire [9:0] data_in311;
  input [9:0] data_in312;
  wire [9:0] data_in312;
  input [9:0] data_in313;
  wire [9:0] data_in313;
  input [9:0] data_in314;
  wire [9:0] data_in314;
  input [9:0] data_in315;
  wire [9:0] data_in315;
  input [9:0] data_in316;
  wire [9:0] data_in316;
  input [9:0] data_in317;
  wire [9:0] data_in317;
  input [9:0] data_in318;
  wire [9:0] data_in318;
  input [9:0] data_in321;
  wire [9:0] data_in321;
  input [9:0] data_in322;
  wire [9:0] data_in322;
  input [9:0] data_in323;
  wire [9:0] data_in323;
  input [9:0] data_in324;
  wire [9:0] data_in324;
  input [9:0] data_in325;
  wire [9:0] data_in325;
  input [9:0] data_in326;
  wire [9:0] data_in326;
  input [9:0] data_in327;
  wire [9:0] data_in327;
  input [9:0] data_in328;
  wire [9:0] data_in328;
  input [9:0] data_in329;
  wire [9:0] data_in329;
  input [9:0] data_in330;
  wire [9:0] data_in330;
  input [9:0] data_in331;
  wire [9:0] data_in331;
  input [9:0] data_in332;
  wire [9:0] data_in332;
  input [9:0] data_in333;
  wire [9:0] data_in333;
  input [9:0] data_in334;
  wire [9:0] data_in334;
  input [9:0] data_in335;
  wire [9:0] data_in335;
  input [9:0] data_in336;
  wire [9:0] data_in336;
  input [9:0] data_in337;
  wire [9:0] data_in337;
  input [9:0] data_in338;
  wire [9:0] data_in338;
  input [9:0] data_in339;
  wire [9:0] data_in339;
  input [9:0] data_in340;
  wire [9:0] data_in340;
  input [9:0] data_in341;
  wire [9:0] data_in341;
  input [9:0] data_in342;
  wire [9:0] data_in342;
  input [9:0] data_in343;
  wire [9:0] data_in343;
  input [9:0] data_in344;
  wire [9:0] data_in344;
  input [9:0] data_in345;
  wire [9:0] data_in345;
  input [9:0] data_in346;
  wire [9:0] data_in346;
  input [9:0] data_in347;
  wire [9:0] data_in347;
  input [9:0] data_in348;
  wire [9:0] data_in348;
  input [9:0] data_in349;
  wire [9:0] data_in349;
  input [9:0] data_in350;
  wire [9:0] data_in350;
  input [9:0] data_in353;
  wire [9:0] data_in353;
  input [9:0] data_in354;
  wire [9:0] data_in354;
  input [9:0] data_in355;
  wire [9:0] data_in355;
  input [9:0] data_in356;
  wire [9:0] data_in356;
  input [9:0] data_in357;
  wire [9:0] data_in357;
  input [9:0] data_in358;
  wire [9:0] data_in358;
  input [9:0] data_in359;
  wire [9:0] data_in359;
  input [9:0] data_in360;
  wire [9:0] data_in360;
  input [9:0] data_in361;
  wire [9:0] data_in361;
  input [9:0] data_in362;
  wire [9:0] data_in362;
  input [9:0] data_in363;
  wire [9:0] data_in363;
  input [9:0] data_in364;
  wire [9:0] data_in364;
  input [9:0] data_in365;
  wire [9:0] data_in365;
  input [9:0] data_in366;
  wire [9:0] data_in366;
  input [9:0] data_in367;
  wire [9:0] data_in367;
  input [9:0] data_in368;
  wire [9:0] data_in368;
  input [9:0] data_in369;
  wire [9:0] data_in369;
  input [9:0] data_in370;
  wire [9:0] data_in370;
  input [9:0] data_in371;
  wire [9:0] data_in371;
  input [9:0] data_in372;
  wire [9:0] data_in372;
  input [9:0] data_in373;
  wire [9:0] data_in373;
  input [9:0] data_in374;
  wire [9:0] data_in374;
  input [9:0] data_in375;
  wire [9:0] data_in375;
  input [9:0] data_in376;
  wire [9:0] data_in376;
  input [9:0] data_in377;
  wire [9:0] data_in377;
  input [9:0] data_in378;
  wire [9:0] data_in378;
  input [9:0] data_in379;
  wire [9:0] data_in379;
  input [9:0] data_in380;
  wire [9:0] data_in380;
  input [9:0] data_in381;
  wire [9:0] data_in381;
  input [9:0] data_in382;
  wire [9:0] data_in382;
  input [9:0] data_in385;
  wire [9:0] data_in385;
  input [9:0] data_in386;
  wire [9:0] data_in386;
  input [9:0] data_in387;
  wire [9:0] data_in387;
  input [9:0] data_in388;
  wire [9:0] data_in388;
  input [9:0] data_in389;
  wire [9:0] data_in389;
  input [9:0] data_in390;
  wire [9:0] data_in390;
  input [9:0] data_in391;
  wire [9:0] data_in391;
  input [9:0] data_in392;
  wire [9:0] data_in392;
  input [9:0] data_in393;
  wire [9:0] data_in393;
  input [9:0] data_in394;
  wire [9:0] data_in394;
  input [9:0] data_in395;
  wire [9:0] data_in395;
  input [9:0] data_in396;
  wire [9:0] data_in396;
  input [9:0] data_in397;
  wire [9:0] data_in397;
  input [9:0] data_in398;
  wire [9:0] data_in398;
  input [9:0] data_in399;
  wire [9:0] data_in399;
  input [9:0] data_in400;
  wire [9:0] data_in400;
  input [9:0] data_in401;
  wire [9:0] data_in401;
  input [9:0] data_in402;
  wire [9:0] data_in402;
  input [9:0] data_in403;
  wire [9:0] data_in403;
  input [9:0] data_in404;
  wire [9:0] data_in404;
  input [9:0] data_in405;
  wire [9:0] data_in405;
  input [9:0] data_in406;
  wire [9:0] data_in406;
  input [9:0] data_in407;
  wire [9:0] data_in407;
  input [9:0] data_in408;
  wire [9:0] data_in408;
  input [9:0] data_in409;
  wire [9:0] data_in409;
  input [9:0] data_in410;
  wire [9:0] data_in410;
  input [9:0] data_in411;
  wire [9:0] data_in411;
  input [9:0] data_in412;
  wire [9:0] data_in412;
  input [9:0] data_in413;
  wire [9:0] data_in413;
  input [9:0] data_in414;
  wire [9:0] data_in414;
  input [9:0] data_in417;
  wire [9:0] data_in417;
  input [9:0] data_in418;
  wire [9:0] data_in418;
  input [9:0] data_in419;
  wire [9:0] data_in419;
  input [9:0] data_in420;
  wire [9:0] data_in420;
  input [9:0] data_in421;
  wire [9:0] data_in421;
  input [9:0] data_in422;
  wire [9:0] data_in422;
  input [9:0] data_in423;
  wire [9:0] data_in423;
  input [9:0] data_in424;
  wire [9:0] data_in424;
  input [9:0] data_in425;
  wire [9:0] data_in425;
  input [9:0] data_in426;
  wire [9:0] data_in426;
  input [9:0] data_in427;
  wire [9:0] data_in427;
  input [9:0] data_in428;
  wire [9:0] data_in428;
  input [9:0] data_in429;
  wire [9:0] data_in429;
  input [9:0] data_in430;
  wire [9:0] data_in430;
  input [9:0] data_in431;
  wire [9:0] data_in431;
  input [9:0] data_in432;
  wire [9:0] data_in432;
  input [9:0] data_in433;
  wire [9:0] data_in433;
  input [9:0] data_in434;
  wire [9:0] data_in434;
  input [9:0] data_in435;
  wire [9:0] data_in435;
  input [9:0] data_in436;
  wire [9:0] data_in436;
  input [9:0] data_in437;
  wire [9:0] data_in437;
  input [9:0] data_in438;
  wire [9:0] data_in438;
  input [9:0] data_in439;
  wire [9:0] data_in439;
  input [9:0] data_in440;
  wire [9:0] data_in440;
  input [9:0] data_in441;
  wire [9:0] data_in441;
  input [9:0] data_in442;
  wire [9:0] data_in442;
  input [9:0] data_in443;
  wire [9:0] data_in443;
  input [9:0] data_in444;
  wire [9:0] data_in444;
  input [9:0] data_in445;
  wire [9:0] data_in445;
  input [9:0] data_in446;
  wire [9:0] data_in446;
  input [9:0] data_in449;
  wire [9:0] data_in449;
  input [9:0] data_in450;
  wire [9:0] data_in450;
  input [9:0] data_in451;
  wire [9:0] data_in451;
  input [9:0] data_in452;
  wire [9:0] data_in452;
  input [9:0] data_in453;
  wire [9:0] data_in453;
  input [9:0] data_in454;
  wire [9:0] data_in454;
  input [9:0] data_in455;
  wire [9:0] data_in455;
  input [9:0] data_in456;
  wire [9:0] data_in456;
  input [9:0] data_in457;
  wire [9:0] data_in457;
  input [9:0] data_in458;
  wire [9:0] data_in458;
  input [9:0] data_in459;
  wire [9:0] data_in459;
  input [9:0] data_in460;
  wire [9:0] data_in460;
  input [9:0] data_in461;
  wire [9:0] data_in461;
  input [9:0] data_in462;
  wire [9:0] data_in462;
  input [9:0] data_in463;
  wire [9:0] data_in463;
  input [9:0] data_in464;
  wire [9:0] data_in464;
  input [9:0] data_in465;
  wire [9:0] data_in465;
  input [9:0] data_in466;
  wire [9:0] data_in466;
  input [9:0] data_in467;
  wire [9:0] data_in467;
  input [9:0] data_in468;
  wire [9:0] data_in468;
  input [9:0] data_in469;
  wire [9:0] data_in469;
  input [9:0] data_in470;
  wire [9:0] data_in470;
  input [9:0] data_in471;
  wire [9:0] data_in471;
  input [9:0] data_in472;
  wire [9:0] data_in472;
  input [9:0] data_in473;
  wire [9:0] data_in473;
  input [9:0] data_in474;
  wire [9:0] data_in474;
  input [9:0] data_in475;
  wire [9:0] data_in475;
  input [9:0] data_in476;
  wire [9:0] data_in476;
  input [9:0] data_in477;
  wire [9:0] data_in477;
  input [9:0] data_in478;
  wire [9:0] data_in478;
  output [9:0] data_out_org33;
  wire [9:0] data_out_org33;
  output [9:0] data_out_org34;
  wire [9:0] data_out_org34;
  output [9:0] data_out_org35;
  wire [9:0] data_out_org35;
  output [9:0] data_out_org36;
  wire [9:0] data_out_org36;
  output [9:0] data_out_org37;
  wire [9:0] data_out_org37;
  output [9:0] data_out_org38;
  wire [9:0] data_out_org38;
  output [9:0] data_out_org39;
  wire [9:0] data_out_org39;
  output [9:0] data_out_org40;
  wire [9:0] data_out_org40;
  output [9:0] data_out_org41;
  wire [9:0] data_out_org41;
  output [9:0] data_out_org42;
  wire [9:0] data_out_org42;
  output [9:0] data_out_org43;
  wire [9:0] data_out_org43;
  output [9:0] data_out_org44;
  wire [9:0] data_out_org44;
  output [9:0] data_out_org45;
  wire [9:0] data_out_org45;
  output [9:0] data_out_org46;
  wire [9:0] data_out_org46;
  output [9:0] data_out_org47;
  wire [9:0] data_out_org47;
  output [9:0] data_out_org48;
  wire [9:0] data_out_org48;
  output [9:0] data_out_org49;
  wire [9:0] data_out_org49;
  output [9:0] data_out_org50;
  wire [9:0] data_out_org50;
  output [9:0] data_out_org51;
  wire [9:0] data_out_org51;
  output [9:0] data_out_org52;
  wire [9:0] data_out_org52;
  output [9:0] data_out_org53;
  wire [9:0] data_out_org53;
  output [9:0] data_out_org54;
  wire [9:0] data_out_org54;
  output [9:0] data_out_org55;
  wire [9:0] data_out_org55;
  output [9:0] data_out_org56;
  wire [9:0] data_out_org56;
  output [9:0] data_out_org57;
  wire [9:0] data_out_org57;
  output [9:0] data_out_org58;
  wire [9:0] data_out_org58;
  output [9:0] data_out_org59;
  wire [9:0] data_out_org59;
  output [9:0] data_out_org60;
  wire [9:0] data_out_org60;
  output [9:0] data_out_org61;
  wire [9:0] data_out_org61;
  output [9:0] data_out_org62;
  wire [9:0] data_out_org62;
  output [9:0] data_out_org65;
  wire [9:0] data_out_org65;
  output [9:0] data_out_org66;
  wire [9:0] data_out_org66;
  output [9:0] data_out_org67;
  wire [9:0] data_out_org67;
  output [9:0] data_out_org68;
  wire [9:0] data_out_org68;
  output [9:0] data_out_org69;
  wire [9:0] data_out_org69;
  output [9:0] data_out_org70;
  wire [9:0] data_out_org70;
  output [9:0] data_out_org71;
  wire [9:0] data_out_org71;
  output [9:0] data_out_org72;
  wire [9:0] data_out_org72;
  output [9:0] data_out_org73;
  wire [9:0] data_out_org73;
  output [9:0] data_out_org74;
  wire [9:0] data_out_org74;
  output [9:0] data_out_org75;
  wire [9:0] data_out_org75;
  output [9:0] data_out_org76;
  wire [9:0] data_out_org76;
  output [9:0] data_out_org77;
  wire [9:0] data_out_org77;
  output [9:0] data_out_org78;
  wire [9:0] data_out_org78;
  output [9:0] data_out_org79;
  wire [9:0] data_out_org79;
  output [9:0] data_out_org80;
  wire [9:0] data_out_org80;
  output [9:0] data_out_org81;
  wire [9:0] data_out_org81;
  output [9:0] data_out_org82;
  wire [9:0] data_out_org82;
  output [9:0] data_out_org83;
  wire [9:0] data_out_org83;
  output [9:0] data_out_org84;
  wire [9:0] data_out_org84;
  output [9:0] data_out_org85;
  wire [9:0] data_out_org85;
  output [9:0] data_out_org86;
  wire [9:0] data_out_org86;
  output [9:0] data_out_org87;
  wire [9:0] data_out_org87;
  output [9:0] data_out_org88;
  wire [9:0] data_out_org88;
  output [9:0] data_out_org89;
  wire [9:0] data_out_org89;
  output [9:0] data_out_org90;
  wire [9:0] data_out_org90;
  output [9:0] data_out_org91;
  wire [9:0] data_out_org91;
  output [9:0] data_out_org92;
  wire [9:0] data_out_org92;
  output [9:0] data_out_org93;
  wire [9:0] data_out_org93;
  output [9:0] data_out_org94;
  wire [9:0] data_out_org94;
  output [9:0] data_out_org97;
  wire [9:0] data_out_org97;
  output [9:0] data_out_org98;
  wire [9:0] data_out_org98;
  output [9:0] data_out_org99;
  wire [9:0] data_out_org99;
  output [9:0] data_out_org100;
  wire [9:0] data_out_org100;
  output [9:0] data_out_org101;
  wire [9:0] data_out_org101;
  output [9:0] data_out_org102;
  wire [9:0] data_out_org102;
  output [9:0] data_out_org103;
  wire [9:0] data_out_org103;
  output [9:0] data_out_org104;
  wire [9:0] data_out_org104;
  output [9:0] data_out_org105;
  wire [9:0] data_out_org105;
  output [9:0] data_out_org106;
  wire [9:0] data_out_org106;
  output [9:0] data_out_org107;
  wire [9:0] data_out_org107;
  output [9:0] data_out_org108;
  wire [9:0] data_out_org108;
  output [9:0] data_out_org109;
  wire [9:0] data_out_org109;
  output [9:0] data_out_org110;
  wire [9:0] data_out_org110;
  output [9:0] data_out_org111;
  wire [9:0] data_out_org111;
  output [9:0] data_out_org112;
  wire [9:0] data_out_org112;
  output [9:0] data_out_org113;
  wire [9:0] data_out_org113;
  output [9:0] data_out_org114;
  wire [9:0] data_out_org114;
  output [9:0] data_out_org115;
  wire [9:0] data_out_org115;
  output [9:0] data_out_org116;
  wire [9:0] data_out_org116;
  output [9:0] data_out_org117;
  wire [9:0] data_out_org117;
  output [9:0] data_out_org118;
  wire [9:0] data_out_org118;
  output [9:0] data_out_org119;
  wire [9:0] data_out_org119;
  output [9:0] data_out_org120;
  wire [9:0] data_out_org120;
  output [9:0] data_out_org121;
  wire [9:0] data_out_org121;
  output [9:0] data_out_org122;
  wire [9:0] data_out_org122;
  output [9:0] data_out_org123;
  wire [9:0] data_out_org123;
  output [9:0] data_out_org124;
  wire [9:0] data_out_org124;
  output [9:0] data_out_org125;
  wire [9:0] data_out_org125;
  output [9:0] data_out_org126;
  wire [9:0] data_out_org126;
  output [9:0] data_out_org129;
  wire [9:0] data_out_org129;
  output [9:0] data_out_org130;
  wire [9:0] data_out_org130;
  output [9:0] data_out_org131;
  wire [9:0] data_out_org131;
  output [9:0] data_out_org132;
  wire [9:0] data_out_org132;
  output [9:0] data_out_org133;
  wire [9:0] data_out_org133;
  output [9:0] data_out_org134;
  wire [9:0] data_out_org134;
  output [9:0] data_out_org135;
  wire [9:0] data_out_org135;
  output [9:0] data_out_org136;
  wire [9:0] data_out_org136;
  output [9:0] data_out_org137;
  wire [9:0] data_out_org137;
  output [9:0] data_out_org138;
  wire [9:0] data_out_org138;
  output [9:0] data_out_org139;
  wire [9:0] data_out_org139;
  output [9:0] data_out_org140;
  wire [9:0] data_out_org140;
  output [9:0] data_out_org141;
  wire [9:0] data_out_org141;
  output [9:0] data_out_org142;
  wire [9:0] data_out_org142;
  output [9:0] data_out_org143;
  wire [9:0] data_out_org143;
  output [9:0] data_out_org144;
  wire [9:0] data_out_org144;
  output [9:0] data_out_org145;
  wire [9:0] data_out_org145;
  output [9:0] data_out_org146;
  wire [9:0] data_out_org146;
  output [9:0] data_out_org147;
  wire [9:0] data_out_org147;
  output [9:0] data_out_org148;
  wire [9:0] data_out_org148;
  output [9:0] data_out_org149;
  wire [9:0] data_out_org149;
  output [9:0] data_out_org150;
  wire [9:0] data_out_org150;
  output [9:0] data_out_org151;
  wire [9:0] data_out_org151;
  output [9:0] data_out_org152;
  wire [9:0] data_out_org152;
  output [9:0] data_out_org153;
  wire [9:0] data_out_org153;
  output [9:0] data_out_org154;
  wire [9:0] data_out_org154;
  output [9:0] data_out_org155;
  wire [9:0] data_out_org155;
  output [9:0] data_out_org156;
  wire [9:0] data_out_org156;
  output [9:0] data_out_org157;
  wire [9:0] data_out_org157;
  output [9:0] data_out_org158;
  wire [9:0] data_out_org158;
  output [9:0] data_out_org161;
  wire [9:0] data_out_org161;
  output [9:0] data_out_org162;
  wire [9:0] data_out_org162;
  output [9:0] data_out_org163;
  wire [9:0] data_out_org163;
  output [9:0] data_out_org164;
  wire [9:0] data_out_org164;
  output [9:0] data_out_org165;
  wire [9:0] data_out_org165;
  output [9:0] data_out_org166;
  wire [9:0] data_out_org166;
  output [9:0] data_out_org167;
  wire [9:0] data_out_org167;
  output [9:0] data_out_org168;
  wire [9:0] data_out_org168;
  output [9:0] data_out_org169;
  wire [9:0] data_out_org169;
  output [9:0] data_out_org170;
  wire [9:0] data_out_org170;
  output [9:0] data_out_org171;
  wire [9:0] data_out_org171;
  output [9:0] data_out_org172;
  wire [9:0] data_out_org172;
  output [9:0] data_out_org173;
  wire [9:0] data_out_org173;
  output [9:0] data_out_org174;
  wire [9:0] data_out_org174;
  output [9:0] data_out_org175;
  wire [9:0] data_out_org175;
  output [9:0] data_out_org176;
  wire [9:0] data_out_org176;
  output [9:0] data_out_org177;
  wire [9:0] data_out_org177;
  output [9:0] data_out_org178;
  wire [9:0] data_out_org178;
  output [9:0] data_out_org179;
  wire [9:0] data_out_org179;
  output [9:0] data_out_org180;
  wire [9:0] data_out_org180;
  output [9:0] data_out_org181;
  wire [9:0] data_out_org181;
  output [9:0] data_out_org182;
  wire [9:0] data_out_org182;
  output [9:0] data_out_org183;
  wire [9:0] data_out_org183;
  output [9:0] data_out_org184;
  wire [9:0] data_out_org184;
  output [9:0] data_out_org185;
  wire [9:0] data_out_org185;
  output [9:0] data_out_org186;
  wire [9:0] data_out_org186;
  output [9:0] data_out_org187;
  wire [9:0] data_out_org187;
  output [9:0] data_out_org188;
  wire [9:0] data_out_org188;
  output [9:0] data_out_org189;
  wire [9:0] data_out_org189;
  output [9:0] data_out_org190;
  wire [9:0] data_out_org190;
  output [9:0] data_out_org193;
  wire [9:0] data_out_org193;
  output [9:0] data_out_org194;
  wire [9:0] data_out_org194;
  output [9:0] data_out_org195;
  wire [9:0] data_out_org195;
  output [9:0] data_out_org196;
  wire [9:0] data_out_org196;
  output [9:0] data_out_org197;
  wire [9:0] data_out_org197;
  output [9:0] data_out_org198;
  wire [9:0] data_out_org198;
  output [9:0] data_out_org199;
  wire [9:0] data_out_org199;
  output [9:0] data_out_org200;
  wire [9:0] data_out_org200;
  output [9:0] data_out_org201;
  wire [9:0] data_out_org201;
  output [9:0] data_out_org202;
  wire [9:0] data_out_org202;
  output [9:0] data_out_org203;
  wire [9:0] data_out_org203;
  output [9:0] data_out_org204;
  wire [9:0] data_out_org204;
  output [9:0] data_out_org205;
  wire [9:0] data_out_org205;
  output [9:0] data_out_org206;
  wire [9:0] data_out_org206;
  output [9:0] data_out_org207;
  wire [9:0] data_out_org207;
  output [9:0] data_out_org208;
  wire [9:0] data_out_org208;
  output [9:0] data_out_org209;
  wire [9:0] data_out_org209;
  output [9:0] data_out_org210;
  wire [9:0] data_out_org210;
  output [9:0] data_out_org211;
  wire [9:0] data_out_org211;
  output [9:0] data_out_org212;
  wire [9:0] data_out_org212;
  output [9:0] data_out_org213;
  wire [9:0] data_out_org213;
  output [9:0] data_out_org214;
  wire [9:0] data_out_org214;
  output [9:0] data_out_org215;
  wire [9:0] data_out_org215;
  output [9:0] data_out_org216;
  wire [9:0] data_out_org216;
  output [9:0] data_out_org217;
  wire [9:0] data_out_org217;
  output [9:0] data_out_org218;
  wire [9:0] data_out_org218;
  output [9:0] data_out_org219;
  wire [9:0] data_out_org219;
  output [9:0] data_out_org220;
  wire [9:0] data_out_org220;
  output [9:0] data_out_org221;
  wire [9:0] data_out_org221;
  output [9:0] data_out_org222;
  wire [9:0] data_out_org222;
  output [9:0] data_out_org225;
  wire [9:0] data_out_org225;
  output [9:0] data_out_org226;
  wire [9:0] data_out_org226;
  output [9:0] data_out_org227;
  wire [9:0] data_out_org227;
  output [9:0] data_out_org228;
  wire [9:0] data_out_org228;
  output [9:0] data_out_org229;
  wire [9:0] data_out_org229;
  output [9:0] data_out_org230;
  wire [9:0] data_out_org230;
  output [9:0] data_out_org231;
  wire [9:0] data_out_org231;
  output [9:0] data_out_org232;
  wire [9:0] data_out_org232;
  output [9:0] data_out_org233;
  wire [9:0] data_out_org233;
  output [9:0] data_out_org234;
  wire [9:0] data_out_org234;
  output [9:0] data_out_org235;
  wire [9:0] data_out_org235;
  output [9:0] data_out_org236;
  wire [9:0] data_out_org236;
  output [9:0] data_out_org237;
  wire [9:0] data_out_org237;
  output [9:0] data_out_org238;
  wire [9:0] data_out_org238;
  output [9:0] data_out_org239;
  wire [9:0] data_out_org239;
  output [9:0] data_out_org240;
  wire [9:0] data_out_org240;
  output [9:0] data_out_org241;
  wire [9:0] data_out_org241;
  output [9:0] data_out_org242;
  wire [9:0] data_out_org242;
  output [9:0] data_out_org243;
  wire [9:0] data_out_org243;
  output [9:0] data_out_org244;
  wire [9:0] data_out_org244;
  output [9:0] data_out_org245;
  wire [9:0] data_out_org245;
  output [9:0] data_out_org246;
  wire [9:0] data_out_org246;
  output [9:0] data_out_org247;
  wire [9:0] data_out_org247;
  output [9:0] data_out_org248;
  wire [9:0] data_out_org248;
  output [9:0] data_out_org249;
  wire [9:0] data_out_org249;
  output [9:0] data_out_org250;
  wire [9:0] data_out_org250;
  output [9:0] data_out_org251;
  wire [9:0] data_out_org251;
  output [9:0] data_out_org252;
  wire [9:0] data_out_org252;
  output [9:0] data_out_org253;
  wire [9:0] data_out_org253;
  output [9:0] data_out_org254;
  wire [9:0] data_out_org254;
  output [9:0] data_out_org257;
  wire [9:0] data_out_org257;
  output [9:0] data_out_org258;
  wire [9:0] data_out_org258;
  output [9:0] data_out_org259;
  wire [9:0] data_out_org259;
  output [9:0] data_out_org260;
  wire [9:0] data_out_org260;
  output [9:0] data_out_org261;
  wire [9:0] data_out_org261;
  output [9:0] data_out_org262;
  wire [9:0] data_out_org262;
  output [9:0] data_out_org263;
  wire [9:0] data_out_org263;
  output [9:0] data_out_org264;
  wire [9:0] data_out_org264;
  output [9:0] data_out_org265;
  wire [9:0] data_out_org265;
  output [9:0] data_out_org266;
  wire [9:0] data_out_org266;
  output [9:0] data_out_org267;
  wire [9:0] data_out_org267;
  output [9:0] data_out_org268;
  wire [9:0] data_out_org268;
  output [9:0] data_out_org269;
  wire [9:0] data_out_org269;
  output [9:0] data_out_org270;
  wire [9:0] data_out_org270;
  output [9:0] data_out_org271;
  wire [9:0] data_out_org271;
  output [9:0] data_out_org272;
  wire [9:0] data_out_org272;
  output [9:0] data_out_org273;
  wire [9:0] data_out_org273;
  output [9:0] data_out_org274;
  wire [9:0] data_out_org274;
  output [9:0] data_out_org275;
  wire [9:0] data_out_org275;
  output [9:0] data_out_org276;
  wire [9:0] data_out_org276;
  output [9:0] data_out_org277;
  wire [9:0] data_out_org277;
  output [9:0] data_out_org278;
  wire [9:0] data_out_org278;
  output [9:0] data_out_org279;
  wire [9:0] data_out_org279;
  output [9:0] data_out_org280;
  wire [9:0] data_out_org280;
  output [9:0] data_out_org281;
  wire [9:0] data_out_org281;
  output [9:0] data_out_org282;
  wire [9:0] data_out_org282;
  output [9:0] data_out_org283;
  wire [9:0] data_out_org283;
  output [9:0] data_out_org284;
  wire [9:0] data_out_org284;
  output [9:0] data_out_org285;
  wire [9:0] data_out_org285;
  output [9:0] data_out_org286;
  wire [9:0] data_out_org286;
  output [9:0] data_out_org289;
  wire [9:0] data_out_org289;
  output [9:0] data_out_org290;
  wire [9:0] data_out_org290;
  output [9:0] data_out_org291;
  wire [9:0] data_out_org291;
  output [9:0] data_out_org292;
  wire [9:0] data_out_org292;
  output [9:0] data_out_org293;
  wire [9:0] data_out_org293;
  output [9:0] data_out_org294;
  wire [9:0] data_out_org294;
  output [9:0] data_out_org295;
  wire [9:0] data_out_org295;
  output [9:0] data_out_org296;
  wire [9:0] data_out_org296;
  output [9:0] data_out_org297;
  wire [9:0] data_out_org297;
  output [9:0] data_out_org298;
  wire [9:0] data_out_org298;
  output [9:0] data_out_org299;
  wire [9:0] data_out_org299;
  output [9:0] data_out_org300;
  wire [9:0] data_out_org300;
  output [9:0] data_out_org301;
  wire [9:0] data_out_org301;
  output [9:0] data_out_org302;
  wire [9:0] data_out_org302;
  output [9:0] data_out_org303;
  wire [9:0] data_out_org303;
  output [9:0] data_out_org304;
  wire [9:0] data_out_org304;
  output [9:0] data_out_org305;
  wire [9:0] data_out_org305;
  output [9:0] data_out_org306;
  wire [9:0] data_out_org306;
  output [9:0] data_out_org307;
  wire [9:0] data_out_org307;
  output [9:0] data_out_org308;
  wire [9:0] data_out_org308;
  output [9:0] data_out_org309;
  wire [9:0] data_out_org309;
  output [9:0] data_out_org310;
  wire [9:0] data_out_org310;
  output [9:0] data_out_org311;
  wire [9:0] data_out_org311;
  output [9:0] data_out_org312;
  wire [9:0] data_out_org312;
  output [9:0] data_out_org313;
  wire [9:0] data_out_org313;
  output [9:0] data_out_org314;
  wire [9:0] data_out_org314;
  output [9:0] data_out_org315;
  wire [9:0] data_out_org315;
  output [9:0] data_out_org316;
  wire [9:0] data_out_org316;
  output [9:0] data_out_org317;
  wire [9:0] data_out_org317;
  output [9:0] data_out_org318;
  wire [9:0] data_out_org318;
  output [9:0] data_out_org321;
  wire [9:0] data_out_org321;
  output [9:0] data_out_org322;
  wire [9:0] data_out_org322;
  output [9:0] data_out_org323;
  wire [9:0] data_out_org323;
  output [9:0] data_out_org324;
  wire [9:0] data_out_org324;
  output [9:0] data_out_org325;
  wire [9:0] data_out_org325;
  output [9:0] data_out_org326;
  wire [9:0] data_out_org326;
  output [9:0] data_out_org327;
  wire [9:0] data_out_org327;
  output [9:0] data_out_org328;
  wire [9:0] data_out_org328;
  output [9:0] data_out_org329;
  wire [9:0] data_out_org329;
  output [9:0] data_out_org330;
  wire [9:0] data_out_org330;
  output [9:0] data_out_org331;
  wire [9:0] data_out_org331;
  output [9:0] data_out_org332;
  wire [9:0] data_out_org332;
  output [9:0] data_out_org333;
  wire [9:0] data_out_org333;
  output [9:0] data_out_org334;
  wire [9:0] data_out_org334;
  output [9:0] data_out_org335;
  wire [9:0] data_out_org335;
  output [9:0] data_out_org336;
  wire [9:0] data_out_org336;
  output [9:0] data_out_org337;
  wire [9:0] data_out_org337;
  output [9:0] data_out_org338;
  wire [9:0] data_out_org338;
  output [9:0] data_out_org339;
  wire [9:0] data_out_org339;
  output [9:0] data_out_org340;
  wire [9:0] data_out_org340;
  output [9:0] data_out_org341;
  wire [9:0] data_out_org341;
  output [9:0] data_out_org342;
  wire [9:0] data_out_org342;
  output [9:0] data_out_org343;
  wire [9:0] data_out_org343;
  output [9:0] data_out_org344;
  wire [9:0] data_out_org344;
  output [9:0] data_out_org345;
  wire [9:0] data_out_org345;
  output [9:0] data_out_org346;
  wire [9:0] data_out_org346;
  output [9:0] data_out_org347;
  wire [9:0] data_out_org347;
  output [9:0] data_out_org348;
  wire [9:0] data_out_org348;
  output [9:0] data_out_org349;
  wire [9:0] data_out_org349;
  output [9:0] data_out_org350;
  wire [9:0] data_out_org350;
  output [9:0] data_out_org353;
  wire [9:0] data_out_org353;
  output [9:0] data_out_org354;
  wire [9:0] data_out_org354;
  output [9:0] data_out_org355;
  wire [9:0] data_out_org355;
  output [9:0] data_out_org356;
  wire [9:0] data_out_org356;
  output [9:0] data_out_org357;
  wire [9:0] data_out_org357;
  output [9:0] data_out_org358;
  wire [9:0] data_out_org358;
  output [9:0] data_out_org359;
  wire [9:0] data_out_org359;
  output [9:0] data_out_org360;
  wire [9:0] data_out_org360;
  output [9:0] data_out_org361;
  wire [9:0] data_out_org361;
  output [9:0] data_out_org362;
  wire [9:0] data_out_org362;
  output [9:0] data_out_org363;
  wire [9:0] data_out_org363;
  output [9:0] data_out_org364;
  wire [9:0] data_out_org364;
  output [9:0] data_out_org365;
  wire [9:0] data_out_org365;
  output [9:0] data_out_org366;
  wire [9:0] data_out_org366;
  output [9:0] data_out_org367;
  wire [9:0] data_out_org367;
  output [9:0] data_out_org368;
  wire [9:0] data_out_org368;
  output [9:0] data_out_org369;
  wire [9:0] data_out_org369;
  output [9:0] data_out_org370;
  wire [9:0] data_out_org370;
  output [9:0] data_out_org371;
  wire [9:0] data_out_org371;
  output [9:0] data_out_org372;
  wire [9:0] data_out_org372;
  output [9:0] data_out_org373;
  wire [9:0] data_out_org373;
  output [9:0] data_out_org374;
  wire [9:0] data_out_org374;
  output [9:0] data_out_org375;
  wire [9:0] data_out_org375;
  output [9:0] data_out_org376;
  wire [9:0] data_out_org376;
  output [9:0] data_out_org377;
  wire [9:0] data_out_org377;
  output [9:0] data_out_org378;
  wire [9:0] data_out_org378;
  output [9:0] data_out_org379;
  wire [9:0] data_out_org379;
  output [9:0] data_out_org380;
  wire [9:0] data_out_org380;
  output [9:0] data_out_org381;
  wire [9:0] data_out_org381;
  output [9:0] data_out_org382;
  wire [9:0] data_out_org382;
  output [9:0] data_out_org385;
  wire [9:0] data_out_org385;
  output [9:0] data_out_org386;
  wire [9:0] data_out_org386;
  output [9:0] data_out_org387;
  wire [9:0] data_out_org387;
  output [9:0] data_out_org388;
  wire [9:0] data_out_org388;
  output [9:0] data_out_org389;
  wire [9:0] data_out_org389;
  output [9:0] data_out_org390;
  wire [9:0] data_out_org390;
  output [9:0] data_out_org391;
  wire [9:0] data_out_org391;
  output [9:0] data_out_org392;
  wire [9:0] data_out_org392;
  output [9:0] data_out_org393;
  wire [9:0] data_out_org393;
  output [9:0] data_out_org394;
  wire [9:0] data_out_org394;
  output [9:0] data_out_org395;
  wire [9:0] data_out_org395;
  output [9:0] data_out_org396;
  wire [9:0] data_out_org396;
  output [9:0] data_out_org397;
  wire [9:0] data_out_org397;
  output [9:0] data_out_org398;
  wire [9:0] data_out_org398;
  output [9:0] data_out_org399;
  wire [9:0] data_out_org399;
  output [9:0] data_out_org400;
  wire [9:0] data_out_org400;
  output [9:0] data_out_org401;
  wire [9:0] data_out_org401;
  output [9:0] data_out_org402;
  wire [9:0] data_out_org402;
  output [9:0] data_out_org403;
  wire [9:0] data_out_org403;
  output [9:0] data_out_org404;
  wire [9:0] data_out_org404;
  output [9:0] data_out_org405;
  wire [9:0] data_out_org405;
  output [9:0] data_out_org406;
  wire [9:0] data_out_org406;
  output [9:0] data_out_org407;
  wire [9:0] data_out_org407;
  output [9:0] data_out_org408;
  wire [9:0] data_out_org408;
  output [9:0] data_out_org409;
  wire [9:0] data_out_org409;
  output [9:0] data_out_org410;
  wire [9:0] data_out_org410;
  output [9:0] data_out_org411;
  wire [9:0] data_out_org411;
  output [9:0] data_out_org412;
  wire [9:0] data_out_org412;
  output [9:0] data_out_org413;
  wire [9:0] data_out_org413;
  output [9:0] data_out_org414;
  wire [9:0] data_out_org414;
  output [9:0] data_out_org417;
  wire [9:0] data_out_org417;
  output [9:0] data_out_org418;
  wire [9:0] data_out_org418;
  output [9:0] data_out_org419;
  wire [9:0] data_out_org419;
  output [9:0] data_out_org420;
  wire [9:0] data_out_org420;
  output [9:0] data_out_org421;
  wire [9:0] data_out_org421;
  output [9:0] data_out_org422;
  wire [9:0] data_out_org422;
  output [9:0] data_out_org423;
  wire [9:0] data_out_org423;
  output [9:0] data_out_org424;
  wire [9:0] data_out_org424;
  output [9:0] data_out_org425;
  wire [9:0] data_out_org425;
  output [9:0] data_out_org426;
  wire [9:0] data_out_org426;
  output [9:0] data_out_org427;
  wire [9:0] data_out_org427;
  output [9:0] data_out_org428;
  wire [9:0] data_out_org428;
  output [9:0] data_out_org429;
  wire [9:0] data_out_org429;
  output [9:0] data_out_org430;
  wire [9:0] data_out_org430;
  output [9:0] data_out_org431;
  wire [9:0] data_out_org431;
  output [9:0] data_out_org432;
  wire [9:0] data_out_org432;
  output [9:0] data_out_org433;
  wire [9:0] data_out_org433;
  output [9:0] data_out_org434;
  wire [9:0] data_out_org434;
  output [9:0] data_out_org435;
  wire [9:0] data_out_org435;
  output [9:0] data_out_org436;
  wire [9:0] data_out_org436;
  output [9:0] data_out_org437;
  wire [9:0] data_out_org437;
  output [9:0] data_out_org438;
  wire [9:0] data_out_org438;
  output [9:0] data_out_org439;
  wire [9:0] data_out_org439;
  output [9:0] data_out_org440;
  wire [9:0] data_out_org440;
  output [9:0] data_out_org441;
  wire [9:0] data_out_org441;
  output [9:0] data_out_org442;
  wire [9:0] data_out_org442;
  output [9:0] data_out_org443;
  wire [9:0] data_out_org443;
  output [9:0] data_out_org444;
  wire [9:0] data_out_org444;
  output [9:0] data_out_org445;
  wire [9:0] data_out_org445;
  output [9:0] data_out_org446;
  wire [9:0] data_out_org446;
  output [9:0] data_out_org449;
  wire [9:0] data_out_org449;
  output [9:0] data_out_org450;
  wire [9:0] data_out_org450;
  output [9:0] data_out_org451;
  wire [9:0] data_out_org451;
  output [9:0] data_out_org452;
  wire [9:0] data_out_org452;
  output [9:0] data_out_org453;
  wire [9:0] data_out_org453;
  output [9:0] data_out_org454;
  wire [9:0] data_out_org454;
  output [9:0] data_out_org455;
  wire [9:0] data_out_org455;
  output [9:0] data_out_org456;
  wire [9:0] data_out_org456;
  output [9:0] data_out_org457;
  wire [9:0] data_out_org457;
  output [9:0] data_out_org458;
  wire [9:0] data_out_org458;
  output [9:0] data_out_org459;
  wire [9:0] data_out_org459;
  output [9:0] data_out_org460;
  wire [9:0] data_out_org460;
  output [9:0] data_out_org461;
  wire [9:0] data_out_org461;
  output [9:0] data_out_org462;
  wire [9:0] data_out_org462;
  output [9:0] data_out_org463;
  wire [9:0] data_out_org463;
  output [9:0] data_out_org464;
  wire [9:0] data_out_org464;
  output [9:0] data_out_org465;
  wire [9:0] data_out_org465;
  output [9:0] data_out_org466;
  wire [9:0] data_out_org466;
  output [9:0] data_out_org467;
  wire [9:0] data_out_org467;
  output [9:0] data_out_org468;
  wire [9:0] data_out_org468;
  output [9:0] data_out_org469;
  wire [9:0] data_out_org469;
  output [9:0] data_out_org470;
  wire [9:0] data_out_org470;
  output [9:0] data_out_org471;
  wire [9:0] data_out_org471;
  output [9:0] data_out_org472;
  wire [9:0] data_out_org472;
  output [9:0] data_out_org473;
  wire [9:0] data_out_org473;
  output [9:0] data_out_org474;
  wire [9:0] data_out_org474;
  output [9:0] data_out_org475;
  wire [9:0] data_out_org475;
  output [9:0] data_out_org476;
  wire [9:0] data_out_org476;
  output [9:0] data_out_org477;
  wire [9:0] data_out_org477;
  output [9:0] data_out_org478;
  wire [9:0] data_out_org478;
  input [9:0] data_in_org33;
  wire [9:0] data_in_org33;
  input [9:0] data_in_org34;
  wire [9:0] data_in_org34;
  input [9:0] data_in_org35;
  wire [9:0] data_in_org35;
  input [9:0] data_in_org36;
  wire [9:0] data_in_org36;
  input [9:0] data_in_org37;
  wire [9:0] data_in_org37;
  input [9:0] data_in_org38;
  wire [9:0] data_in_org38;
  input [9:0] data_in_org39;
  wire [9:0] data_in_org39;
  input [9:0] data_in_org40;
  wire [9:0] data_in_org40;
  input [9:0] data_in_org41;
  wire [9:0] data_in_org41;
  input [9:0] data_in_org42;
  wire [9:0] data_in_org42;
  input [9:0] data_in_org43;
  wire [9:0] data_in_org43;
  input [9:0] data_in_org44;
  wire [9:0] data_in_org44;
  input [9:0] data_in_org45;
  wire [9:0] data_in_org45;
  input [9:0] data_in_org46;
  wire [9:0] data_in_org46;
  input [9:0] data_in_org47;
  wire [9:0] data_in_org47;
  input [9:0] data_in_org48;
  wire [9:0] data_in_org48;
  input [9:0] data_in_org49;
  wire [9:0] data_in_org49;
  input [9:0] data_in_org50;
  wire [9:0] data_in_org50;
  input [9:0] data_in_org51;
  wire [9:0] data_in_org51;
  input [9:0] data_in_org52;
  wire [9:0] data_in_org52;
  input [9:0] data_in_org53;
  wire [9:0] data_in_org53;
  input [9:0] data_in_org54;
  wire [9:0] data_in_org54;
  input [9:0] data_in_org55;
  wire [9:0] data_in_org55;
  input [9:0] data_in_org56;
  wire [9:0] data_in_org56;
  input [9:0] data_in_org57;
  wire [9:0] data_in_org57;
  input [9:0] data_in_org58;
  wire [9:0] data_in_org58;
  input [9:0] data_in_org59;
  wire [9:0] data_in_org59;
  input [9:0] data_in_org60;
  wire [9:0] data_in_org60;
  input [9:0] data_in_org61;
  wire [9:0] data_in_org61;
  input [9:0] data_in_org62;
  wire [9:0] data_in_org62;
  input [9:0] data_in_org65;
  wire [9:0] data_in_org65;
  input [9:0] data_in_org66;
  wire [9:0] data_in_org66;
  input [9:0] data_in_org67;
  wire [9:0] data_in_org67;
  input [9:0] data_in_org68;
  wire [9:0] data_in_org68;
  input [9:0] data_in_org69;
  wire [9:0] data_in_org69;
  input [9:0] data_in_org70;
  wire [9:0] data_in_org70;
  input [9:0] data_in_org71;
  wire [9:0] data_in_org71;
  input [9:0] data_in_org72;
  wire [9:0] data_in_org72;
  input [9:0] data_in_org73;
  wire [9:0] data_in_org73;
  input [9:0] data_in_org74;
  wire [9:0] data_in_org74;
  input [9:0] data_in_org75;
  wire [9:0] data_in_org75;
  input [9:0] data_in_org76;
  wire [9:0] data_in_org76;
  input [9:0] data_in_org77;
  wire [9:0] data_in_org77;
  input [9:0] data_in_org78;
  wire [9:0] data_in_org78;
  input [9:0] data_in_org79;
  wire [9:0] data_in_org79;
  input [9:0] data_in_org80;
  wire [9:0] data_in_org80;
  input [9:0] data_in_org81;
  wire [9:0] data_in_org81;
  input [9:0] data_in_org82;
  wire [9:0] data_in_org82;
  input [9:0] data_in_org83;
  wire [9:0] data_in_org83;
  input [9:0] data_in_org84;
  wire [9:0] data_in_org84;
  input [9:0] data_in_org85;
  wire [9:0] data_in_org85;
  input [9:0] data_in_org86;
  wire [9:0] data_in_org86;
  input [9:0] data_in_org87;
  wire [9:0] data_in_org87;
  input [9:0] data_in_org88;
  wire [9:0] data_in_org88;
  input [9:0] data_in_org89;
  wire [9:0] data_in_org89;
  input [9:0] data_in_org90;
  wire [9:0] data_in_org90;
  input [9:0] data_in_org91;
  wire [9:0] data_in_org91;
  input [9:0] data_in_org92;
  wire [9:0] data_in_org92;
  input [9:0] data_in_org93;
  wire [9:0] data_in_org93;
  input [9:0] data_in_org94;
  wire [9:0] data_in_org94;
  input [9:0] data_in_org97;
  wire [9:0] data_in_org97;
  input [9:0] data_in_org98;
  wire [9:0] data_in_org98;
  input [9:0] data_in_org99;
  wire [9:0] data_in_org99;
  input [9:0] data_in_org100;
  wire [9:0] data_in_org100;
  input [9:0] data_in_org101;
  wire [9:0] data_in_org101;
  input [9:0] data_in_org102;
  wire [9:0] data_in_org102;
  input [9:0] data_in_org103;
  wire [9:0] data_in_org103;
  input [9:0] data_in_org104;
  wire [9:0] data_in_org104;
  input [9:0] data_in_org105;
  wire [9:0] data_in_org105;
  input [9:0] data_in_org106;
  wire [9:0] data_in_org106;
  input [9:0] data_in_org107;
  wire [9:0] data_in_org107;
  input [9:0] data_in_org108;
  wire [9:0] data_in_org108;
  input [9:0] data_in_org109;
  wire [9:0] data_in_org109;
  input [9:0] data_in_org110;
  wire [9:0] data_in_org110;
  input [9:0] data_in_org111;
  wire [9:0] data_in_org111;
  input [9:0] data_in_org112;
  wire [9:0] data_in_org112;
  input [9:0] data_in_org113;
  wire [9:0] data_in_org113;
  input [9:0] data_in_org114;
  wire [9:0] data_in_org114;
  input [9:0] data_in_org115;
  wire [9:0] data_in_org115;
  input [9:0] data_in_org116;
  wire [9:0] data_in_org116;
  input [9:0] data_in_org117;
  wire [9:0] data_in_org117;
  input [9:0] data_in_org118;
  wire [9:0] data_in_org118;
  input [9:0] data_in_org119;
  wire [9:0] data_in_org119;
  input [9:0] data_in_org120;
  wire [9:0] data_in_org120;
  input [9:0] data_in_org121;
  wire [9:0] data_in_org121;
  input [9:0] data_in_org122;
  wire [9:0] data_in_org122;
  input [9:0] data_in_org123;
  wire [9:0] data_in_org123;
  input [9:0] data_in_org124;
  wire [9:0] data_in_org124;
  input [9:0] data_in_org125;
  wire [9:0] data_in_org125;
  input [9:0] data_in_org126;
  wire [9:0] data_in_org126;
  input [9:0] data_in_org129;
  wire [9:0] data_in_org129;
  input [9:0] data_in_org130;
  wire [9:0] data_in_org130;
  input [9:0] data_in_org131;
  wire [9:0] data_in_org131;
  input [9:0] data_in_org132;
  wire [9:0] data_in_org132;
  input [9:0] data_in_org133;
  wire [9:0] data_in_org133;
  input [9:0] data_in_org134;
  wire [9:0] data_in_org134;
  input [9:0] data_in_org135;
  wire [9:0] data_in_org135;
  input [9:0] data_in_org136;
  wire [9:0] data_in_org136;
  input [9:0] data_in_org137;
  wire [9:0] data_in_org137;
  input [9:0] data_in_org138;
  wire [9:0] data_in_org138;
  input [9:0] data_in_org139;
  wire [9:0] data_in_org139;
  input [9:0] data_in_org140;
  wire [9:0] data_in_org140;
  input [9:0] data_in_org141;
  wire [9:0] data_in_org141;
  input [9:0] data_in_org142;
  wire [9:0] data_in_org142;
  input [9:0] data_in_org143;
  wire [9:0] data_in_org143;
  input [9:0] data_in_org144;
  wire [9:0] data_in_org144;
  input [9:0] data_in_org145;
  wire [9:0] data_in_org145;
  input [9:0] data_in_org146;
  wire [9:0] data_in_org146;
  input [9:0] data_in_org147;
  wire [9:0] data_in_org147;
  input [9:0] data_in_org148;
  wire [9:0] data_in_org148;
  input [9:0] data_in_org149;
  wire [9:0] data_in_org149;
  input [9:0] data_in_org150;
  wire [9:0] data_in_org150;
  input [9:0] data_in_org151;
  wire [9:0] data_in_org151;
  input [9:0] data_in_org152;
  wire [9:0] data_in_org152;
  input [9:0] data_in_org153;
  wire [9:0] data_in_org153;
  input [9:0] data_in_org154;
  wire [9:0] data_in_org154;
  input [9:0] data_in_org155;
  wire [9:0] data_in_org155;
  input [9:0] data_in_org156;
  wire [9:0] data_in_org156;
  input [9:0] data_in_org157;
  wire [9:0] data_in_org157;
  input [9:0] data_in_org158;
  wire [9:0] data_in_org158;
  input [9:0] data_in_org161;
  wire [9:0] data_in_org161;
  input [9:0] data_in_org162;
  wire [9:0] data_in_org162;
  input [9:0] data_in_org163;
  wire [9:0] data_in_org163;
  input [9:0] data_in_org164;
  wire [9:0] data_in_org164;
  input [9:0] data_in_org165;
  wire [9:0] data_in_org165;
  input [9:0] data_in_org166;
  wire [9:0] data_in_org166;
  input [9:0] data_in_org167;
  wire [9:0] data_in_org167;
  input [9:0] data_in_org168;
  wire [9:0] data_in_org168;
  input [9:0] data_in_org169;
  wire [9:0] data_in_org169;
  input [9:0] data_in_org170;
  wire [9:0] data_in_org170;
  input [9:0] data_in_org171;
  wire [9:0] data_in_org171;
  input [9:0] data_in_org172;
  wire [9:0] data_in_org172;
  input [9:0] data_in_org173;
  wire [9:0] data_in_org173;
  input [9:0] data_in_org174;
  wire [9:0] data_in_org174;
  input [9:0] data_in_org175;
  wire [9:0] data_in_org175;
  input [9:0] data_in_org176;
  wire [9:0] data_in_org176;
  input [9:0] data_in_org177;
  wire [9:0] data_in_org177;
  input [9:0] data_in_org178;
  wire [9:0] data_in_org178;
  input [9:0] data_in_org179;
  wire [9:0] data_in_org179;
  input [9:0] data_in_org180;
  wire [9:0] data_in_org180;
  input [9:0] data_in_org181;
  wire [9:0] data_in_org181;
  input [9:0] data_in_org182;
  wire [9:0] data_in_org182;
  input [9:0] data_in_org183;
  wire [9:0] data_in_org183;
  input [9:0] data_in_org184;
  wire [9:0] data_in_org184;
  input [9:0] data_in_org185;
  wire [9:0] data_in_org185;
  input [9:0] data_in_org186;
  wire [9:0] data_in_org186;
  input [9:0] data_in_org187;
  wire [9:0] data_in_org187;
  input [9:0] data_in_org188;
  wire [9:0] data_in_org188;
  input [9:0] data_in_org189;
  wire [9:0] data_in_org189;
  input [9:0] data_in_org190;
  wire [9:0] data_in_org190;
  input [9:0] data_in_org193;
  wire [9:0] data_in_org193;
  input [9:0] data_in_org194;
  wire [9:0] data_in_org194;
  input [9:0] data_in_org195;
  wire [9:0] data_in_org195;
  input [9:0] data_in_org196;
  wire [9:0] data_in_org196;
  input [9:0] data_in_org197;
  wire [9:0] data_in_org197;
  input [9:0] data_in_org198;
  wire [9:0] data_in_org198;
  input [9:0] data_in_org199;
  wire [9:0] data_in_org199;
  input [9:0] data_in_org200;
  wire [9:0] data_in_org200;
  input [9:0] data_in_org201;
  wire [9:0] data_in_org201;
  input [9:0] data_in_org202;
  wire [9:0] data_in_org202;
  input [9:0] data_in_org203;
  wire [9:0] data_in_org203;
  input [9:0] data_in_org204;
  wire [9:0] data_in_org204;
  input [9:0] data_in_org205;
  wire [9:0] data_in_org205;
  input [9:0] data_in_org206;
  wire [9:0] data_in_org206;
  input [9:0] data_in_org207;
  wire [9:0] data_in_org207;
  input [9:0] data_in_org208;
  wire [9:0] data_in_org208;
  input [9:0] data_in_org209;
  wire [9:0] data_in_org209;
  input [9:0] data_in_org210;
  wire [9:0] data_in_org210;
  input [9:0] data_in_org211;
  wire [9:0] data_in_org211;
  input [9:0] data_in_org212;
  wire [9:0] data_in_org212;
  input [9:0] data_in_org213;
  wire [9:0] data_in_org213;
  input [9:0] data_in_org214;
  wire [9:0] data_in_org214;
  input [9:0] data_in_org215;
  wire [9:0] data_in_org215;
  input [9:0] data_in_org216;
  wire [9:0] data_in_org216;
  input [9:0] data_in_org217;
  wire [9:0] data_in_org217;
  input [9:0] data_in_org218;
  wire [9:0] data_in_org218;
  input [9:0] data_in_org219;
  wire [9:0] data_in_org219;
  input [9:0] data_in_org220;
  wire [9:0] data_in_org220;
  input [9:0] data_in_org221;
  wire [9:0] data_in_org221;
  input [9:0] data_in_org222;
  wire [9:0] data_in_org222;
  input [9:0] data_in_org225;
  wire [9:0] data_in_org225;
  input [9:0] data_in_org226;
  wire [9:0] data_in_org226;
  input [9:0] data_in_org227;
  wire [9:0] data_in_org227;
  input [9:0] data_in_org228;
  wire [9:0] data_in_org228;
  input [9:0] data_in_org229;
  wire [9:0] data_in_org229;
  input [9:0] data_in_org230;
  wire [9:0] data_in_org230;
  input [9:0] data_in_org231;
  wire [9:0] data_in_org231;
  input [9:0] data_in_org232;
  wire [9:0] data_in_org232;
  input [9:0] data_in_org233;
  wire [9:0] data_in_org233;
  input [9:0] data_in_org234;
  wire [9:0] data_in_org234;
  input [9:0] data_in_org235;
  wire [9:0] data_in_org235;
  input [9:0] data_in_org236;
  wire [9:0] data_in_org236;
  input [9:0] data_in_org237;
  wire [9:0] data_in_org237;
  input [9:0] data_in_org238;
  wire [9:0] data_in_org238;
  input [9:0] data_in_org239;
  wire [9:0] data_in_org239;
  input [9:0] data_in_org240;
  wire [9:0] data_in_org240;
  input [9:0] data_in_org241;
  wire [9:0] data_in_org241;
  input [9:0] data_in_org242;
  wire [9:0] data_in_org242;
  input [9:0] data_in_org243;
  wire [9:0] data_in_org243;
  input [9:0] data_in_org244;
  wire [9:0] data_in_org244;
  input [9:0] data_in_org245;
  wire [9:0] data_in_org245;
  input [9:0] data_in_org246;
  wire [9:0] data_in_org246;
  input [9:0] data_in_org247;
  wire [9:0] data_in_org247;
  input [9:0] data_in_org248;
  wire [9:0] data_in_org248;
  input [9:0] data_in_org249;
  wire [9:0] data_in_org249;
  input [9:0] data_in_org250;
  wire [9:0] data_in_org250;
  input [9:0] data_in_org251;
  wire [9:0] data_in_org251;
  input [9:0] data_in_org252;
  wire [9:0] data_in_org252;
  input [9:0] data_in_org253;
  wire [9:0] data_in_org253;
  input [9:0] data_in_org254;
  wire [9:0] data_in_org254;
  input [9:0] data_in_org257;
  wire [9:0] data_in_org257;
  input [9:0] data_in_org258;
  wire [9:0] data_in_org258;
  input [9:0] data_in_org259;
  wire [9:0] data_in_org259;
  input [9:0] data_in_org260;
  wire [9:0] data_in_org260;
  input [9:0] data_in_org261;
  wire [9:0] data_in_org261;
  input [9:0] data_in_org262;
  wire [9:0] data_in_org262;
  input [9:0] data_in_org263;
  wire [9:0] data_in_org263;
  input [9:0] data_in_org264;
  wire [9:0] data_in_org264;
  input [9:0] data_in_org265;
  wire [9:0] data_in_org265;
  input [9:0] data_in_org266;
  wire [9:0] data_in_org266;
  input [9:0] data_in_org267;
  wire [9:0] data_in_org267;
  input [9:0] data_in_org268;
  wire [9:0] data_in_org268;
  input [9:0] data_in_org269;
  wire [9:0] data_in_org269;
  input [9:0] data_in_org270;
  wire [9:0] data_in_org270;
  input [9:0] data_in_org271;
  wire [9:0] data_in_org271;
  input [9:0] data_in_org272;
  wire [9:0] data_in_org272;
  input [9:0] data_in_org273;
  wire [9:0] data_in_org273;
  input [9:0] data_in_org274;
  wire [9:0] data_in_org274;
  input [9:0] data_in_org275;
  wire [9:0] data_in_org275;
  input [9:0] data_in_org276;
  wire [9:0] data_in_org276;
  input [9:0] data_in_org277;
  wire [9:0] data_in_org277;
  input [9:0] data_in_org278;
  wire [9:0] data_in_org278;
  input [9:0] data_in_org279;
  wire [9:0] data_in_org279;
  input [9:0] data_in_org280;
  wire [9:0] data_in_org280;
  input [9:0] data_in_org281;
  wire [9:0] data_in_org281;
  input [9:0] data_in_org282;
  wire [9:0] data_in_org282;
  input [9:0] data_in_org283;
  wire [9:0] data_in_org283;
  input [9:0] data_in_org284;
  wire [9:0] data_in_org284;
  input [9:0] data_in_org285;
  wire [9:0] data_in_org285;
  input [9:0] data_in_org286;
  wire [9:0] data_in_org286;
  input [9:0] data_in_org289;
  wire [9:0] data_in_org289;
  input [9:0] data_in_org290;
  wire [9:0] data_in_org290;
  input [9:0] data_in_org291;
  wire [9:0] data_in_org291;
  input [9:0] data_in_org292;
  wire [9:0] data_in_org292;
  input [9:0] data_in_org293;
  wire [9:0] data_in_org293;
  input [9:0] data_in_org294;
  wire [9:0] data_in_org294;
  input [9:0] data_in_org295;
  wire [9:0] data_in_org295;
  input [9:0] data_in_org296;
  wire [9:0] data_in_org296;
  input [9:0] data_in_org297;
  wire [9:0] data_in_org297;
  input [9:0] data_in_org298;
  wire [9:0] data_in_org298;
  input [9:0] data_in_org299;
  wire [9:0] data_in_org299;
  input [9:0] data_in_org300;
  wire [9:0] data_in_org300;
  input [9:0] data_in_org301;
  wire [9:0] data_in_org301;
  input [9:0] data_in_org302;
  wire [9:0] data_in_org302;
  input [9:0] data_in_org303;
  wire [9:0] data_in_org303;
  input [9:0] data_in_org304;
  wire [9:0] data_in_org304;
  input [9:0] data_in_org305;
  wire [9:0] data_in_org305;
  input [9:0] data_in_org306;
  wire [9:0] data_in_org306;
  input [9:0] data_in_org307;
  wire [9:0] data_in_org307;
  input [9:0] data_in_org308;
  wire [9:0] data_in_org308;
  input [9:0] data_in_org309;
  wire [9:0] data_in_org309;
  input [9:0] data_in_org310;
  wire [9:0] data_in_org310;
  input [9:0] data_in_org311;
  wire [9:0] data_in_org311;
  input [9:0] data_in_org312;
  wire [9:0] data_in_org312;
  input [9:0] data_in_org313;
  wire [9:0] data_in_org313;
  input [9:0] data_in_org314;
  wire [9:0] data_in_org314;
  input [9:0] data_in_org315;
  wire [9:0] data_in_org315;
  input [9:0] data_in_org316;
  wire [9:0] data_in_org316;
  input [9:0] data_in_org317;
  wire [9:0] data_in_org317;
  input [9:0] data_in_org318;
  wire [9:0] data_in_org318;
  input [9:0] data_in_org321;
  wire [9:0] data_in_org321;
  input [9:0] data_in_org322;
  wire [9:0] data_in_org322;
  input [9:0] data_in_org323;
  wire [9:0] data_in_org323;
  input [9:0] data_in_org324;
  wire [9:0] data_in_org324;
  input [9:0] data_in_org325;
  wire [9:0] data_in_org325;
  input [9:0] data_in_org326;
  wire [9:0] data_in_org326;
  input [9:0] data_in_org327;
  wire [9:0] data_in_org327;
  input [9:0] data_in_org328;
  wire [9:0] data_in_org328;
  input [9:0] data_in_org329;
  wire [9:0] data_in_org329;
  input [9:0] data_in_org330;
  wire [9:0] data_in_org330;
  input [9:0] data_in_org331;
  wire [9:0] data_in_org331;
  input [9:0] data_in_org332;
  wire [9:0] data_in_org332;
  input [9:0] data_in_org333;
  wire [9:0] data_in_org333;
  input [9:0] data_in_org334;
  wire [9:0] data_in_org334;
  input [9:0] data_in_org335;
  wire [9:0] data_in_org335;
  input [9:0] data_in_org336;
  wire [9:0] data_in_org336;
  input [9:0] data_in_org337;
  wire [9:0] data_in_org337;
  input [9:0] data_in_org338;
  wire [9:0] data_in_org338;
  input [9:0] data_in_org339;
  wire [9:0] data_in_org339;
  input [9:0] data_in_org340;
  wire [9:0] data_in_org340;
  input [9:0] data_in_org341;
  wire [9:0] data_in_org341;
  input [9:0] data_in_org342;
  wire [9:0] data_in_org342;
  input [9:0] data_in_org343;
  wire [9:0] data_in_org343;
  input [9:0] data_in_org344;
  wire [9:0] data_in_org344;
  input [9:0] data_in_org345;
  wire [9:0] data_in_org345;
  input [9:0] data_in_org346;
  wire [9:0] data_in_org346;
  input [9:0] data_in_org347;
  wire [9:0] data_in_org347;
  input [9:0] data_in_org348;
  wire [9:0] data_in_org348;
  input [9:0] data_in_org349;
  wire [9:0] data_in_org349;
  input [9:0] data_in_org350;
  wire [9:0] data_in_org350;
  input [9:0] data_in_org353;
  wire [9:0] data_in_org353;
  input [9:0] data_in_org354;
  wire [9:0] data_in_org354;
  input [9:0] data_in_org355;
  wire [9:0] data_in_org355;
  input [9:0] data_in_org356;
  wire [9:0] data_in_org356;
  input [9:0] data_in_org357;
  wire [9:0] data_in_org357;
  input [9:0] data_in_org358;
  wire [9:0] data_in_org358;
  input [9:0] data_in_org359;
  wire [9:0] data_in_org359;
  input [9:0] data_in_org360;
  wire [9:0] data_in_org360;
  input [9:0] data_in_org361;
  wire [9:0] data_in_org361;
  input [9:0] data_in_org362;
  wire [9:0] data_in_org362;
  input [9:0] data_in_org363;
  wire [9:0] data_in_org363;
  input [9:0] data_in_org364;
  wire [9:0] data_in_org364;
  input [9:0] data_in_org365;
  wire [9:0] data_in_org365;
  input [9:0] data_in_org366;
  wire [9:0] data_in_org366;
  input [9:0] data_in_org367;
  wire [9:0] data_in_org367;
  input [9:0] data_in_org368;
  wire [9:0] data_in_org368;
  input [9:0] data_in_org369;
  wire [9:0] data_in_org369;
  input [9:0] data_in_org370;
  wire [9:0] data_in_org370;
  input [9:0] data_in_org371;
  wire [9:0] data_in_org371;
  input [9:0] data_in_org372;
  wire [9:0] data_in_org372;
  input [9:0] data_in_org373;
  wire [9:0] data_in_org373;
  input [9:0] data_in_org374;
  wire [9:0] data_in_org374;
  input [9:0] data_in_org375;
  wire [9:0] data_in_org375;
  input [9:0] data_in_org376;
  wire [9:0] data_in_org376;
  input [9:0] data_in_org377;
  wire [9:0] data_in_org377;
  input [9:0] data_in_org378;
  wire [9:0] data_in_org378;
  input [9:0] data_in_org379;
  wire [9:0] data_in_org379;
  input [9:0] data_in_org380;
  wire [9:0] data_in_org380;
  input [9:0] data_in_org381;
  wire [9:0] data_in_org381;
  input [9:0] data_in_org382;
  wire [9:0] data_in_org382;
  input [9:0] data_in_org385;
  wire [9:0] data_in_org385;
  input [9:0] data_in_org386;
  wire [9:0] data_in_org386;
  input [9:0] data_in_org387;
  wire [9:0] data_in_org387;
  input [9:0] data_in_org388;
  wire [9:0] data_in_org388;
  input [9:0] data_in_org389;
  wire [9:0] data_in_org389;
  input [9:0] data_in_org390;
  wire [9:0] data_in_org390;
  input [9:0] data_in_org391;
  wire [9:0] data_in_org391;
  input [9:0] data_in_org392;
  wire [9:0] data_in_org392;
  input [9:0] data_in_org393;
  wire [9:0] data_in_org393;
  input [9:0] data_in_org394;
  wire [9:0] data_in_org394;
  input [9:0] data_in_org395;
  wire [9:0] data_in_org395;
  input [9:0] data_in_org396;
  wire [9:0] data_in_org396;
  input [9:0] data_in_org397;
  wire [9:0] data_in_org397;
  input [9:0] data_in_org398;
  wire [9:0] data_in_org398;
  input [9:0] data_in_org399;
  wire [9:0] data_in_org399;
  input [9:0] data_in_org400;
  wire [9:0] data_in_org400;
  input [9:0] data_in_org401;
  wire [9:0] data_in_org401;
  input [9:0] data_in_org402;
  wire [9:0] data_in_org402;
  input [9:0] data_in_org403;
  wire [9:0] data_in_org403;
  input [9:0] data_in_org404;
  wire [9:0] data_in_org404;
  input [9:0] data_in_org405;
  wire [9:0] data_in_org405;
  input [9:0] data_in_org406;
  wire [9:0] data_in_org406;
  input [9:0] data_in_org407;
  wire [9:0] data_in_org407;
  input [9:0] data_in_org408;
  wire [9:0] data_in_org408;
  input [9:0] data_in_org409;
  wire [9:0] data_in_org409;
  input [9:0] data_in_org410;
  wire [9:0] data_in_org410;
  input [9:0] data_in_org411;
  wire [9:0] data_in_org411;
  input [9:0] data_in_org412;
  wire [9:0] data_in_org412;
  input [9:0] data_in_org413;
  wire [9:0] data_in_org413;
  input [9:0] data_in_org414;
  wire [9:0] data_in_org414;
  input [9:0] data_in_org417;
  wire [9:0] data_in_org417;
  input [9:0] data_in_org418;
  wire [9:0] data_in_org418;
  input [9:0] data_in_org419;
  wire [9:0] data_in_org419;
  input [9:0] data_in_org420;
  wire [9:0] data_in_org420;
  input [9:0] data_in_org421;
  wire [9:0] data_in_org421;
  input [9:0] data_in_org422;
  wire [9:0] data_in_org422;
  input [9:0] data_in_org423;
  wire [9:0] data_in_org423;
  input [9:0] data_in_org424;
  wire [9:0] data_in_org424;
  input [9:0] data_in_org425;
  wire [9:0] data_in_org425;
  input [9:0] data_in_org426;
  wire [9:0] data_in_org426;
  input [9:0] data_in_org427;
  wire [9:0] data_in_org427;
  input [9:0] data_in_org428;
  wire [9:0] data_in_org428;
  input [9:0] data_in_org429;
  wire [9:0] data_in_org429;
  input [9:0] data_in_org430;
  wire [9:0] data_in_org430;
  input [9:0] data_in_org431;
  wire [9:0] data_in_org431;
  input [9:0] data_in_org432;
  wire [9:0] data_in_org432;
  input [9:0] data_in_org433;
  wire [9:0] data_in_org433;
  input [9:0] data_in_org434;
  wire [9:0] data_in_org434;
  input [9:0] data_in_org435;
  wire [9:0] data_in_org435;
  input [9:0] data_in_org436;
  wire [9:0] data_in_org436;
  input [9:0] data_in_org437;
  wire [9:0] data_in_org437;
  input [9:0] data_in_org438;
  wire [9:0] data_in_org438;
  input [9:0] data_in_org439;
  wire [9:0] data_in_org439;
  input [9:0] data_in_org440;
  wire [9:0] data_in_org440;
  input [9:0] data_in_org441;
  wire [9:0] data_in_org441;
  input [9:0] data_in_org442;
  wire [9:0] data_in_org442;
  input [9:0] data_in_org443;
  wire [9:0] data_in_org443;
  input [9:0] data_in_org444;
  wire [9:0] data_in_org444;
  input [9:0] data_in_org445;
  wire [9:0] data_in_org445;
  input [9:0] data_in_org446;
  wire [9:0] data_in_org446;
  input [9:0] data_in_org449;
  wire [9:0] data_in_org449;
  input [9:0] data_in_org450;
  wire [9:0] data_in_org450;
  input [9:0] data_in_org451;
  wire [9:0] data_in_org451;
  input [9:0] data_in_org452;
  wire [9:0] data_in_org452;
  input [9:0] data_in_org453;
  wire [9:0] data_in_org453;
  input [9:0] data_in_org454;
  wire [9:0] data_in_org454;
  input [9:0] data_in_org455;
  wire [9:0] data_in_org455;
  input [9:0] data_in_org456;
  wire [9:0] data_in_org456;
  input [9:0] data_in_org457;
  wire [9:0] data_in_org457;
  input [9:0] data_in_org458;
  wire [9:0] data_in_org458;
  input [9:0] data_in_org459;
  wire [9:0] data_in_org459;
  input [9:0] data_in_org460;
  wire [9:0] data_in_org460;
  input [9:0] data_in_org461;
  wire [9:0] data_in_org461;
  input [9:0] data_in_org462;
  wire [9:0] data_in_org462;
  input [9:0] data_in_org463;
  wire [9:0] data_in_org463;
  input [9:0] data_in_org464;
  wire [9:0] data_in_org464;
  input [9:0] data_in_org465;
  wire [9:0] data_in_org465;
  input [9:0] data_in_org466;
  wire [9:0] data_in_org466;
  input [9:0] data_in_org467;
  wire [9:0] data_in_org467;
  input [9:0] data_in_org468;
  wire [9:0] data_in_org468;
  input [9:0] data_in_org469;
  wire [9:0] data_in_org469;
  input [9:0] data_in_org470;
  wire [9:0] data_in_org470;
  input [9:0] data_in_org471;
  wire [9:0] data_in_org471;
  input [9:0] data_in_org472;
  wire [9:0] data_in_org472;
  input [9:0] data_in_org473;
  wire [9:0] data_in_org473;
  input [9:0] data_in_org474;
  wire [9:0] data_in_org474;
  input [9:0] data_in_org475;
  wire [9:0] data_in_org475;
  input [9:0] data_in_org476;
  wire [9:0] data_in_org476;
  input [9:0] data_in_org477;
  wire [9:0] data_in_org477;
  input [9:0] data_in_org478;
  wire [9:0] data_in_org478;
  output [9:0] data_out33;
  wire [9:0] data_out33;
  output [9:0] data_out34;
  wire [9:0] data_out34;
  output [9:0] data_out35;
  wire [9:0] data_out35;
  output [9:0] data_out36;
  wire [9:0] data_out36;
  output [9:0] data_out37;
  wire [9:0] data_out37;
  output [9:0] data_out38;
  wire [9:0] data_out38;
  output [9:0] data_out39;
  wire [9:0] data_out39;
  output [9:0] data_out40;
  wire [9:0] data_out40;
  output [9:0] data_out41;
  wire [9:0] data_out41;
  output [9:0] data_out42;
  wire [9:0] data_out42;
  output [9:0] data_out43;
  wire [9:0] data_out43;
  output [9:0] data_out44;
  wire [9:0] data_out44;
  output [9:0] data_out45;
  wire [9:0] data_out45;
  output [9:0] data_out46;
  wire [9:0] data_out46;
  output [9:0] data_out47;
  wire [9:0] data_out47;
  output [9:0] data_out48;
  wire [9:0] data_out48;
  output [9:0] data_out49;
  wire [9:0] data_out49;
  output [9:0] data_out50;
  wire [9:0] data_out50;
  output [9:0] data_out51;
  wire [9:0] data_out51;
  output [9:0] data_out52;
  wire [9:0] data_out52;
  output [9:0] data_out53;
  wire [9:0] data_out53;
  output [9:0] data_out54;
  wire [9:0] data_out54;
  output [9:0] data_out55;
  wire [9:0] data_out55;
  output [9:0] data_out56;
  wire [9:0] data_out56;
  output [9:0] data_out57;
  wire [9:0] data_out57;
  output [9:0] data_out58;
  wire [9:0] data_out58;
  output [9:0] data_out59;
  wire [9:0] data_out59;
  output [9:0] data_out60;
  wire [9:0] data_out60;
  output [9:0] data_out61;
  wire [9:0] data_out61;
  output [9:0] data_out62;
  wire [9:0] data_out62;
  output [9:0] data_out65;
  wire [9:0] data_out65;
  output [9:0] data_out66;
  wire [9:0] data_out66;
  output [9:0] data_out67;
  wire [9:0] data_out67;
  output [9:0] data_out68;
  wire [9:0] data_out68;
  output [9:0] data_out69;
  wire [9:0] data_out69;
  output [9:0] data_out70;
  wire [9:0] data_out70;
  output [9:0] data_out71;
  wire [9:0] data_out71;
  output [9:0] data_out72;
  wire [9:0] data_out72;
  output [9:0] data_out73;
  wire [9:0] data_out73;
  output [9:0] data_out74;
  wire [9:0] data_out74;
  output [9:0] data_out75;
  wire [9:0] data_out75;
  output [9:0] data_out76;
  wire [9:0] data_out76;
  output [9:0] data_out77;
  wire [9:0] data_out77;
  output [9:0] data_out78;
  wire [9:0] data_out78;
  output [9:0] data_out79;
  wire [9:0] data_out79;
  output [9:0] data_out80;
  wire [9:0] data_out80;
  output [9:0] data_out81;
  wire [9:0] data_out81;
  output [9:0] data_out82;
  wire [9:0] data_out82;
  output [9:0] data_out83;
  wire [9:0] data_out83;
  output [9:0] data_out84;
  wire [9:0] data_out84;
  output [9:0] data_out85;
  wire [9:0] data_out85;
  output [9:0] data_out86;
  wire [9:0] data_out86;
  output [9:0] data_out87;
  wire [9:0] data_out87;
  output [9:0] data_out88;
  wire [9:0] data_out88;
  output [9:0] data_out89;
  wire [9:0] data_out89;
  output [9:0] data_out90;
  wire [9:0] data_out90;
  output [9:0] data_out91;
  wire [9:0] data_out91;
  output [9:0] data_out92;
  wire [9:0] data_out92;
  output [9:0] data_out93;
  wire [9:0] data_out93;
  output [9:0] data_out94;
  wire [9:0] data_out94;
  output [9:0] data_out97;
  wire [9:0] data_out97;
  output [9:0] data_out98;
  wire [9:0] data_out98;
  output [9:0] data_out99;
  wire [9:0] data_out99;
  output [9:0] data_out100;
  wire [9:0] data_out100;
  output [9:0] data_out101;
  wire [9:0] data_out101;
  output [9:0] data_out102;
  wire [9:0] data_out102;
  output [9:0] data_out103;
  wire [9:0] data_out103;
  output [9:0] data_out104;
  wire [9:0] data_out104;
  output [9:0] data_out105;
  wire [9:0] data_out105;
  output [9:0] data_out106;
  wire [9:0] data_out106;
  output [9:0] data_out107;
  wire [9:0] data_out107;
  output [9:0] data_out108;
  wire [9:0] data_out108;
  output [9:0] data_out109;
  wire [9:0] data_out109;
  output [9:0] data_out110;
  wire [9:0] data_out110;
  output [9:0] data_out111;
  wire [9:0] data_out111;
  output [9:0] data_out112;
  wire [9:0] data_out112;
  output [9:0] data_out113;
  wire [9:0] data_out113;
  output [9:0] data_out114;
  wire [9:0] data_out114;
  output [9:0] data_out115;
  wire [9:0] data_out115;
  output [9:0] data_out116;
  wire [9:0] data_out116;
  output [9:0] data_out117;
  wire [9:0] data_out117;
  output [9:0] data_out118;
  wire [9:0] data_out118;
  output [9:0] data_out119;
  wire [9:0] data_out119;
  output [9:0] data_out120;
  wire [9:0] data_out120;
  output [9:0] data_out121;
  wire [9:0] data_out121;
  output [9:0] data_out122;
  wire [9:0] data_out122;
  output [9:0] data_out123;
  wire [9:0] data_out123;
  output [9:0] data_out124;
  wire [9:0] data_out124;
  output [9:0] data_out125;
  wire [9:0] data_out125;
  output [9:0] data_out126;
  wire [9:0] data_out126;
  output [9:0] data_out129;
  wire [9:0] data_out129;
  output [9:0] data_out130;
  wire [9:0] data_out130;
  output [9:0] data_out131;
  wire [9:0] data_out131;
  output [9:0] data_out132;
  wire [9:0] data_out132;
  output [9:0] data_out133;
  wire [9:0] data_out133;
  output [9:0] data_out134;
  wire [9:0] data_out134;
  output [9:0] data_out135;
  wire [9:0] data_out135;
  output [9:0] data_out136;
  wire [9:0] data_out136;
  output [9:0] data_out137;
  wire [9:0] data_out137;
  output [9:0] data_out138;
  wire [9:0] data_out138;
  output [9:0] data_out139;
  wire [9:0] data_out139;
  output [9:0] data_out140;
  wire [9:0] data_out140;
  output [9:0] data_out141;
  wire [9:0] data_out141;
  output [9:0] data_out142;
  wire [9:0] data_out142;
  output [9:0] data_out143;
  wire [9:0] data_out143;
  output [9:0] data_out144;
  wire [9:0] data_out144;
  output [9:0] data_out145;
  wire [9:0] data_out145;
  output [9:0] data_out146;
  wire [9:0] data_out146;
  output [9:0] data_out147;
  wire [9:0] data_out147;
  output [9:0] data_out148;
  wire [9:0] data_out148;
  output [9:0] data_out149;
  wire [9:0] data_out149;
  output [9:0] data_out150;
  wire [9:0] data_out150;
  output [9:0] data_out151;
  wire [9:0] data_out151;
  output [9:0] data_out152;
  wire [9:0] data_out152;
  output [9:0] data_out153;
  wire [9:0] data_out153;
  output [9:0] data_out154;
  wire [9:0] data_out154;
  output [9:0] data_out155;
  wire [9:0] data_out155;
  output [9:0] data_out156;
  wire [9:0] data_out156;
  output [9:0] data_out157;
  wire [9:0] data_out157;
  output [9:0] data_out158;
  wire [9:0] data_out158;
  output [9:0] data_out161;
  wire [9:0] data_out161;
  output [9:0] data_out162;
  wire [9:0] data_out162;
  output [9:0] data_out163;
  wire [9:0] data_out163;
  output [9:0] data_out164;
  wire [9:0] data_out164;
  output [9:0] data_out165;
  wire [9:0] data_out165;
  output [9:0] data_out166;
  wire [9:0] data_out166;
  output [9:0] data_out167;
  wire [9:0] data_out167;
  output [9:0] data_out168;
  wire [9:0] data_out168;
  output [9:0] data_out169;
  wire [9:0] data_out169;
  output [9:0] data_out170;
  wire [9:0] data_out170;
  output [9:0] data_out171;
  wire [9:0] data_out171;
  output [9:0] data_out172;
  wire [9:0] data_out172;
  output [9:0] data_out173;
  wire [9:0] data_out173;
  output [9:0] data_out174;
  wire [9:0] data_out174;
  output [9:0] data_out175;
  wire [9:0] data_out175;
  output [9:0] data_out176;
  wire [9:0] data_out176;
  output [9:0] data_out177;
  wire [9:0] data_out177;
  output [9:0] data_out178;
  wire [9:0] data_out178;
  output [9:0] data_out179;
  wire [9:0] data_out179;
  output [9:0] data_out180;
  wire [9:0] data_out180;
  output [9:0] data_out181;
  wire [9:0] data_out181;
  output [9:0] data_out182;
  wire [9:0] data_out182;
  output [9:0] data_out183;
  wire [9:0] data_out183;
  output [9:0] data_out184;
  wire [9:0] data_out184;
  output [9:0] data_out185;
  wire [9:0] data_out185;
  output [9:0] data_out186;
  wire [9:0] data_out186;
  output [9:0] data_out187;
  wire [9:0] data_out187;
  output [9:0] data_out188;
  wire [9:0] data_out188;
  output [9:0] data_out189;
  wire [9:0] data_out189;
  output [9:0] data_out190;
  wire [9:0] data_out190;
  output [9:0] data_out193;
  wire [9:0] data_out193;
  output [9:0] data_out194;
  wire [9:0] data_out194;
  output [9:0] data_out195;
  wire [9:0] data_out195;
  output [9:0] data_out196;
  wire [9:0] data_out196;
  output [9:0] data_out197;
  wire [9:0] data_out197;
  output [9:0] data_out198;
  wire [9:0] data_out198;
  output [9:0] data_out199;
  wire [9:0] data_out199;
  output [9:0] data_out200;
  wire [9:0] data_out200;
  output [9:0] data_out201;
  wire [9:0] data_out201;
  output [9:0] data_out202;
  wire [9:0] data_out202;
  output [9:0] data_out203;
  wire [9:0] data_out203;
  output [9:0] data_out204;
  wire [9:0] data_out204;
  output [9:0] data_out205;
  wire [9:0] data_out205;
  output [9:0] data_out206;
  wire [9:0] data_out206;
  output [9:0] data_out207;
  wire [9:0] data_out207;
  output [9:0] data_out208;
  wire [9:0] data_out208;
  output [9:0] data_out209;
  wire [9:0] data_out209;
  output [9:0] data_out210;
  wire [9:0] data_out210;
  output [9:0] data_out211;
  wire [9:0] data_out211;
  output [9:0] data_out212;
  wire [9:0] data_out212;
  output [9:0] data_out213;
  wire [9:0] data_out213;
  output [9:0] data_out214;
  wire [9:0] data_out214;
  output [9:0] data_out215;
  wire [9:0] data_out215;
  output [9:0] data_out216;
  wire [9:0] data_out216;
  output [9:0] data_out217;
  wire [9:0] data_out217;
  output [9:0] data_out218;
  wire [9:0] data_out218;
  output [9:0] data_out219;
  wire [9:0] data_out219;
  output [9:0] data_out220;
  wire [9:0] data_out220;
  output [9:0] data_out221;
  wire [9:0] data_out221;
  output [9:0] data_out222;
  wire [9:0] data_out222;
  output [9:0] data_out225;
  wire [9:0] data_out225;
  output [9:0] data_out226;
  wire [9:0] data_out226;
  output [9:0] data_out227;
  wire [9:0] data_out227;
  output [9:0] data_out228;
  wire [9:0] data_out228;
  output [9:0] data_out229;
  wire [9:0] data_out229;
  output [9:0] data_out230;
  wire [9:0] data_out230;
  output [9:0] data_out231;
  wire [9:0] data_out231;
  output [9:0] data_out232;
  wire [9:0] data_out232;
  output [9:0] data_out233;
  wire [9:0] data_out233;
  output [9:0] data_out234;
  wire [9:0] data_out234;
  output [9:0] data_out235;
  wire [9:0] data_out235;
  output [9:0] data_out236;
  wire [9:0] data_out236;
  output [9:0] data_out237;
  wire [9:0] data_out237;
  output [9:0] data_out238;
  wire [9:0] data_out238;
  output [9:0] data_out239;
  wire [9:0] data_out239;
  output [9:0] data_out240;
  wire [9:0] data_out240;
  output [9:0] data_out241;
  wire [9:0] data_out241;
  output [9:0] data_out242;
  wire [9:0] data_out242;
  output [9:0] data_out243;
  wire [9:0] data_out243;
  output [9:0] data_out244;
  wire [9:0] data_out244;
  output [9:0] data_out245;
  wire [9:0] data_out245;
  output [9:0] data_out246;
  wire [9:0] data_out246;
  output [9:0] data_out247;
  wire [9:0] data_out247;
  output [9:0] data_out248;
  wire [9:0] data_out248;
  output [9:0] data_out249;
  wire [9:0] data_out249;
  output [9:0] data_out250;
  wire [9:0] data_out250;
  output [9:0] data_out251;
  wire [9:0] data_out251;
  output [9:0] data_out252;
  wire [9:0] data_out252;
  output [9:0] data_out253;
  wire [9:0] data_out253;
  output [9:0] data_out254;
  wire [9:0] data_out254;
  output [9:0] data_out257;
  wire [9:0] data_out257;
  output [9:0] data_out258;
  wire [9:0] data_out258;
  output [9:0] data_out259;
  wire [9:0] data_out259;
  output [9:0] data_out260;
  wire [9:0] data_out260;
  output [9:0] data_out261;
  wire [9:0] data_out261;
  output [9:0] data_out262;
  wire [9:0] data_out262;
  output [9:0] data_out263;
  wire [9:0] data_out263;
  output [9:0] data_out264;
  wire [9:0] data_out264;
  output [9:0] data_out265;
  wire [9:0] data_out265;
  output [9:0] data_out266;
  wire [9:0] data_out266;
  output [9:0] data_out267;
  wire [9:0] data_out267;
  output [9:0] data_out268;
  wire [9:0] data_out268;
  output [9:0] data_out269;
  wire [9:0] data_out269;
  output [9:0] data_out270;
  wire [9:0] data_out270;
  output [9:0] data_out271;
  wire [9:0] data_out271;
  output [9:0] data_out272;
  wire [9:0] data_out272;
  output [9:0] data_out273;
  wire [9:0] data_out273;
  output [9:0] data_out274;
  wire [9:0] data_out274;
  output [9:0] data_out275;
  wire [9:0] data_out275;
  output [9:0] data_out276;
  wire [9:0] data_out276;
  output [9:0] data_out277;
  wire [9:0] data_out277;
  output [9:0] data_out278;
  wire [9:0] data_out278;
  output [9:0] data_out279;
  wire [9:0] data_out279;
  output [9:0] data_out280;
  wire [9:0] data_out280;
  output [9:0] data_out281;
  wire [9:0] data_out281;
  output [9:0] data_out282;
  wire [9:0] data_out282;
  output [9:0] data_out283;
  wire [9:0] data_out283;
  output [9:0] data_out284;
  wire [9:0] data_out284;
  output [9:0] data_out285;
  wire [9:0] data_out285;
  output [9:0] data_out286;
  wire [9:0] data_out286;
  output [9:0] data_out289;
  wire [9:0] data_out289;
  output [9:0] data_out290;
  wire [9:0] data_out290;
  output [9:0] data_out291;
  wire [9:0] data_out291;
  output [9:0] data_out292;
  wire [9:0] data_out292;
  output [9:0] data_out293;
  wire [9:0] data_out293;
  output [9:0] data_out294;
  wire [9:0] data_out294;
  output [9:0] data_out295;
  wire [9:0] data_out295;
  output [9:0] data_out296;
  wire [9:0] data_out296;
  output [9:0] data_out297;
  wire [9:0] data_out297;
  output [9:0] data_out298;
  wire [9:0] data_out298;
  output [9:0] data_out299;
  wire [9:0] data_out299;
  output [9:0] data_out300;
  wire [9:0] data_out300;
  output [9:0] data_out301;
  wire [9:0] data_out301;
  output [9:0] data_out302;
  wire [9:0] data_out302;
  output [9:0] data_out303;
  wire [9:0] data_out303;
  output [9:0] data_out304;
  wire [9:0] data_out304;
  output [9:0] data_out305;
  wire [9:0] data_out305;
  output [9:0] data_out306;
  wire [9:0] data_out306;
  output [9:0] data_out307;
  wire [9:0] data_out307;
  output [9:0] data_out308;
  wire [9:0] data_out308;
  output [9:0] data_out309;
  wire [9:0] data_out309;
  output [9:0] data_out310;
  wire [9:0] data_out310;
  output [9:0] data_out311;
  wire [9:0] data_out311;
  output [9:0] data_out312;
  wire [9:0] data_out312;
  output [9:0] data_out313;
  wire [9:0] data_out313;
  output [9:0] data_out314;
  wire [9:0] data_out314;
  output [9:0] data_out315;
  wire [9:0] data_out315;
  output [9:0] data_out316;
  wire [9:0] data_out316;
  output [9:0] data_out317;
  wire [9:0] data_out317;
  output [9:0] data_out318;
  wire [9:0] data_out318;
  output [9:0] data_out321;
  wire [9:0] data_out321;
  output [9:0] data_out322;
  wire [9:0] data_out322;
  output [9:0] data_out323;
  wire [9:0] data_out323;
  output [9:0] data_out324;
  wire [9:0] data_out324;
  output [9:0] data_out325;
  wire [9:0] data_out325;
  output [9:0] data_out326;
  wire [9:0] data_out326;
  output [9:0] data_out327;
  wire [9:0] data_out327;
  output [9:0] data_out328;
  wire [9:0] data_out328;
  output [9:0] data_out329;
  wire [9:0] data_out329;
  output [9:0] data_out330;
  wire [9:0] data_out330;
  output [9:0] data_out331;
  wire [9:0] data_out331;
  output [9:0] data_out332;
  wire [9:0] data_out332;
  output [9:0] data_out333;
  wire [9:0] data_out333;
  output [9:0] data_out334;
  wire [9:0] data_out334;
  output [9:0] data_out335;
  wire [9:0] data_out335;
  output [9:0] data_out336;
  wire [9:0] data_out336;
  output [9:0] data_out337;
  wire [9:0] data_out337;
  output [9:0] data_out338;
  wire [9:0] data_out338;
  output [9:0] data_out339;
  wire [9:0] data_out339;
  output [9:0] data_out340;
  wire [9:0] data_out340;
  output [9:0] data_out341;
  wire [9:0] data_out341;
  output [9:0] data_out342;
  wire [9:0] data_out342;
  output [9:0] data_out343;
  wire [9:0] data_out343;
  output [9:0] data_out344;
  wire [9:0] data_out344;
  output [9:0] data_out345;
  wire [9:0] data_out345;
  output [9:0] data_out346;
  wire [9:0] data_out346;
  output [9:0] data_out347;
  wire [9:0] data_out347;
  output [9:0] data_out348;
  wire [9:0] data_out348;
  output [9:0] data_out349;
  wire [9:0] data_out349;
  output [9:0] data_out350;
  wire [9:0] data_out350;
  output [9:0] data_out353;
  wire [9:0] data_out353;
  output [9:0] data_out354;
  wire [9:0] data_out354;
  output [9:0] data_out355;
  wire [9:0] data_out355;
  output [9:0] data_out356;
  wire [9:0] data_out356;
  output [9:0] data_out357;
  wire [9:0] data_out357;
  output [9:0] data_out358;
  wire [9:0] data_out358;
  output [9:0] data_out359;
  wire [9:0] data_out359;
  output [9:0] data_out360;
  wire [9:0] data_out360;
  output [9:0] data_out361;
  wire [9:0] data_out361;
  output [9:0] data_out362;
  wire [9:0] data_out362;
  output [9:0] data_out363;
  wire [9:0] data_out363;
  output [9:0] data_out364;
  wire [9:0] data_out364;
  output [9:0] data_out365;
  wire [9:0] data_out365;
  output [9:0] data_out366;
  wire [9:0] data_out366;
  output [9:0] data_out367;
  wire [9:0] data_out367;
  output [9:0] data_out368;
  wire [9:0] data_out368;
  output [9:0] data_out369;
  wire [9:0] data_out369;
  output [9:0] data_out370;
  wire [9:0] data_out370;
  output [9:0] data_out371;
  wire [9:0] data_out371;
  output [9:0] data_out372;
  wire [9:0] data_out372;
  output [9:0] data_out373;
  wire [9:0] data_out373;
  output [9:0] data_out374;
  wire [9:0] data_out374;
  output [9:0] data_out375;
  wire [9:0] data_out375;
  output [9:0] data_out376;
  wire [9:0] data_out376;
  output [9:0] data_out377;
  wire [9:0] data_out377;
  output [9:0] data_out378;
  wire [9:0] data_out378;
  output [9:0] data_out379;
  wire [9:0] data_out379;
  output [9:0] data_out380;
  wire [9:0] data_out380;
  output [9:0] data_out381;
  wire [9:0] data_out381;
  output [9:0] data_out382;
  wire [9:0] data_out382;
  output [9:0] data_out385;
  wire [9:0] data_out385;
  output [9:0] data_out386;
  wire [9:0] data_out386;
  output [9:0] data_out387;
  wire [9:0] data_out387;
  output [9:0] data_out388;
  wire [9:0] data_out388;
  output [9:0] data_out389;
  wire [9:0] data_out389;
  output [9:0] data_out390;
  wire [9:0] data_out390;
  output [9:0] data_out391;
  wire [9:0] data_out391;
  output [9:0] data_out392;
  wire [9:0] data_out392;
  output [9:0] data_out393;
  wire [9:0] data_out393;
  output [9:0] data_out394;
  wire [9:0] data_out394;
  output [9:0] data_out395;
  wire [9:0] data_out395;
  output [9:0] data_out396;
  wire [9:0] data_out396;
  output [9:0] data_out397;
  wire [9:0] data_out397;
  output [9:0] data_out398;
  wire [9:0] data_out398;
  output [9:0] data_out399;
  wire [9:0] data_out399;
  output [9:0] data_out400;
  wire [9:0] data_out400;
  output [9:0] data_out401;
  wire [9:0] data_out401;
  output [9:0] data_out402;
  wire [9:0] data_out402;
  output [9:0] data_out403;
  wire [9:0] data_out403;
  output [9:0] data_out404;
  wire [9:0] data_out404;
  output [9:0] data_out405;
  wire [9:0] data_out405;
  output [9:0] data_out406;
  wire [9:0] data_out406;
  output [9:0] data_out407;
  wire [9:0] data_out407;
  output [9:0] data_out408;
  wire [9:0] data_out408;
  output [9:0] data_out409;
  wire [9:0] data_out409;
  output [9:0] data_out410;
  wire [9:0] data_out410;
  output [9:0] data_out411;
  wire [9:0] data_out411;
  output [9:0] data_out412;
  wire [9:0] data_out412;
  output [9:0] data_out413;
  wire [9:0] data_out413;
  output [9:0] data_out414;
  wire [9:0] data_out414;
  output [9:0] data_out417;
  wire [9:0] data_out417;
  output [9:0] data_out418;
  wire [9:0] data_out418;
  output [9:0] data_out419;
  wire [9:0] data_out419;
  output [9:0] data_out420;
  wire [9:0] data_out420;
  output [9:0] data_out421;
  wire [9:0] data_out421;
  output [9:0] data_out422;
  wire [9:0] data_out422;
  output [9:0] data_out423;
  wire [9:0] data_out423;
  output [9:0] data_out424;
  wire [9:0] data_out424;
  output [9:0] data_out425;
  wire [9:0] data_out425;
  output [9:0] data_out426;
  wire [9:0] data_out426;
  output [9:0] data_out427;
  wire [9:0] data_out427;
  output [9:0] data_out428;
  wire [9:0] data_out428;
  output [9:0] data_out429;
  wire [9:0] data_out429;
  output [9:0] data_out430;
  wire [9:0] data_out430;
  output [9:0] data_out431;
  wire [9:0] data_out431;
  output [9:0] data_out432;
  wire [9:0] data_out432;
  output [9:0] data_out433;
  wire [9:0] data_out433;
  output [9:0] data_out434;
  wire [9:0] data_out434;
  output [9:0] data_out435;
  wire [9:0] data_out435;
  output [9:0] data_out436;
  wire [9:0] data_out436;
  output [9:0] data_out437;
  wire [9:0] data_out437;
  output [9:0] data_out438;
  wire [9:0] data_out438;
  output [9:0] data_out439;
  wire [9:0] data_out439;
  output [9:0] data_out440;
  wire [9:0] data_out440;
  output [9:0] data_out441;
  wire [9:0] data_out441;
  output [9:0] data_out442;
  wire [9:0] data_out442;
  output [9:0] data_out443;
  wire [9:0] data_out443;
  output [9:0] data_out444;
  wire [9:0] data_out444;
  output [9:0] data_out445;
  wire [9:0] data_out445;
  output [9:0] data_out446;
  wire [9:0] data_out446;
  output [9:0] data_out449;
  wire [9:0] data_out449;
  output [9:0] data_out450;
  wire [9:0] data_out450;
  output [9:0] data_out451;
  wire [9:0] data_out451;
  output [9:0] data_out452;
  wire [9:0] data_out452;
  output [9:0] data_out453;
  wire [9:0] data_out453;
  output [9:0] data_out454;
  wire [9:0] data_out454;
  output [9:0] data_out455;
  wire [9:0] data_out455;
  output [9:0] data_out456;
  wire [9:0] data_out456;
  output [9:0] data_out457;
  wire [9:0] data_out457;
  output [9:0] data_out458;
  wire [9:0] data_out458;
  output [9:0] data_out459;
  wire [9:0] data_out459;
  output [9:0] data_out460;
  wire [9:0] data_out460;
  output [9:0] data_out461;
  wire [9:0] data_out461;
  output [9:0] data_out462;
  wire [9:0] data_out462;
  output [9:0] data_out463;
  wire [9:0] data_out463;
  output [9:0] data_out464;
  wire [9:0] data_out464;
  output [9:0] data_out465;
  wire [9:0] data_out465;
  output [9:0] data_out466;
  wire [9:0] data_out466;
  output [9:0] data_out467;
  wire [9:0] data_out467;
  output [9:0] data_out468;
  wire [9:0] data_out468;
  output [9:0] data_out469;
  wire [9:0] data_out469;
  output [9:0] data_out470;
  wire [9:0] data_out470;
  output [9:0] data_out471;
  wire [9:0] data_out471;
  output [9:0] data_out472;
  wire [9:0] data_out472;
  output [9:0] data_out473;
  wire [9:0] data_out473;
  output [9:0] data_out474;
  wire [9:0] data_out474;
  output [9:0] data_out475;
  wire [9:0] data_out475;
  output [9:0] data_out476;
  wire [9:0] data_out476;
  output [9:0] data_out477;
  wire [9:0] data_out477;
  output [9:0] data_out478;
  wire [9:0] data_out478;
  output [9:0] data_out_index33;
  wire [9:0] data_out_index33;
  output [9:0] data_out_index34;
  wire [9:0] data_out_index34;
  output [9:0] data_out_index35;
  wire [9:0] data_out_index35;
  output [9:0] data_out_index36;
  wire [9:0] data_out_index36;
  output [9:0] data_out_index37;
  wire [9:0] data_out_index37;
  output [9:0] data_out_index38;
  wire [9:0] data_out_index38;
  output [9:0] data_out_index39;
  wire [9:0] data_out_index39;
  output [9:0] data_out_index40;
  wire [9:0] data_out_index40;
  output [9:0] data_out_index41;
  wire [9:0] data_out_index41;
  output [9:0] data_out_index42;
  wire [9:0] data_out_index42;
  output [9:0] data_out_index43;
  wire [9:0] data_out_index43;
  output [9:0] data_out_index44;
  wire [9:0] data_out_index44;
  output [9:0] data_out_index45;
  wire [9:0] data_out_index45;
  output [9:0] data_out_index46;
  wire [9:0] data_out_index46;
  output [9:0] data_out_index47;
  wire [9:0] data_out_index47;
  output [9:0] data_out_index48;
  wire [9:0] data_out_index48;
  output [9:0] data_out_index49;
  wire [9:0] data_out_index49;
  output [9:0] data_out_index50;
  wire [9:0] data_out_index50;
  output [9:0] data_out_index51;
  wire [9:0] data_out_index51;
  output [9:0] data_out_index52;
  wire [9:0] data_out_index52;
  output [9:0] data_out_index53;
  wire [9:0] data_out_index53;
  output [9:0] data_out_index54;
  wire [9:0] data_out_index54;
  output [9:0] data_out_index55;
  wire [9:0] data_out_index55;
  output [9:0] data_out_index56;
  wire [9:0] data_out_index56;
  output [9:0] data_out_index57;
  wire [9:0] data_out_index57;
  output [9:0] data_out_index58;
  wire [9:0] data_out_index58;
  output [9:0] data_out_index59;
  wire [9:0] data_out_index59;
  output [9:0] data_out_index60;
  wire [9:0] data_out_index60;
  output [9:0] data_out_index61;
  wire [9:0] data_out_index61;
  output [9:0] data_out_index62;
  wire [9:0] data_out_index62;
  output [9:0] data_out_index65;
  wire [9:0] data_out_index65;
  output [9:0] data_out_index66;
  wire [9:0] data_out_index66;
  output [9:0] data_out_index67;
  wire [9:0] data_out_index67;
  output [9:0] data_out_index68;
  wire [9:0] data_out_index68;
  output [9:0] data_out_index69;
  wire [9:0] data_out_index69;
  output [9:0] data_out_index70;
  wire [9:0] data_out_index70;
  output [9:0] data_out_index71;
  wire [9:0] data_out_index71;
  output [9:0] data_out_index72;
  wire [9:0] data_out_index72;
  output [9:0] data_out_index73;
  wire [9:0] data_out_index73;
  output [9:0] data_out_index74;
  wire [9:0] data_out_index74;
  output [9:0] data_out_index75;
  wire [9:0] data_out_index75;
  output [9:0] data_out_index76;
  wire [9:0] data_out_index76;
  output [9:0] data_out_index77;
  wire [9:0] data_out_index77;
  output [9:0] data_out_index78;
  wire [9:0] data_out_index78;
  output [9:0] data_out_index79;
  wire [9:0] data_out_index79;
  output [9:0] data_out_index80;
  wire [9:0] data_out_index80;
  output [9:0] data_out_index81;
  wire [9:0] data_out_index81;
  output [9:0] data_out_index82;
  wire [9:0] data_out_index82;
  output [9:0] data_out_index83;
  wire [9:0] data_out_index83;
  output [9:0] data_out_index84;
  wire [9:0] data_out_index84;
  output [9:0] data_out_index85;
  wire [9:0] data_out_index85;
  output [9:0] data_out_index86;
  wire [9:0] data_out_index86;
  output [9:0] data_out_index87;
  wire [9:0] data_out_index87;
  output [9:0] data_out_index88;
  wire [9:0] data_out_index88;
  output [9:0] data_out_index89;
  wire [9:0] data_out_index89;
  output [9:0] data_out_index90;
  wire [9:0] data_out_index90;
  output [9:0] data_out_index91;
  wire [9:0] data_out_index91;
  output [9:0] data_out_index92;
  wire [9:0] data_out_index92;
  output [9:0] data_out_index93;
  wire [9:0] data_out_index93;
  output [9:0] data_out_index94;
  wire [9:0] data_out_index94;
  output [9:0] data_out_index97;
  wire [9:0] data_out_index97;
  output [9:0] data_out_index98;
  wire [9:0] data_out_index98;
  output [9:0] data_out_index99;
  wire [9:0] data_out_index99;
  output [9:0] data_out_index100;
  wire [9:0] data_out_index100;
  output [9:0] data_out_index101;
  wire [9:0] data_out_index101;
  output [9:0] data_out_index102;
  wire [9:0] data_out_index102;
  output [9:0] data_out_index103;
  wire [9:0] data_out_index103;
  output [9:0] data_out_index104;
  wire [9:0] data_out_index104;
  output [9:0] data_out_index105;
  wire [9:0] data_out_index105;
  output [9:0] data_out_index106;
  wire [9:0] data_out_index106;
  output [9:0] data_out_index107;
  wire [9:0] data_out_index107;
  output [9:0] data_out_index108;
  wire [9:0] data_out_index108;
  output [9:0] data_out_index109;
  wire [9:0] data_out_index109;
  output [9:0] data_out_index110;
  wire [9:0] data_out_index110;
  output [9:0] data_out_index111;
  wire [9:0] data_out_index111;
  output [9:0] data_out_index112;
  wire [9:0] data_out_index112;
  output [9:0] data_out_index113;
  wire [9:0] data_out_index113;
  output [9:0] data_out_index114;
  wire [9:0] data_out_index114;
  output [9:0] data_out_index115;
  wire [9:0] data_out_index115;
  output [9:0] data_out_index116;
  wire [9:0] data_out_index116;
  output [9:0] data_out_index117;
  wire [9:0] data_out_index117;
  output [9:0] data_out_index118;
  wire [9:0] data_out_index118;
  output [9:0] data_out_index119;
  wire [9:0] data_out_index119;
  output [9:0] data_out_index120;
  wire [9:0] data_out_index120;
  output [9:0] data_out_index121;
  wire [9:0] data_out_index121;
  output [9:0] data_out_index122;
  wire [9:0] data_out_index122;
  output [9:0] data_out_index123;
  wire [9:0] data_out_index123;
  output [9:0] data_out_index124;
  wire [9:0] data_out_index124;
  output [9:0] data_out_index125;
  wire [9:0] data_out_index125;
  output [9:0] data_out_index126;
  wire [9:0] data_out_index126;
  output [9:0] data_out_index129;
  wire [9:0] data_out_index129;
  output [9:0] data_out_index130;
  wire [9:0] data_out_index130;
  output [9:0] data_out_index131;
  wire [9:0] data_out_index131;
  output [9:0] data_out_index132;
  wire [9:0] data_out_index132;
  output [9:0] data_out_index133;
  wire [9:0] data_out_index133;
  output [9:0] data_out_index134;
  wire [9:0] data_out_index134;
  output [9:0] data_out_index135;
  wire [9:0] data_out_index135;
  output [9:0] data_out_index136;
  wire [9:0] data_out_index136;
  output [9:0] data_out_index137;
  wire [9:0] data_out_index137;
  output [9:0] data_out_index138;
  wire [9:0] data_out_index138;
  output [9:0] data_out_index139;
  wire [9:0] data_out_index139;
  output [9:0] data_out_index140;
  wire [9:0] data_out_index140;
  output [9:0] data_out_index141;
  wire [9:0] data_out_index141;
  output [9:0] data_out_index142;
  wire [9:0] data_out_index142;
  output [9:0] data_out_index143;
  wire [9:0] data_out_index143;
  output [9:0] data_out_index144;
  wire [9:0] data_out_index144;
  output [9:0] data_out_index145;
  wire [9:0] data_out_index145;
  output [9:0] data_out_index146;
  wire [9:0] data_out_index146;
  output [9:0] data_out_index147;
  wire [9:0] data_out_index147;
  output [9:0] data_out_index148;
  wire [9:0] data_out_index148;
  output [9:0] data_out_index149;
  wire [9:0] data_out_index149;
  output [9:0] data_out_index150;
  wire [9:0] data_out_index150;
  output [9:0] data_out_index151;
  wire [9:0] data_out_index151;
  output [9:0] data_out_index152;
  wire [9:0] data_out_index152;
  output [9:0] data_out_index153;
  wire [9:0] data_out_index153;
  output [9:0] data_out_index154;
  wire [9:0] data_out_index154;
  output [9:0] data_out_index155;
  wire [9:0] data_out_index155;
  output [9:0] data_out_index156;
  wire [9:0] data_out_index156;
  output [9:0] data_out_index157;
  wire [9:0] data_out_index157;
  output [9:0] data_out_index158;
  wire [9:0] data_out_index158;
  output [9:0] data_out_index161;
  wire [9:0] data_out_index161;
  output [9:0] data_out_index162;
  wire [9:0] data_out_index162;
  output [9:0] data_out_index163;
  wire [9:0] data_out_index163;
  output [9:0] data_out_index164;
  wire [9:0] data_out_index164;
  output [9:0] data_out_index165;
  wire [9:0] data_out_index165;
  output [9:0] data_out_index166;
  wire [9:0] data_out_index166;
  output [9:0] data_out_index167;
  wire [9:0] data_out_index167;
  output [9:0] data_out_index168;
  wire [9:0] data_out_index168;
  output [9:0] data_out_index169;
  wire [9:0] data_out_index169;
  output [9:0] data_out_index170;
  wire [9:0] data_out_index170;
  output [9:0] data_out_index171;
  wire [9:0] data_out_index171;
  output [9:0] data_out_index172;
  wire [9:0] data_out_index172;
  output [9:0] data_out_index173;
  wire [9:0] data_out_index173;
  output [9:0] data_out_index174;
  wire [9:0] data_out_index174;
  output [9:0] data_out_index175;
  wire [9:0] data_out_index175;
  output [9:0] data_out_index176;
  wire [9:0] data_out_index176;
  output [9:0] data_out_index177;
  wire [9:0] data_out_index177;
  output [9:0] data_out_index178;
  wire [9:0] data_out_index178;
  output [9:0] data_out_index179;
  wire [9:0] data_out_index179;
  output [9:0] data_out_index180;
  wire [9:0] data_out_index180;
  output [9:0] data_out_index181;
  wire [9:0] data_out_index181;
  output [9:0] data_out_index182;
  wire [9:0] data_out_index182;
  output [9:0] data_out_index183;
  wire [9:0] data_out_index183;
  output [9:0] data_out_index184;
  wire [9:0] data_out_index184;
  output [9:0] data_out_index185;
  wire [9:0] data_out_index185;
  output [9:0] data_out_index186;
  wire [9:0] data_out_index186;
  output [9:0] data_out_index187;
  wire [9:0] data_out_index187;
  output [9:0] data_out_index188;
  wire [9:0] data_out_index188;
  output [9:0] data_out_index189;
  wire [9:0] data_out_index189;
  output [9:0] data_out_index190;
  wire [9:0] data_out_index190;
  output [9:0] data_out_index193;
  wire [9:0] data_out_index193;
  output [9:0] data_out_index194;
  wire [9:0] data_out_index194;
  output [9:0] data_out_index195;
  wire [9:0] data_out_index195;
  output [9:0] data_out_index196;
  wire [9:0] data_out_index196;
  output [9:0] data_out_index197;
  wire [9:0] data_out_index197;
  output [9:0] data_out_index198;
  wire [9:0] data_out_index198;
  output [9:0] data_out_index199;
  wire [9:0] data_out_index199;
  output [9:0] data_out_index200;
  wire [9:0] data_out_index200;
  output [9:0] data_out_index201;
  wire [9:0] data_out_index201;
  output [9:0] data_out_index202;
  wire [9:0] data_out_index202;
  output [9:0] data_out_index203;
  wire [9:0] data_out_index203;
  output [9:0] data_out_index204;
  wire [9:0] data_out_index204;
  output [9:0] data_out_index205;
  wire [9:0] data_out_index205;
  output [9:0] data_out_index206;
  wire [9:0] data_out_index206;
  output [9:0] data_out_index207;
  wire [9:0] data_out_index207;
  output [9:0] data_out_index208;
  wire [9:0] data_out_index208;
  output [9:0] data_out_index209;
  wire [9:0] data_out_index209;
  output [9:0] data_out_index210;
  wire [9:0] data_out_index210;
  output [9:0] data_out_index211;
  wire [9:0] data_out_index211;
  output [9:0] data_out_index212;
  wire [9:0] data_out_index212;
  output [9:0] data_out_index213;
  wire [9:0] data_out_index213;
  output [9:0] data_out_index214;
  wire [9:0] data_out_index214;
  output [9:0] data_out_index215;
  wire [9:0] data_out_index215;
  output [9:0] data_out_index216;
  wire [9:0] data_out_index216;
  output [9:0] data_out_index217;
  wire [9:0] data_out_index217;
  output [9:0] data_out_index218;
  wire [9:0] data_out_index218;
  output [9:0] data_out_index219;
  wire [9:0] data_out_index219;
  output [9:0] data_out_index220;
  wire [9:0] data_out_index220;
  output [9:0] data_out_index221;
  wire [9:0] data_out_index221;
  output [9:0] data_out_index222;
  wire [9:0] data_out_index222;
  output [9:0] data_out_index225;
  wire [9:0] data_out_index225;
  output [9:0] data_out_index226;
  wire [9:0] data_out_index226;
  output [9:0] data_out_index227;
  wire [9:0] data_out_index227;
  output [9:0] data_out_index228;
  wire [9:0] data_out_index228;
  output [9:0] data_out_index229;
  wire [9:0] data_out_index229;
  output [9:0] data_out_index230;
  wire [9:0] data_out_index230;
  output [9:0] data_out_index231;
  wire [9:0] data_out_index231;
  output [9:0] data_out_index232;
  wire [9:0] data_out_index232;
  output [9:0] data_out_index233;
  wire [9:0] data_out_index233;
  output [9:0] data_out_index234;
  wire [9:0] data_out_index234;
  output [9:0] data_out_index235;
  wire [9:0] data_out_index235;
  output [9:0] data_out_index236;
  wire [9:0] data_out_index236;
  output [9:0] data_out_index237;
  wire [9:0] data_out_index237;
  output [9:0] data_out_index238;
  wire [9:0] data_out_index238;
  output [9:0] data_out_index239;
  wire [9:0] data_out_index239;
  output [9:0] data_out_index240;
  wire [9:0] data_out_index240;
  output [9:0] data_out_index241;
  wire [9:0] data_out_index241;
  output [9:0] data_out_index242;
  wire [9:0] data_out_index242;
  output [9:0] data_out_index243;
  wire [9:0] data_out_index243;
  output [9:0] data_out_index244;
  wire [9:0] data_out_index244;
  output [9:0] data_out_index245;
  wire [9:0] data_out_index245;
  output [9:0] data_out_index246;
  wire [9:0] data_out_index246;
  output [9:0] data_out_index247;
  wire [9:0] data_out_index247;
  output [9:0] data_out_index248;
  wire [9:0] data_out_index248;
  output [9:0] data_out_index249;
  wire [9:0] data_out_index249;
  output [9:0] data_out_index250;
  wire [9:0] data_out_index250;
  output [9:0] data_out_index251;
  wire [9:0] data_out_index251;
  output [9:0] data_out_index252;
  wire [9:0] data_out_index252;
  output [9:0] data_out_index253;
  wire [9:0] data_out_index253;
  output [9:0] data_out_index254;
  wire [9:0] data_out_index254;
  output [9:0] data_out_index257;
  wire [9:0] data_out_index257;
  output [9:0] data_out_index258;
  wire [9:0] data_out_index258;
  output [9:0] data_out_index259;
  wire [9:0] data_out_index259;
  output [9:0] data_out_index260;
  wire [9:0] data_out_index260;
  output [9:0] data_out_index261;
  wire [9:0] data_out_index261;
  output [9:0] data_out_index262;
  wire [9:0] data_out_index262;
  output [9:0] data_out_index263;
  wire [9:0] data_out_index263;
  output [9:0] data_out_index264;
  wire [9:0] data_out_index264;
  output [9:0] data_out_index265;
  wire [9:0] data_out_index265;
  output [9:0] data_out_index266;
  wire [9:0] data_out_index266;
  output [9:0] data_out_index267;
  wire [9:0] data_out_index267;
  output [9:0] data_out_index268;
  wire [9:0] data_out_index268;
  output [9:0] data_out_index269;
  wire [9:0] data_out_index269;
  output [9:0] data_out_index270;
  wire [9:0] data_out_index270;
  output [9:0] data_out_index271;
  wire [9:0] data_out_index271;
  output [9:0] data_out_index272;
  wire [9:0] data_out_index272;
  output [9:0] data_out_index273;
  wire [9:0] data_out_index273;
  output [9:0] data_out_index274;
  wire [9:0] data_out_index274;
  output [9:0] data_out_index275;
  wire [9:0] data_out_index275;
  output [9:0] data_out_index276;
  wire [9:0] data_out_index276;
  output [9:0] data_out_index277;
  wire [9:0] data_out_index277;
  output [9:0] data_out_index278;
  wire [9:0] data_out_index278;
  output [9:0] data_out_index279;
  wire [9:0] data_out_index279;
  output [9:0] data_out_index280;
  wire [9:0] data_out_index280;
  output [9:0] data_out_index281;
  wire [9:0] data_out_index281;
  output [9:0] data_out_index282;
  wire [9:0] data_out_index282;
  output [9:0] data_out_index283;
  wire [9:0] data_out_index283;
  output [9:0] data_out_index284;
  wire [9:0] data_out_index284;
  output [9:0] data_out_index285;
  wire [9:0] data_out_index285;
  output [9:0] data_out_index286;
  wire [9:0] data_out_index286;
  output [9:0] data_out_index289;
  wire [9:0] data_out_index289;
  output [9:0] data_out_index290;
  wire [9:0] data_out_index290;
  output [9:0] data_out_index291;
  wire [9:0] data_out_index291;
  output [9:0] data_out_index292;
  wire [9:0] data_out_index292;
  output [9:0] data_out_index293;
  wire [9:0] data_out_index293;
  output [9:0] data_out_index294;
  wire [9:0] data_out_index294;
  output [9:0] data_out_index295;
  wire [9:0] data_out_index295;
  output [9:0] data_out_index296;
  wire [9:0] data_out_index296;
  output [9:0] data_out_index297;
  wire [9:0] data_out_index297;
  output [9:0] data_out_index298;
  wire [9:0] data_out_index298;
  output [9:0] data_out_index299;
  wire [9:0] data_out_index299;
  output [9:0] data_out_index300;
  wire [9:0] data_out_index300;
  output [9:0] data_out_index301;
  wire [9:0] data_out_index301;
  output [9:0] data_out_index302;
  wire [9:0] data_out_index302;
  output [9:0] data_out_index303;
  wire [9:0] data_out_index303;
  output [9:0] data_out_index304;
  wire [9:0] data_out_index304;
  output [9:0] data_out_index305;
  wire [9:0] data_out_index305;
  output [9:0] data_out_index306;
  wire [9:0] data_out_index306;
  output [9:0] data_out_index307;
  wire [9:0] data_out_index307;
  output [9:0] data_out_index308;
  wire [9:0] data_out_index308;
  output [9:0] data_out_index309;
  wire [9:0] data_out_index309;
  output [9:0] data_out_index310;
  wire [9:0] data_out_index310;
  output [9:0] data_out_index311;
  wire [9:0] data_out_index311;
  output [9:0] data_out_index312;
  wire [9:0] data_out_index312;
  output [9:0] data_out_index313;
  wire [9:0] data_out_index313;
  output [9:0] data_out_index314;
  wire [9:0] data_out_index314;
  output [9:0] data_out_index315;
  wire [9:0] data_out_index315;
  output [9:0] data_out_index316;
  wire [9:0] data_out_index316;
  output [9:0] data_out_index317;
  wire [9:0] data_out_index317;
  output [9:0] data_out_index318;
  wire [9:0] data_out_index318;
  output [9:0] data_out_index321;
  wire [9:0] data_out_index321;
  output [9:0] data_out_index322;
  wire [9:0] data_out_index322;
  output [9:0] data_out_index323;
  wire [9:0] data_out_index323;
  output [9:0] data_out_index324;
  wire [9:0] data_out_index324;
  output [9:0] data_out_index325;
  wire [9:0] data_out_index325;
  output [9:0] data_out_index326;
  wire [9:0] data_out_index326;
  output [9:0] data_out_index327;
  wire [9:0] data_out_index327;
  output [9:0] data_out_index328;
  wire [9:0] data_out_index328;
  output [9:0] data_out_index329;
  wire [9:0] data_out_index329;
  output [9:0] data_out_index330;
  wire [9:0] data_out_index330;
  output [9:0] data_out_index331;
  wire [9:0] data_out_index331;
  output [9:0] data_out_index332;
  wire [9:0] data_out_index332;
  output [9:0] data_out_index333;
  wire [9:0] data_out_index333;
  output [9:0] data_out_index334;
  wire [9:0] data_out_index334;
  output [9:0] data_out_index335;
  wire [9:0] data_out_index335;
  output [9:0] data_out_index336;
  wire [9:0] data_out_index336;
  output [9:0] data_out_index337;
  wire [9:0] data_out_index337;
  output [9:0] data_out_index338;
  wire [9:0] data_out_index338;
  output [9:0] data_out_index339;
  wire [9:0] data_out_index339;
  output [9:0] data_out_index340;
  wire [9:0] data_out_index340;
  output [9:0] data_out_index341;
  wire [9:0] data_out_index341;
  output [9:0] data_out_index342;
  wire [9:0] data_out_index342;
  output [9:0] data_out_index343;
  wire [9:0] data_out_index343;
  output [9:0] data_out_index344;
  wire [9:0] data_out_index344;
  output [9:0] data_out_index345;
  wire [9:0] data_out_index345;
  output [9:0] data_out_index346;
  wire [9:0] data_out_index346;
  output [9:0] data_out_index347;
  wire [9:0] data_out_index347;
  output [9:0] data_out_index348;
  wire [9:0] data_out_index348;
  output [9:0] data_out_index349;
  wire [9:0] data_out_index349;
  output [9:0] data_out_index350;
  wire [9:0] data_out_index350;
  output [9:0] data_out_index353;
  wire [9:0] data_out_index353;
  output [9:0] data_out_index354;
  wire [9:0] data_out_index354;
  output [9:0] data_out_index355;
  wire [9:0] data_out_index355;
  output [9:0] data_out_index356;
  wire [9:0] data_out_index356;
  output [9:0] data_out_index357;
  wire [9:0] data_out_index357;
  output [9:0] data_out_index358;
  wire [9:0] data_out_index358;
  output [9:0] data_out_index359;
  wire [9:0] data_out_index359;
  output [9:0] data_out_index360;
  wire [9:0] data_out_index360;
  output [9:0] data_out_index361;
  wire [9:0] data_out_index361;
  output [9:0] data_out_index362;
  wire [9:0] data_out_index362;
  output [9:0] data_out_index363;
  wire [9:0] data_out_index363;
  output [9:0] data_out_index364;
  wire [9:0] data_out_index364;
  output [9:0] data_out_index365;
  wire [9:0] data_out_index365;
  output [9:0] data_out_index366;
  wire [9:0] data_out_index366;
  output [9:0] data_out_index367;
  wire [9:0] data_out_index367;
  output [9:0] data_out_index368;
  wire [9:0] data_out_index368;
  output [9:0] data_out_index369;
  wire [9:0] data_out_index369;
  output [9:0] data_out_index370;
  wire [9:0] data_out_index370;
  output [9:0] data_out_index371;
  wire [9:0] data_out_index371;
  output [9:0] data_out_index372;
  wire [9:0] data_out_index372;
  output [9:0] data_out_index373;
  wire [9:0] data_out_index373;
  output [9:0] data_out_index374;
  wire [9:0] data_out_index374;
  output [9:0] data_out_index375;
  wire [9:0] data_out_index375;
  output [9:0] data_out_index376;
  wire [9:0] data_out_index376;
  output [9:0] data_out_index377;
  wire [9:0] data_out_index377;
  output [9:0] data_out_index378;
  wire [9:0] data_out_index378;
  output [9:0] data_out_index379;
  wire [9:0] data_out_index379;
  output [9:0] data_out_index380;
  wire [9:0] data_out_index380;
  output [9:0] data_out_index381;
  wire [9:0] data_out_index381;
  output [9:0] data_out_index382;
  wire [9:0] data_out_index382;
  output [9:0] data_out_index385;
  wire [9:0] data_out_index385;
  output [9:0] data_out_index386;
  wire [9:0] data_out_index386;
  output [9:0] data_out_index387;
  wire [9:0] data_out_index387;
  output [9:0] data_out_index388;
  wire [9:0] data_out_index388;
  output [9:0] data_out_index389;
  wire [9:0] data_out_index389;
  output [9:0] data_out_index390;
  wire [9:0] data_out_index390;
  output [9:0] data_out_index391;
  wire [9:0] data_out_index391;
  output [9:0] data_out_index392;
  wire [9:0] data_out_index392;
  output [9:0] data_out_index393;
  wire [9:0] data_out_index393;
  output [9:0] data_out_index394;
  wire [9:0] data_out_index394;
  output [9:0] data_out_index395;
  wire [9:0] data_out_index395;
  output [9:0] data_out_index396;
  wire [9:0] data_out_index396;
  output [9:0] data_out_index397;
  wire [9:0] data_out_index397;
  output [9:0] data_out_index398;
  wire [9:0] data_out_index398;
  output [9:0] data_out_index399;
  wire [9:0] data_out_index399;
  output [9:0] data_out_index400;
  wire [9:0] data_out_index400;
  output [9:0] data_out_index401;
  wire [9:0] data_out_index401;
  output [9:0] data_out_index402;
  wire [9:0] data_out_index402;
  output [9:0] data_out_index403;
  wire [9:0] data_out_index403;
  output [9:0] data_out_index404;
  wire [9:0] data_out_index404;
  output [9:0] data_out_index405;
  wire [9:0] data_out_index405;
  output [9:0] data_out_index406;
  wire [9:0] data_out_index406;
  output [9:0] data_out_index407;
  wire [9:0] data_out_index407;
  output [9:0] data_out_index408;
  wire [9:0] data_out_index408;
  output [9:0] data_out_index409;
  wire [9:0] data_out_index409;
  output [9:0] data_out_index410;
  wire [9:0] data_out_index410;
  output [9:0] data_out_index411;
  wire [9:0] data_out_index411;
  output [9:0] data_out_index412;
  wire [9:0] data_out_index412;
  output [9:0] data_out_index413;
  wire [9:0] data_out_index413;
  output [9:0] data_out_index414;
  wire [9:0] data_out_index414;
  output [9:0] data_out_index417;
  wire [9:0] data_out_index417;
  output [9:0] data_out_index418;
  wire [9:0] data_out_index418;
  output [9:0] data_out_index419;
  wire [9:0] data_out_index419;
  output [9:0] data_out_index420;
  wire [9:0] data_out_index420;
  output [9:0] data_out_index421;
  wire [9:0] data_out_index421;
  output [9:0] data_out_index422;
  wire [9:0] data_out_index422;
  output [9:0] data_out_index423;
  wire [9:0] data_out_index423;
  output [9:0] data_out_index424;
  wire [9:0] data_out_index424;
  output [9:0] data_out_index425;
  wire [9:0] data_out_index425;
  output [9:0] data_out_index426;
  wire [9:0] data_out_index426;
  output [9:0] data_out_index427;
  wire [9:0] data_out_index427;
  output [9:0] data_out_index428;
  wire [9:0] data_out_index428;
  output [9:0] data_out_index429;
  wire [9:0] data_out_index429;
  output [9:0] data_out_index430;
  wire [9:0] data_out_index430;
  output [9:0] data_out_index431;
  wire [9:0] data_out_index431;
  output [9:0] data_out_index432;
  wire [9:0] data_out_index432;
  output [9:0] data_out_index433;
  wire [9:0] data_out_index433;
  output [9:0] data_out_index434;
  wire [9:0] data_out_index434;
  output [9:0] data_out_index435;
  wire [9:0] data_out_index435;
  output [9:0] data_out_index436;
  wire [9:0] data_out_index436;
  output [9:0] data_out_index437;
  wire [9:0] data_out_index437;
  output [9:0] data_out_index438;
  wire [9:0] data_out_index438;
  output [9:0] data_out_index439;
  wire [9:0] data_out_index439;
  output [9:0] data_out_index440;
  wire [9:0] data_out_index440;
  output [9:0] data_out_index441;
  wire [9:0] data_out_index441;
  output [9:0] data_out_index442;
  wire [9:0] data_out_index442;
  output [9:0] data_out_index443;
  wire [9:0] data_out_index443;
  output [9:0] data_out_index444;
  wire [9:0] data_out_index444;
  output [9:0] data_out_index445;
  wire [9:0] data_out_index445;
  output [9:0] data_out_index446;
  wire [9:0] data_out_index446;
  output [9:0] data_out_index449;
  wire [9:0] data_out_index449;
  output [9:0] data_out_index450;
  wire [9:0] data_out_index450;
  output [9:0] data_out_index451;
  wire [9:0] data_out_index451;
  output [9:0] data_out_index452;
  wire [9:0] data_out_index452;
  output [9:0] data_out_index453;
  wire [9:0] data_out_index453;
  output [9:0] data_out_index454;
  wire [9:0] data_out_index454;
  output [9:0] data_out_index455;
  wire [9:0] data_out_index455;
  output [9:0] data_out_index456;
  wire [9:0] data_out_index456;
  output [9:0] data_out_index457;
  wire [9:0] data_out_index457;
  output [9:0] data_out_index458;
  wire [9:0] data_out_index458;
  output [9:0] data_out_index459;
  wire [9:0] data_out_index459;
  output [9:0] data_out_index460;
  wire [9:0] data_out_index460;
  output [9:0] data_out_index461;
  wire [9:0] data_out_index461;
  output [9:0] data_out_index462;
  wire [9:0] data_out_index462;
  output [9:0] data_out_index463;
  wire [9:0] data_out_index463;
  output [9:0] data_out_index464;
  wire [9:0] data_out_index464;
  output [9:0] data_out_index465;
  wire [9:0] data_out_index465;
  output [9:0] data_out_index466;
  wire [9:0] data_out_index466;
  output [9:0] data_out_index467;
  wire [9:0] data_out_index467;
  output [9:0] data_out_index468;
  wire [9:0] data_out_index468;
  output [9:0] data_out_index469;
  wire [9:0] data_out_index469;
  output [9:0] data_out_index470;
  wire [9:0] data_out_index470;
  output [9:0] data_out_index471;
  wire [9:0] data_out_index471;
  output [9:0] data_out_index472;
  wire [9:0] data_out_index472;
  output [9:0] data_out_index473;
  wire [9:0] data_out_index473;
  output [9:0] data_out_index474;
  wire [9:0] data_out_index474;
  output [9:0] data_out_index475;
  wire [9:0] data_out_index475;
  output [9:0] data_out_index476;
  wire [9:0] data_out_index476;
  output [9:0] data_out_index477;
  wire [9:0] data_out_index477;
  output [9:0] data_out_index478;
  wire [9:0] data_out_index478;
  input [1:0] sg_in33;
  wire [1:0] sg_in33;
  input [1:0] sg_in34;
  wire [1:0] sg_in34;
  input [1:0] sg_in35;
  wire [1:0] sg_in35;
  input [1:0] sg_in36;
  wire [1:0] sg_in36;
  input [1:0] sg_in37;
  wire [1:0] sg_in37;
  input [1:0] sg_in38;
  wire [1:0] sg_in38;
  input [1:0] sg_in39;
  wire [1:0] sg_in39;
  input [1:0] sg_in40;
  wire [1:0] sg_in40;
  input [1:0] sg_in41;
  wire [1:0] sg_in41;
  input [1:0] sg_in42;
  wire [1:0] sg_in42;
  input [1:0] sg_in43;
  wire [1:0] sg_in43;
  input [1:0] sg_in44;
  wire [1:0] sg_in44;
  input [1:0] sg_in45;
  wire [1:0] sg_in45;
  input [1:0] sg_in46;
  wire [1:0] sg_in46;
  input [1:0] sg_in47;
  wire [1:0] sg_in47;
  input [1:0] sg_in48;
  wire [1:0] sg_in48;
  input [1:0] sg_in49;
  wire [1:0] sg_in49;
  input [1:0] sg_in50;
  wire [1:0] sg_in50;
  input [1:0] sg_in51;
  wire [1:0] sg_in51;
  input [1:0] sg_in52;
  wire [1:0] sg_in52;
  input [1:0] sg_in53;
  wire [1:0] sg_in53;
  input [1:0] sg_in54;
  wire [1:0] sg_in54;
  input [1:0] sg_in55;
  wire [1:0] sg_in55;
  input [1:0] sg_in56;
  wire [1:0] sg_in56;
  input [1:0] sg_in57;
  wire [1:0] sg_in57;
  input [1:0] sg_in58;
  wire [1:0] sg_in58;
  input [1:0] sg_in59;
  wire [1:0] sg_in59;
  input [1:0] sg_in60;
  wire [1:0] sg_in60;
  input [1:0] sg_in61;
  wire [1:0] sg_in61;
  input [1:0] sg_in62;
  wire [1:0] sg_in62;
  input [1:0] sg_in65;
  wire [1:0] sg_in65;
  input [1:0] sg_in66;
  wire [1:0] sg_in66;
  input [1:0] sg_in67;
  wire [1:0] sg_in67;
  input [1:0] sg_in68;
  wire [1:0] sg_in68;
  input [1:0] sg_in69;
  wire [1:0] sg_in69;
  input [1:0] sg_in70;
  wire [1:0] sg_in70;
  input [1:0] sg_in71;
  wire [1:0] sg_in71;
  input [1:0] sg_in72;
  wire [1:0] sg_in72;
  input [1:0] sg_in73;
  wire [1:0] sg_in73;
  input [1:0] sg_in74;
  wire [1:0] sg_in74;
  input [1:0] sg_in75;
  wire [1:0] sg_in75;
  input [1:0] sg_in76;
  wire [1:0] sg_in76;
  input [1:0] sg_in77;
  wire [1:0] sg_in77;
  input [1:0] sg_in78;
  wire [1:0] sg_in78;
  input [1:0] sg_in79;
  wire [1:0] sg_in79;
  input [1:0] sg_in80;
  wire [1:0] sg_in80;
  input [1:0] sg_in81;
  wire [1:0] sg_in81;
  input [1:0] sg_in82;
  wire [1:0] sg_in82;
  input [1:0] sg_in83;
  wire [1:0] sg_in83;
  input [1:0] sg_in84;
  wire [1:0] sg_in84;
  input [1:0] sg_in85;
  wire [1:0] sg_in85;
  input [1:0] sg_in86;
  wire [1:0] sg_in86;
  input [1:0] sg_in87;
  wire [1:0] sg_in87;
  input [1:0] sg_in88;
  wire [1:0] sg_in88;
  input [1:0] sg_in89;
  wire [1:0] sg_in89;
  input [1:0] sg_in90;
  wire [1:0] sg_in90;
  input [1:0] sg_in91;
  wire [1:0] sg_in91;
  input [1:0] sg_in92;
  wire [1:0] sg_in92;
  input [1:0] sg_in93;
  wire [1:0] sg_in93;
  input [1:0] sg_in94;
  wire [1:0] sg_in94;
  input [1:0] sg_in97;
  wire [1:0] sg_in97;
  input [1:0] sg_in98;
  wire [1:0] sg_in98;
  input [1:0] sg_in99;
  wire [1:0] sg_in99;
  input [1:0] sg_in100;
  wire [1:0] sg_in100;
  input [1:0] sg_in101;
  wire [1:0] sg_in101;
  input [1:0] sg_in102;
  wire [1:0] sg_in102;
  input [1:0] sg_in103;
  wire [1:0] sg_in103;
  input [1:0] sg_in104;
  wire [1:0] sg_in104;
  input [1:0] sg_in105;
  wire [1:0] sg_in105;
  input [1:0] sg_in106;
  wire [1:0] sg_in106;
  input [1:0] sg_in107;
  wire [1:0] sg_in107;
  input [1:0] sg_in108;
  wire [1:0] sg_in108;
  input [1:0] sg_in109;
  wire [1:0] sg_in109;
  input [1:0] sg_in110;
  wire [1:0] sg_in110;
  input [1:0] sg_in111;
  wire [1:0] sg_in111;
  input [1:0] sg_in112;
  wire [1:0] sg_in112;
  input [1:0] sg_in113;
  wire [1:0] sg_in113;
  input [1:0] sg_in114;
  wire [1:0] sg_in114;
  input [1:0] sg_in115;
  wire [1:0] sg_in115;
  input [1:0] sg_in116;
  wire [1:0] sg_in116;
  input [1:0] sg_in117;
  wire [1:0] sg_in117;
  input [1:0] sg_in118;
  wire [1:0] sg_in118;
  input [1:0] sg_in119;
  wire [1:0] sg_in119;
  input [1:0] sg_in120;
  wire [1:0] sg_in120;
  input [1:0] sg_in121;
  wire [1:0] sg_in121;
  input [1:0] sg_in122;
  wire [1:0] sg_in122;
  input [1:0] sg_in123;
  wire [1:0] sg_in123;
  input [1:0] sg_in124;
  wire [1:0] sg_in124;
  input [1:0] sg_in125;
  wire [1:0] sg_in125;
  input [1:0] sg_in126;
  wire [1:0] sg_in126;
  input [1:0] sg_in129;
  wire [1:0] sg_in129;
  input [1:0] sg_in130;
  wire [1:0] sg_in130;
  input [1:0] sg_in131;
  wire [1:0] sg_in131;
  input [1:0] sg_in132;
  wire [1:0] sg_in132;
  input [1:0] sg_in133;
  wire [1:0] sg_in133;
  input [1:0] sg_in134;
  wire [1:0] sg_in134;
  input [1:0] sg_in135;
  wire [1:0] sg_in135;
  input [1:0] sg_in136;
  wire [1:0] sg_in136;
  input [1:0] sg_in137;
  wire [1:0] sg_in137;
  input [1:0] sg_in138;
  wire [1:0] sg_in138;
  input [1:0] sg_in139;
  wire [1:0] sg_in139;
  input [1:0] sg_in140;
  wire [1:0] sg_in140;
  input [1:0] sg_in141;
  wire [1:0] sg_in141;
  input [1:0] sg_in142;
  wire [1:0] sg_in142;
  input [1:0] sg_in143;
  wire [1:0] sg_in143;
  input [1:0] sg_in144;
  wire [1:0] sg_in144;
  input [1:0] sg_in145;
  wire [1:0] sg_in145;
  input [1:0] sg_in146;
  wire [1:0] sg_in146;
  input [1:0] sg_in147;
  wire [1:0] sg_in147;
  input [1:0] sg_in148;
  wire [1:0] sg_in148;
  input [1:0] sg_in149;
  wire [1:0] sg_in149;
  input [1:0] sg_in150;
  wire [1:0] sg_in150;
  input [1:0] sg_in151;
  wire [1:0] sg_in151;
  input [1:0] sg_in152;
  wire [1:0] sg_in152;
  input [1:0] sg_in153;
  wire [1:0] sg_in153;
  input [1:0] sg_in154;
  wire [1:0] sg_in154;
  input [1:0] sg_in155;
  wire [1:0] sg_in155;
  input [1:0] sg_in156;
  wire [1:0] sg_in156;
  input [1:0] sg_in157;
  wire [1:0] sg_in157;
  input [1:0] sg_in158;
  wire [1:0] sg_in158;
  input [1:0] sg_in161;
  wire [1:0] sg_in161;
  input [1:0] sg_in162;
  wire [1:0] sg_in162;
  input [1:0] sg_in163;
  wire [1:0] sg_in163;
  input [1:0] sg_in164;
  wire [1:0] sg_in164;
  input [1:0] sg_in165;
  wire [1:0] sg_in165;
  input [1:0] sg_in166;
  wire [1:0] sg_in166;
  input [1:0] sg_in167;
  wire [1:0] sg_in167;
  input [1:0] sg_in168;
  wire [1:0] sg_in168;
  input [1:0] sg_in169;
  wire [1:0] sg_in169;
  input [1:0] sg_in170;
  wire [1:0] sg_in170;
  input [1:0] sg_in171;
  wire [1:0] sg_in171;
  input [1:0] sg_in172;
  wire [1:0] sg_in172;
  input [1:0] sg_in173;
  wire [1:0] sg_in173;
  input [1:0] sg_in174;
  wire [1:0] sg_in174;
  input [1:0] sg_in175;
  wire [1:0] sg_in175;
  input [1:0] sg_in176;
  wire [1:0] sg_in176;
  input [1:0] sg_in177;
  wire [1:0] sg_in177;
  input [1:0] sg_in178;
  wire [1:0] sg_in178;
  input [1:0] sg_in179;
  wire [1:0] sg_in179;
  input [1:0] sg_in180;
  wire [1:0] sg_in180;
  input [1:0] sg_in181;
  wire [1:0] sg_in181;
  input [1:0] sg_in182;
  wire [1:0] sg_in182;
  input [1:0] sg_in183;
  wire [1:0] sg_in183;
  input [1:0] sg_in184;
  wire [1:0] sg_in184;
  input [1:0] sg_in185;
  wire [1:0] sg_in185;
  input [1:0] sg_in186;
  wire [1:0] sg_in186;
  input [1:0] sg_in187;
  wire [1:0] sg_in187;
  input [1:0] sg_in188;
  wire [1:0] sg_in188;
  input [1:0] sg_in189;
  wire [1:0] sg_in189;
  input [1:0] sg_in190;
  wire [1:0] sg_in190;
  input [1:0] sg_in193;
  wire [1:0] sg_in193;
  input [1:0] sg_in194;
  wire [1:0] sg_in194;
  input [1:0] sg_in195;
  wire [1:0] sg_in195;
  input [1:0] sg_in196;
  wire [1:0] sg_in196;
  input [1:0] sg_in197;
  wire [1:0] sg_in197;
  input [1:0] sg_in198;
  wire [1:0] sg_in198;
  input [1:0] sg_in199;
  wire [1:0] sg_in199;
  input [1:0] sg_in200;
  wire [1:0] sg_in200;
  input [1:0] sg_in201;
  wire [1:0] sg_in201;
  input [1:0] sg_in202;
  wire [1:0] sg_in202;
  input [1:0] sg_in203;
  wire [1:0] sg_in203;
  input [1:0] sg_in204;
  wire [1:0] sg_in204;
  input [1:0] sg_in205;
  wire [1:0] sg_in205;
  input [1:0] sg_in206;
  wire [1:0] sg_in206;
  input [1:0] sg_in207;
  wire [1:0] sg_in207;
  input [1:0] sg_in208;
  wire [1:0] sg_in208;
  input [1:0] sg_in209;
  wire [1:0] sg_in209;
  input [1:0] sg_in210;
  wire [1:0] sg_in210;
  input [1:0] sg_in211;
  wire [1:0] sg_in211;
  input [1:0] sg_in212;
  wire [1:0] sg_in212;
  input [1:0] sg_in213;
  wire [1:0] sg_in213;
  input [1:0] sg_in214;
  wire [1:0] sg_in214;
  input [1:0] sg_in215;
  wire [1:0] sg_in215;
  input [1:0] sg_in216;
  wire [1:0] sg_in216;
  input [1:0] sg_in217;
  wire [1:0] sg_in217;
  input [1:0] sg_in218;
  wire [1:0] sg_in218;
  input [1:0] sg_in219;
  wire [1:0] sg_in219;
  input [1:0] sg_in220;
  wire [1:0] sg_in220;
  input [1:0] sg_in221;
  wire [1:0] sg_in221;
  input [1:0] sg_in222;
  wire [1:0] sg_in222;
  input [1:0] sg_in225;
  wire [1:0] sg_in225;
  input [1:0] sg_in226;
  wire [1:0] sg_in226;
  input [1:0] sg_in227;
  wire [1:0] sg_in227;
  input [1:0] sg_in228;
  wire [1:0] sg_in228;
  input [1:0] sg_in229;
  wire [1:0] sg_in229;
  input [1:0] sg_in230;
  wire [1:0] sg_in230;
  input [1:0] sg_in231;
  wire [1:0] sg_in231;
  input [1:0] sg_in232;
  wire [1:0] sg_in232;
  input [1:0] sg_in233;
  wire [1:0] sg_in233;
  input [1:0] sg_in234;
  wire [1:0] sg_in234;
  input [1:0] sg_in235;
  wire [1:0] sg_in235;
  input [1:0] sg_in236;
  wire [1:0] sg_in236;
  input [1:0] sg_in237;
  wire [1:0] sg_in237;
  input [1:0] sg_in238;
  wire [1:0] sg_in238;
  input [1:0] sg_in239;
  wire [1:0] sg_in239;
  input [1:0] sg_in240;
  wire [1:0] sg_in240;
  input [1:0] sg_in241;
  wire [1:0] sg_in241;
  input [1:0] sg_in242;
  wire [1:0] sg_in242;
  input [1:0] sg_in243;
  wire [1:0] sg_in243;
  input [1:0] sg_in244;
  wire [1:0] sg_in244;
  input [1:0] sg_in245;
  wire [1:0] sg_in245;
  input [1:0] sg_in246;
  wire [1:0] sg_in246;
  input [1:0] sg_in247;
  wire [1:0] sg_in247;
  input [1:0] sg_in248;
  wire [1:0] sg_in248;
  input [1:0] sg_in249;
  wire [1:0] sg_in249;
  input [1:0] sg_in250;
  wire [1:0] sg_in250;
  input [1:0] sg_in251;
  wire [1:0] sg_in251;
  input [1:0] sg_in252;
  wire [1:0] sg_in252;
  input [1:0] sg_in253;
  wire [1:0] sg_in253;
  input [1:0] sg_in254;
  wire [1:0] sg_in254;
  input [1:0] sg_in257;
  wire [1:0] sg_in257;
  input [1:0] sg_in258;
  wire [1:0] sg_in258;
  input [1:0] sg_in259;
  wire [1:0] sg_in259;
  input [1:0] sg_in260;
  wire [1:0] sg_in260;
  input [1:0] sg_in261;
  wire [1:0] sg_in261;
  input [1:0] sg_in262;
  wire [1:0] sg_in262;
  input [1:0] sg_in263;
  wire [1:0] sg_in263;
  input [1:0] sg_in264;
  wire [1:0] sg_in264;
  input [1:0] sg_in265;
  wire [1:0] sg_in265;
  input [1:0] sg_in266;
  wire [1:0] sg_in266;
  input [1:0] sg_in267;
  wire [1:0] sg_in267;
  input [1:0] sg_in268;
  wire [1:0] sg_in268;
  input [1:0] sg_in269;
  wire [1:0] sg_in269;
  input [1:0] sg_in270;
  wire [1:0] sg_in270;
  input [1:0] sg_in271;
  wire [1:0] sg_in271;
  input [1:0] sg_in272;
  wire [1:0] sg_in272;
  input [1:0] sg_in273;
  wire [1:0] sg_in273;
  input [1:0] sg_in274;
  wire [1:0] sg_in274;
  input [1:0] sg_in275;
  wire [1:0] sg_in275;
  input [1:0] sg_in276;
  wire [1:0] sg_in276;
  input [1:0] sg_in277;
  wire [1:0] sg_in277;
  input [1:0] sg_in278;
  wire [1:0] sg_in278;
  input [1:0] sg_in279;
  wire [1:0] sg_in279;
  input [1:0] sg_in280;
  wire [1:0] sg_in280;
  input [1:0] sg_in281;
  wire [1:0] sg_in281;
  input [1:0] sg_in282;
  wire [1:0] sg_in282;
  input [1:0] sg_in283;
  wire [1:0] sg_in283;
  input [1:0] sg_in284;
  wire [1:0] sg_in284;
  input [1:0] sg_in285;
  wire [1:0] sg_in285;
  input [1:0] sg_in286;
  wire [1:0] sg_in286;
  input [1:0] sg_in289;
  wire [1:0] sg_in289;
  input [1:0] sg_in290;
  wire [1:0] sg_in290;
  input [1:0] sg_in291;
  wire [1:0] sg_in291;
  input [1:0] sg_in292;
  wire [1:0] sg_in292;
  input [1:0] sg_in293;
  wire [1:0] sg_in293;
  input [1:0] sg_in294;
  wire [1:0] sg_in294;
  input [1:0] sg_in295;
  wire [1:0] sg_in295;
  input [1:0] sg_in296;
  wire [1:0] sg_in296;
  input [1:0] sg_in297;
  wire [1:0] sg_in297;
  input [1:0] sg_in298;
  wire [1:0] sg_in298;
  input [1:0] sg_in299;
  wire [1:0] sg_in299;
  input [1:0] sg_in300;
  wire [1:0] sg_in300;
  input [1:0] sg_in301;
  wire [1:0] sg_in301;
  input [1:0] sg_in302;
  wire [1:0] sg_in302;
  input [1:0] sg_in303;
  wire [1:0] sg_in303;
  input [1:0] sg_in304;
  wire [1:0] sg_in304;
  input [1:0] sg_in305;
  wire [1:0] sg_in305;
  input [1:0] sg_in306;
  wire [1:0] sg_in306;
  input [1:0] sg_in307;
  wire [1:0] sg_in307;
  input [1:0] sg_in308;
  wire [1:0] sg_in308;
  input [1:0] sg_in309;
  wire [1:0] sg_in309;
  input [1:0] sg_in310;
  wire [1:0] sg_in310;
  input [1:0] sg_in311;
  wire [1:0] sg_in311;
  input [1:0] sg_in312;
  wire [1:0] sg_in312;
  input [1:0] sg_in313;
  wire [1:0] sg_in313;
  input [1:0] sg_in314;
  wire [1:0] sg_in314;
  input [1:0] sg_in315;
  wire [1:0] sg_in315;
  input [1:0] sg_in316;
  wire [1:0] sg_in316;
  input [1:0] sg_in317;
  wire [1:0] sg_in317;
  input [1:0] sg_in318;
  wire [1:0] sg_in318;
  input [1:0] sg_in321;
  wire [1:0] sg_in321;
  input [1:0] sg_in322;
  wire [1:0] sg_in322;
  input [1:0] sg_in323;
  wire [1:0] sg_in323;
  input [1:0] sg_in324;
  wire [1:0] sg_in324;
  input [1:0] sg_in325;
  wire [1:0] sg_in325;
  input [1:0] sg_in326;
  wire [1:0] sg_in326;
  input [1:0] sg_in327;
  wire [1:0] sg_in327;
  input [1:0] sg_in328;
  wire [1:0] sg_in328;
  input [1:0] sg_in329;
  wire [1:0] sg_in329;
  input [1:0] sg_in330;
  wire [1:0] sg_in330;
  input [1:0] sg_in331;
  wire [1:0] sg_in331;
  input [1:0] sg_in332;
  wire [1:0] sg_in332;
  input [1:0] sg_in333;
  wire [1:0] sg_in333;
  input [1:0] sg_in334;
  wire [1:0] sg_in334;
  input [1:0] sg_in335;
  wire [1:0] sg_in335;
  input [1:0] sg_in336;
  wire [1:0] sg_in336;
  input [1:0] sg_in337;
  wire [1:0] sg_in337;
  input [1:0] sg_in338;
  wire [1:0] sg_in338;
  input [1:0] sg_in339;
  wire [1:0] sg_in339;
  input [1:0] sg_in340;
  wire [1:0] sg_in340;
  input [1:0] sg_in341;
  wire [1:0] sg_in341;
  input [1:0] sg_in342;
  wire [1:0] sg_in342;
  input [1:0] sg_in343;
  wire [1:0] sg_in343;
  input [1:0] sg_in344;
  wire [1:0] sg_in344;
  input [1:0] sg_in345;
  wire [1:0] sg_in345;
  input [1:0] sg_in346;
  wire [1:0] sg_in346;
  input [1:0] sg_in347;
  wire [1:0] sg_in347;
  input [1:0] sg_in348;
  wire [1:0] sg_in348;
  input [1:0] sg_in349;
  wire [1:0] sg_in349;
  input [1:0] sg_in350;
  wire [1:0] sg_in350;
  input [1:0] sg_in353;
  wire [1:0] sg_in353;
  input [1:0] sg_in354;
  wire [1:0] sg_in354;
  input [1:0] sg_in355;
  wire [1:0] sg_in355;
  input [1:0] sg_in356;
  wire [1:0] sg_in356;
  input [1:0] sg_in357;
  wire [1:0] sg_in357;
  input [1:0] sg_in358;
  wire [1:0] sg_in358;
  input [1:0] sg_in359;
  wire [1:0] sg_in359;
  input [1:0] sg_in360;
  wire [1:0] sg_in360;
  input [1:0] sg_in361;
  wire [1:0] sg_in361;
  input [1:0] sg_in362;
  wire [1:0] sg_in362;
  input [1:0] sg_in363;
  wire [1:0] sg_in363;
  input [1:0] sg_in364;
  wire [1:0] sg_in364;
  input [1:0] sg_in365;
  wire [1:0] sg_in365;
  input [1:0] sg_in366;
  wire [1:0] sg_in366;
  input [1:0] sg_in367;
  wire [1:0] sg_in367;
  input [1:0] sg_in368;
  wire [1:0] sg_in368;
  input [1:0] sg_in369;
  wire [1:0] sg_in369;
  input [1:0] sg_in370;
  wire [1:0] sg_in370;
  input [1:0] sg_in371;
  wire [1:0] sg_in371;
  input [1:0] sg_in372;
  wire [1:0] sg_in372;
  input [1:0] sg_in373;
  wire [1:0] sg_in373;
  input [1:0] sg_in374;
  wire [1:0] sg_in374;
  input [1:0] sg_in375;
  wire [1:0] sg_in375;
  input [1:0] sg_in376;
  wire [1:0] sg_in376;
  input [1:0] sg_in377;
  wire [1:0] sg_in377;
  input [1:0] sg_in378;
  wire [1:0] sg_in378;
  input [1:0] sg_in379;
  wire [1:0] sg_in379;
  input [1:0] sg_in380;
  wire [1:0] sg_in380;
  input [1:0] sg_in381;
  wire [1:0] sg_in381;
  input [1:0] sg_in382;
  wire [1:0] sg_in382;
  input [1:0] sg_in385;
  wire [1:0] sg_in385;
  input [1:0] sg_in386;
  wire [1:0] sg_in386;
  input [1:0] sg_in387;
  wire [1:0] sg_in387;
  input [1:0] sg_in388;
  wire [1:0] sg_in388;
  input [1:0] sg_in389;
  wire [1:0] sg_in389;
  input [1:0] sg_in390;
  wire [1:0] sg_in390;
  input [1:0] sg_in391;
  wire [1:0] sg_in391;
  input [1:0] sg_in392;
  wire [1:0] sg_in392;
  input [1:0] sg_in393;
  wire [1:0] sg_in393;
  input [1:0] sg_in394;
  wire [1:0] sg_in394;
  input [1:0] sg_in395;
  wire [1:0] sg_in395;
  input [1:0] sg_in396;
  wire [1:0] sg_in396;
  input [1:0] sg_in397;
  wire [1:0] sg_in397;
  input [1:0] sg_in398;
  wire [1:0] sg_in398;
  input [1:0] sg_in399;
  wire [1:0] sg_in399;
  input [1:0] sg_in400;
  wire [1:0] sg_in400;
  input [1:0] sg_in401;
  wire [1:0] sg_in401;
  input [1:0] sg_in402;
  wire [1:0] sg_in402;
  input [1:0] sg_in403;
  wire [1:0] sg_in403;
  input [1:0] sg_in404;
  wire [1:0] sg_in404;
  input [1:0] sg_in405;
  wire [1:0] sg_in405;
  input [1:0] sg_in406;
  wire [1:0] sg_in406;
  input [1:0] sg_in407;
  wire [1:0] sg_in407;
  input [1:0] sg_in408;
  wire [1:0] sg_in408;
  input [1:0] sg_in409;
  wire [1:0] sg_in409;
  input [1:0] sg_in410;
  wire [1:0] sg_in410;
  input [1:0] sg_in411;
  wire [1:0] sg_in411;
  input [1:0] sg_in412;
  wire [1:0] sg_in412;
  input [1:0] sg_in413;
  wire [1:0] sg_in413;
  input [1:0] sg_in414;
  wire [1:0] sg_in414;
  input [1:0] sg_in417;
  wire [1:0] sg_in417;
  input [1:0] sg_in418;
  wire [1:0] sg_in418;
  input [1:0] sg_in419;
  wire [1:0] sg_in419;
  input [1:0] sg_in420;
  wire [1:0] sg_in420;
  input [1:0] sg_in421;
  wire [1:0] sg_in421;
  input [1:0] sg_in422;
  wire [1:0] sg_in422;
  input [1:0] sg_in423;
  wire [1:0] sg_in423;
  input [1:0] sg_in424;
  wire [1:0] sg_in424;
  input [1:0] sg_in425;
  wire [1:0] sg_in425;
  input [1:0] sg_in426;
  wire [1:0] sg_in426;
  input [1:0] sg_in427;
  wire [1:0] sg_in427;
  input [1:0] sg_in428;
  wire [1:0] sg_in428;
  input [1:0] sg_in429;
  wire [1:0] sg_in429;
  input [1:0] sg_in430;
  wire [1:0] sg_in430;
  input [1:0] sg_in431;
  wire [1:0] sg_in431;
  input [1:0] sg_in432;
  wire [1:0] sg_in432;
  input [1:0] sg_in433;
  wire [1:0] sg_in433;
  input [1:0] sg_in434;
  wire [1:0] sg_in434;
  input [1:0] sg_in435;
  wire [1:0] sg_in435;
  input [1:0] sg_in436;
  wire [1:0] sg_in436;
  input [1:0] sg_in437;
  wire [1:0] sg_in437;
  input [1:0] sg_in438;
  wire [1:0] sg_in438;
  input [1:0] sg_in439;
  wire [1:0] sg_in439;
  input [1:0] sg_in440;
  wire [1:0] sg_in440;
  input [1:0] sg_in441;
  wire [1:0] sg_in441;
  input [1:0] sg_in442;
  wire [1:0] sg_in442;
  input [1:0] sg_in443;
  wire [1:0] sg_in443;
  input [1:0] sg_in444;
  wire [1:0] sg_in444;
  input [1:0] sg_in445;
  wire [1:0] sg_in445;
  input [1:0] sg_in446;
  wire [1:0] sg_in446;
  input [1:0] sg_in449;
  wire [1:0] sg_in449;
  input [1:0] sg_in450;
  wire [1:0] sg_in450;
  input [1:0] sg_in451;
  wire [1:0] sg_in451;
  input [1:0] sg_in452;
  wire [1:0] sg_in452;
  input [1:0] sg_in453;
  wire [1:0] sg_in453;
  input [1:0] sg_in454;
  wire [1:0] sg_in454;
  input [1:0] sg_in455;
  wire [1:0] sg_in455;
  input [1:0] sg_in456;
  wire [1:0] sg_in456;
  input [1:0] sg_in457;
  wire [1:0] sg_in457;
  input [1:0] sg_in458;
  wire [1:0] sg_in458;
  input [1:0] sg_in459;
  wire [1:0] sg_in459;
  input [1:0] sg_in460;
  wire [1:0] sg_in460;
  input [1:0] sg_in461;
  wire [1:0] sg_in461;
  input [1:0] sg_in462;
  wire [1:0] sg_in462;
  input [1:0] sg_in463;
  wire [1:0] sg_in463;
  input [1:0] sg_in464;
  wire [1:0] sg_in464;
  input [1:0] sg_in465;
  wire [1:0] sg_in465;
  input [1:0] sg_in466;
  wire [1:0] sg_in466;
  input [1:0] sg_in467;
  wire [1:0] sg_in467;
  input [1:0] sg_in468;
  wire [1:0] sg_in468;
  input [1:0] sg_in469;
  wire [1:0] sg_in469;
  input [1:0] sg_in470;
  wire [1:0] sg_in470;
  input [1:0] sg_in471;
  wire [1:0] sg_in471;
  input [1:0] sg_in472;
  wire [1:0] sg_in472;
  input [1:0] sg_in473;
  wire [1:0] sg_in473;
  input [1:0] sg_in474;
  wire [1:0] sg_in474;
  input [1:0] sg_in475;
  wire [1:0] sg_in475;
  input [1:0] sg_in476;
  wire [1:0] sg_in476;
  input [1:0] sg_in477;
  wire [1:0] sg_in477;
  input [1:0] sg_in478;
  wire [1:0] sg_in478;
  output [1:0] sg_out33;
  wire [1:0] sg_out33;
  output [1:0] sg_out34;
  wire [1:0] sg_out34;
  output [1:0] sg_out35;
  wire [1:0] sg_out35;
  output [1:0] sg_out36;
  wire [1:0] sg_out36;
  output [1:0] sg_out37;
  wire [1:0] sg_out37;
  output [1:0] sg_out38;
  wire [1:0] sg_out38;
  output [1:0] sg_out39;
  wire [1:0] sg_out39;
  output [1:0] sg_out40;
  wire [1:0] sg_out40;
  output [1:0] sg_out41;
  wire [1:0] sg_out41;
  output [1:0] sg_out42;
  wire [1:0] sg_out42;
  output [1:0] sg_out43;
  wire [1:0] sg_out43;
  output [1:0] sg_out44;
  wire [1:0] sg_out44;
  output [1:0] sg_out45;
  wire [1:0] sg_out45;
  output [1:0] sg_out46;
  wire [1:0] sg_out46;
  output [1:0] sg_out47;
  wire [1:0] sg_out47;
  output [1:0] sg_out48;
  wire [1:0] sg_out48;
  output [1:0] sg_out49;
  wire [1:0] sg_out49;
  output [1:0] sg_out50;
  wire [1:0] sg_out50;
  output [1:0] sg_out51;
  wire [1:0] sg_out51;
  output [1:0] sg_out52;
  wire [1:0] sg_out52;
  output [1:0] sg_out53;
  wire [1:0] sg_out53;
  output [1:0] sg_out54;
  wire [1:0] sg_out54;
  output [1:0] sg_out55;
  wire [1:0] sg_out55;
  output [1:0] sg_out56;
  wire [1:0] sg_out56;
  output [1:0] sg_out57;
  wire [1:0] sg_out57;
  output [1:0] sg_out58;
  wire [1:0] sg_out58;
  output [1:0] sg_out59;
  wire [1:0] sg_out59;
  output [1:0] sg_out60;
  wire [1:0] sg_out60;
  output [1:0] sg_out61;
  wire [1:0] sg_out61;
  output [9:0] sg_out62;
  wire [9:0] sg_out62;
  output [1:0] sg_out65;
  wire [1:0] sg_out65;
  output [1:0] sg_out66;
  wire [1:0] sg_out66;
  output [1:0] sg_out67;
  wire [1:0] sg_out67;
  output [1:0] sg_out68;
  wire [1:0] sg_out68;
  output [1:0] sg_out69;
  wire [1:0] sg_out69;
  output [1:0] sg_out70;
  wire [1:0] sg_out70;
  output [1:0] sg_out71;
  wire [1:0] sg_out71;
  output [1:0] sg_out72;
  wire [1:0] sg_out72;
  output [1:0] sg_out73;
  wire [1:0] sg_out73;
  output [1:0] sg_out74;
  wire [1:0] sg_out74;
  output [1:0] sg_out75;
  wire [1:0] sg_out75;
  output [1:0] sg_out76;
  wire [1:0] sg_out76;
  output [1:0] sg_out77;
  wire [1:0] sg_out77;
  output [1:0] sg_out78;
  wire [1:0] sg_out78;
  output [1:0] sg_out79;
  wire [1:0] sg_out79;
  output [1:0] sg_out80;
  wire [1:0] sg_out80;
  output [1:0] sg_out81;
  wire [1:0] sg_out81;
  output [1:0] sg_out82;
  wire [1:0] sg_out82;
  output [1:0] sg_out83;
  wire [1:0] sg_out83;
  output [1:0] sg_out84;
  wire [1:0] sg_out84;
  output [1:0] sg_out85;
  wire [1:0] sg_out85;
  output [1:0] sg_out86;
  wire [1:0] sg_out86;
  output [1:0] sg_out87;
  wire [1:0] sg_out87;
  output [1:0] sg_out88;
  wire [1:0] sg_out88;
  output [1:0] sg_out89;
  wire [1:0] sg_out89;
  output [1:0] sg_out90;
  wire [1:0] sg_out90;
  output [1:0] sg_out91;
  wire [1:0] sg_out91;
  output [1:0] sg_out92;
  wire [1:0] sg_out92;
  output [1:0] sg_out93;
  wire [1:0] sg_out93;
  output [1:0] sg_out94;
  wire [1:0] sg_out94;
  output [1:0] sg_out97;
  wire [1:0] sg_out97;
  output [1:0] sg_out98;
  wire [1:0] sg_out98;
  output [1:0] sg_out99;
  wire [1:0] sg_out99;
  output [1:0] sg_out100;
  wire [1:0] sg_out100;
  output [1:0] sg_out101;
  wire [1:0] sg_out101;
  output [1:0] sg_out102;
  wire [1:0] sg_out102;
  output [1:0] sg_out103;
  wire [1:0] sg_out103;
  output [1:0] sg_out104;
  wire [1:0] sg_out104;
  output [1:0] sg_out105;
  wire [1:0] sg_out105;
  output [1:0] sg_out106;
  wire [1:0] sg_out106;
  output [1:0] sg_out107;
  wire [1:0] sg_out107;
  output [1:0] sg_out108;
  wire [1:0] sg_out108;
  output [1:0] sg_out109;
  wire [1:0] sg_out109;
  output [1:0] sg_out110;
  wire [1:0] sg_out110;
  output [1:0] sg_out111;
  wire [1:0] sg_out111;
  output [1:0] sg_out112;
  wire [1:0] sg_out112;
  output [1:0] sg_out113;
  wire [1:0] sg_out113;
  output [1:0] sg_out114;
  wire [1:0] sg_out114;
  output [1:0] sg_out115;
  wire [1:0] sg_out115;
  output [1:0] sg_out116;
  wire [1:0] sg_out116;
  output [1:0] sg_out117;
  wire [1:0] sg_out117;
  output [1:0] sg_out118;
  wire [1:0] sg_out118;
  output [1:0] sg_out119;
  wire [1:0] sg_out119;
  output [1:0] sg_out120;
  wire [1:0] sg_out120;
  output [1:0] sg_out121;
  wire [1:0] sg_out121;
  output [1:0] sg_out122;
  wire [1:0] sg_out122;
  output [1:0] sg_out123;
  wire [1:0] sg_out123;
  output [1:0] sg_out124;
  wire [1:0] sg_out124;
  output [1:0] sg_out125;
  wire [1:0] sg_out125;
  output [1:0] sg_out126;
  wire [1:0] sg_out126;
  output [1:0] sg_out129;
  wire [1:0] sg_out129;
  output [1:0] sg_out130;
  wire [1:0] sg_out130;
  output [1:0] sg_out131;
  wire [1:0] sg_out131;
  output [1:0] sg_out132;
  wire [1:0] sg_out132;
  output [1:0] sg_out133;
  wire [1:0] sg_out133;
  output [1:0] sg_out134;
  wire [1:0] sg_out134;
  output [1:0] sg_out135;
  wire [1:0] sg_out135;
  output [1:0] sg_out136;
  wire [1:0] sg_out136;
  output [1:0] sg_out137;
  wire [1:0] sg_out137;
  output [1:0] sg_out138;
  wire [1:0] sg_out138;
  output [1:0] sg_out139;
  wire [1:0] sg_out139;
  output [1:0] sg_out140;
  wire [1:0] sg_out140;
  output [1:0] sg_out141;
  wire [1:0] sg_out141;
  output [1:0] sg_out142;
  wire [1:0] sg_out142;
  output [1:0] sg_out143;
  wire [1:0] sg_out143;
  output [1:0] sg_out144;
  wire [1:0] sg_out144;
  output [1:0] sg_out145;
  wire [1:0] sg_out145;
  output [1:0] sg_out146;
  wire [1:0] sg_out146;
  output [1:0] sg_out147;
  wire [1:0] sg_out147;
  output [1:0] sg_out148;
  wire [1:0] sg_out148;
  output [1:0] sg_out149;
  wire [1:0] sg_out149;
  output [1:0] sg_out150;
  wire [1:0] sg_out150;
  output [1:0] sg_out151;
  wire [1:0] sg_out151;
  output [1:0] sg_out152;
  wire [1:0] sg_out152;
  output [1:0] sg_out153;
  wire [1:0] sg_out153;
  output [1:0] sg_out154;
  wire [1:0] sg_out154;
  output [1:0] sg_out155;
  wire [1:0] sg_out155;
  output [1:0] sg_out156;
  wire [1:0] sg_out156;
  output [1:0] sg_out157;
  wire [1:0] sg_out157;
  output [1:0] sg_out158;
  wire [1:0] sg_out158;
  output [1:0] sg_out161;
  wire [1:0] sg_out161;
  output [1:0] sg_out162;
  wire [1:0] sg_out162;
  output [1:0] sg_out163;
  wire [1:0] sg_out163;
  output [1:0] sg_out164;
  wire [1:0] sg_out164;
  output [1:0] sg_out165;
  wire [1:0] sg_out165;
  output [1:0] sg_out166;
  wire [1:0] sg_out166;
  output [1:0] sg_out167;
  wire [1:0] sg_out167;
  output [1:0] sg_out168;
  wire [1:0] sg_out168;
  output [1:0] sg_out169;
  wire [1:0] sg_out169;
  output [1:0] sg_out170;
  wire [1:0] sg_out170;
  output [1:0] sg_out171;
  wire [1:0] sg_out171;
  output [1:0] sg_out172;
  wire [1:0] sg_out172;
  output [1:0] sg_out173;
  wire [1:0] sg_out173;
  output [1:0] sg_out174;
  wire [1:0] sg_out174;
  output [1:0] sg_out175;
  wire [1:0] sg_out175;
  output [1:0] sg_out176;
  wire [1:0] sg_out176;
  output [1:0] sg_out177;
  wire [1:0] sg_out177;
  output [1:0] sg_out178;
  wire [1:0] sg_out178;
  output [1:0] sg_out179;
  wire [1:0] sg_out179;
  output [1:0] sg_out180;
  wire [1:0] sg_out180;
  output [1:0] sg_out181;
  wire [1:0] sg_out181;
  output [1:0] sg_out182;
  wire [1:0] sg_out182;
  output [1:0] sg_out183;
  wire [1:0] sg_out183;
  output [1:0] sg_out184;
  wire [1:0] sg_out184;
  output [1:0] sg_out185;
  wire [1:0] sg_out185;
  output [1:0] sg_out186;
  wire [1:0] sg_out186;
  output [1:0] sg_out187;
  wire [1:0] sg_out187;
  output [1:0] sg_out188;
  wire [1:0] sg_out188;
  output [1:0] sg_out189;
  wire [1:0] sg_out189;
  output [1:0] sg_out190;
  wire [1:0] sg_out190;
  output [1:0] sg_out193;
  wire [1:0] sg_out193;
  output [1:0] sg_out194;
  wire [1:0] sg_out194;
  output [1:0] sg_out195;
  wire [1:0] sg_out195;
  output [1:0] sg_out196;
  wire [1:0] sg_out196;
  output [1:0] sg_out197;
  wire [1:0] sg_out197;
  output [1:0] sg_out198;
  wire [1:0] sg_out198;
  output [1:0] sg_out199;
  wire [1:0] sg_out199;
  output [1:0] sg_out200;
  wire [1:0] sg_out200;
  output [1:0] sg_out201;
  wire [1:0] sg_out201;
  output [1:0] sg_out202;
  wire [1:0] sg_out202;
  output [1:0] sg_out203;
  wire [1:0] sg_out203;
  output [1:0] sg_out204;
  wire [1:0] sg_out204;
  output [1:0] sg_out205;
  wire [1:0] sg_out205;
  output [1:0] sg_out206;
  wire [1:0] sg_out206;
  output [1:0] sg_out207;
  wire [1:0] sg_out207;
  output [1:0] sg_out208;
  wire [1:0] sg_out208;
  output [1:0] sg_out209;
  wire [1:0] sg_out209;
  output [1:0] sg_out210;
  wire [1:0] sg_out210;
  output [1:0] sg_out211;
  wire [1:0] sg_out211;
  output [1:0] sg_out212;
  wire [1:0] sg_out212;
  output [1:0] sg_out213;
  wire [1:0] sg_out213;
  output [1:0] sg_out214;
  wire [1:0] sg_out214;
  output [1:0] sg_out215;
  wire [1:0] sg_out215;
  output [1:0] sg_out216;
  wire [1:0] sg_out216;
  output [1:0] sg_out217;
  wire [1:0] sg_out217;
  output [1:0] sg_out218;
  wire [1:0] sg_out218;
  output [1:0] sg_out219;
  wire [1:0] sg_out219;
  output [1:0] sg_out220;
  wire [1:0] sg_out220;
  output [1:0] sg_out221;
  wire [1:0] sg_out221;
  output [1:0] sg_out222;
  wire [1:0] sg_out222;
  output [1:0] sg_out225;
  wire [1:0] sg_out225;
  output [1:0] sg_out226;
  wire [1:0] sg_out226;
  output [1:0] sg_out227;
  wire [1:0] sg_out227;
  output [1:0] sg_out228;
  wire [1:0] sg_out228;
  output [1:0] sg_out229;
  wire [1:0] sg_out229;
  output [1:0] sg_out230;
  wire [1:0] sg_out230;
  output [1:0] sg_out231;
  wire [1:0] sg_out231;
  output [1:0] sg_out232;
  wire [1:0] sg_out232;
  output [1:0] sg_out233;
  wire [1:0] sg_out233;
  output [1:0] sg_out234;
  wire [1:0] sg_out234;
  output [1:0] sg_out235;
  wire [1:0] sg_out235;
  output [1:0] sg_out236;
  wire [1:0] sg_out236;
  output [1:0] sg_out237;
  wire [1:0] sg_out237;
  output [1:0] sg_out238;
  wire [1:0] sg_out238;
  output [1:0] sg_out239;
  wire [1:0] sg_out239;
  output [1:0] sg_out240;
  wire [1:0] sg_out240;
  output [1:0] sg_out241;
  wire [1:0] sg_out241;
  output [1:0] sg_out242;
  wire [1:0] sg_out242;
  output [1:0] sg_out243;
  wire [1:0] sg_out243;
  output [1:0] sg_out244;
  wire [1:0] sg_out244;
  output [1:0] sg_out245;
  wire [1:0] sg_out245;
  output [1:0] sg_out246;
  wire [1:0] sg_out246;
  output [1:0] sg_out247;
  wire [1:0] sg_out247;
  output [1:0] sg_out248;
  wire [1:0] sg_out248;
  output [1:0] sg_out249;
  wire [1:0] sg_out249;
  output [1:0] sg_out250;
  wire [1:0] sg_out250;
  output [1:0] sg_out251;
  wire [1:0] sg_out251;
  output [1:0] sg_out252;
  wire [1:0] sg_out252;
  output [1:0] sg_out253;
  wire [1:0] sg_out253;
  output [1:0] sg_out254;
  wire [1:0] sg_out254;
  output [1:0] sg_out257;
  wire [1:0] sg_out257;
  output [1:0] sg_out258;
  wire [1:0] sg_out258;
  output [1:0] sg_out259;
  wire [1:0] sg_out259;
  output [1:0] sg_out260;
  wire [1:0] sg_out260;
  output [1:0] sg_out261;
  wire [1:0] sg_out261;
  output [1:0] sg_out262;
  wire [1:0] sg_out262;
  output [1:0] sg_out263;
  wire [1:0] sg_out263;
  output [1:0] sg_out264;
  wire [1:0] sg_out264;
  output [1:0] sg_out265;
  wire [1:0] sg_out265;
  output [1:0] sg_out266;
  wire [1:0] sg_out266;
  output [1:0] sg_out267;
  wire [1:0] sg_out267;
  output [1:0] sg_out268;
  wire [1:0] sg_out268;
  output [1:0] sg_out269;
  wire [1:0] sg_out269;
  output [1:0] sg_out270;
  wire [1:0] sg_out270;
  output [1:0] sg_out271;
  wire [1:0] sg_out271;
  output [1:0] sg_out272;
  wire [1:0] sg_out272;
  output [1:0] sg_out273;
  wire [1:0] sg_out273;
  output [1:0] sg_out274;
  wire [1:0] sg_out274;
  output [1:0] sg_out275;
  wire [1:0] sg_out275;
  output [1:0] sg_out276;
  wire [1:0] sg_out276;
  output [1:0] sg_out277;
  wire [1:0] sg_out277;
  output [1:0] sg_out278;
  wire [1:0] sg_out278;
  output [1:0] sg_out279;
  wire [1:0] sg_out279;
  output [1:0] sg_out280;
  wire [1:0] sg_out280;
  output [1:0] sg_out281;
  wire [1:0] sg_out281;
  output [1:0] sg_out282;
  wire [1:0] sg_out282;
  output [1:0] sg_out283;
  wire [1:0] sg_out283;
  output [1:0] sg_out284;
  wire [1:0] sg_out284;
  output [1:0] sg_out285;
  wire [1:0] sg_out285;
  output [1:0] sg_out286;
  wire [1:0] sg_out286;
  output [1:0] sg_out289;
  wire [1:0] sg_out289;
  output [1:0] sg_out290;
  wire [1:0] sg_out290;
  output [1:0] sg_out291;
  wire [1:0] sg_out291;
  output [1:0] sg_out292;
  wire [1:0] sg_out292;
  output [1:0] sg_out293;
  wire [1:0] sg_out293;
  output [1:0] sg_out294;
  wire [1:0] sg_out294;
  output [1:0] sg_out295;
  wire [1:0] sg_out295;
  output [1:0] sg_out296;
  wire [1:0] sg_out296;
  output [1:0] sg_out297;
  wire [1:0] sg_out297;
  output [1:0] sg_out298;
  wire [1:0] sg_out298;
  output [1:0] sg_out299;
  wire [1:0] sg_out299;
  output [1:0] sg_out300;
  wire [1:0] sg_out300;
  output [1:0] sg_out301;
  wire [1:0] sg_out301;
  output [1:0] sg_out302;
  wire [1:0] sg_out302;
  output [1:0] sg_out303;
  wire [1:0] sg_out303;
  output [1:0] sg_out304;
  wire [1:0] sg_out304;
  output [1:0] sg_out305;
  wire [1:0] sg_out305;
  output [1:0] sg_out306;
  wire [1:0] sg_out306;
  output [1:0] sg_out307;
  wire [1:0] sg_out307;
  output [1:0] sg_out308;
  wire [1:0] sg_out308;
  output [1:0] sg_out309;
  wire [1:0] sg_out309;
  output [1:0] sg_out310;
  wire [1:0] sg_out310;
  output [1:0] sg_out311;
  wire [1:0] sg_out311;
  output [1:0] sg_out312;
  wire [1:0] sg_out312;
  output [1:0] sg_out313;
  wire [1:0] sg_out313;
  output [1:0] sg_out314;
  wire [1:0] sg_out314;
  output [1:0] sg_out315;
  wire [1:0] sg_out315;
  output [1:0] sg_out316;
  wire [1:0] sg_out316;
  output [1:0] sg_out317;
  wire [1:0] sg_out317;
  output [1:0] sg_out318;
  wire [1:0] sg_out318;
  output [1:0] sg_out321;
  wire [1:0] sg_out321;
  output [1:0] sg_out322;
  wire [1:0] sg_out322;
  output [1:0] sg_out323;
  wire [1:0] sg_out323;
  output [1:0] sg_out324;
  wire [1:0] sg_out324;
  output [1:0] sg_out325;
  wire [1:0] sg_out325;
  output [1:0] sg_out326;
  wire [1:0] sg_out326;
  output [1:0] sg_out327;
  wire [1:0] sg_out327;
  output [1:0] sg_out328;
  wire [1:0] sg_out328;
  output [1:0] sg_out329;
  wire [1:0] sg_out329;
  output [1:0] sg_out330;
  wire [1:0] sg_out330;
  output [1:0] sg_out331;
  wire [1:0] sg_out331;
  output [1:0] sg_out332;
  wire [1:0] sg_out332;
  output [1:0] sg_out333;
  wire [1:0] sg_out333;
  output [1:0] sg_out334;
  wire [1:0] sg_out334;
  output [1:0] sg_out335;
  wire [1:0] sg_out335;
  output [1:0] sg_out336;
  wire [1:0] sg_out336;
  output [1:0] sg_out337;
  wire [1:0] sg_out337;
  output [1:0] sg_out338;
  wire [1:0] sg_out338;
  output [1:0] sg_out339;
  wire [1:0] sg_out339;
  output [1:0] sg_out340;
  wire [1:0] sg_out340;
  output [1:0] sg_out341;
  wire [1:0] sg_out341;
  output [1:0] sg_out342;
  wire [1:0] sg_out342;
  output [1:0] sg_out343;
  wire [1:0] sg_out343;
  output [1:0] sg_out344;
  wire [1:0] sg_out344;
  output [1:0] sg_out345;
  wire [1:0] sg_out345;
  output [1:0] sg_out346;
  wire [1:0] sg_out346;
  output [1:0] sg_out347;
  wire [1:0] sg_out347;
  output [1:0] sg_out348;
  wire [1:0] sg_out348;
  output [1:0] sg_out349;
  wire [1:0] sg_out349;
  output [1:0] sg_out350;
  wire [1:0] sg_out350;
  output [1:0] sg_out353;
  wire [1:0] sg_out353;
  output [1:0] sg_out354;
  wire [1:0] sg_out354;
  output [1:0] sg_out355;
  wire [1:0] sg_out355;
  output [1:0] sg_out356;
  wire [1:0] sg_out356;
  output [1:0] sg_out357;
  wire [1:0] sg_out357;
  output [1:0] sg_out358;
  wire [1:0] sg_out358;
  output [1:0] sg_out359;
  wire [1:0] sg_out359;
  output [1:0] sg_out360;
  wire [1:0] sg_out360;
  output [1:0] sg_out361;
  wire [1:0] sg_out361;
  output [1:0] sg_out362;
  wire [1:0] sg_out362;
  output [1:0] sg_out363;
  wire [1:0] sg_out363;
  output [1:0] sg_out364;
  wire [1:0] sg_out364;
  output [1:0] sg_out365;
  wire [1:0] sg_out365;
  output [1:0] sg_out366;
  wire [1:0] sg_out366;
  output [1:0] sg_out367;
  wire [1:0] sg_out367;
  output [1:0] sg_out368;
  wire [1:0] sg_out368;
  output [1:0] sg_out369;
  wire [1:0] sg_out369;
  output [1:0] sg_out370;
  wire [1:0] sg_out370;
  output [1:0] sg_out371;
  wire [1:0] sg_out371;
  output [1:0] sg_out372;
  wire [1:0] sg_out372;
  output [1:0] sg_out373;
  wire [1:0] sg_out373;
  output [1:0] sg_out374;
  wire [1:0] sg_out374;
  output [1:0] sg_out375;
  wire [1:0] sg_out375;
  output [1:0] sg_out376;
  wire [1:0] sg_out376;
  output [1:0] sg_out377;
  wire [1:0] sg_out377;
  output [1:0] sg_out378;
  wire [1:0] sg_out378;
  output [1:0] sg_out379;
  wire [1:0] sg_out379;
  output [1:0] sg_out380;
  wire [1:0] sg_out380;
  output [1:0] sg_out381;
  wire [1:0] sg_out381;
  output [1:0] sg_out382;
  wire [1:0] sg_out382;
  output [1:0] sg_out385;
  wire [1:0] sg_out385;
  output [1:0] sg_out386;
  wire [1:0] sg_out386;
  output [1:0] sg_out387;
  wire [1:0] sg_out387;
  output [1:0] sg_out388;
  wire [1:0] sg_out388;
  output [1:0] sg_out389;
  wire [1:0] sg_out389;
  output [1:0] sg_out390;
  wire [1:0] sg_out390;
  output [1:0] sg_out391;
  wire [1:0] sg_out391;
  output [1:0] sg_out392;
  wire [1:0] sg_out392;
  output [1:0] sg_out393;
  wire [1:0] sg_out393;
  output [1:0] sg_out394;
  wire [1:0] sg_out394;
  output [1:0] sg_out395;
  wire [1:0] sg_out395;
  output [1:0] sg_out396;
  wire [1:0] sg_out396;
  output [1:0] sg_out397;
  wire [1:0] sg_out397;
  output [1:0] sg_out398;
  wire [1:0] sg_out398;
  output [1:0] sg_out399;
  wire [1:0] sg_out399;
  output [1:0] sg_out400;
  wire [1:0] sg_out400;
  output [1:0] sg_out401;
  wire [1:0] sg_out401;
  output [1:0] sg_out402;
  wire [1:0] sg_out402;
  output [1:0] sg_out403;
  wire [1:0] sg_out403;
  output [1:0] sg_out404;
  wire [1:0] sg_out404;
  output [1:0] sg_out405;
  wire [1:0] sg_out405;
  output [1:0] sg_out406;
  wire [1:0] sg_out406;
  output [1:0] sg_out407;
  wire [1:0] sg_out407;
  output [1:0] sg_out408;
  wire [1:0] sg_out408;
  output [1:0] sg_out409;
  wire [1:0] sg_out409;
  output [1:0] sg_out410;
  wire [1:0] sg_out410;
  output [1:0] sg_out411;
  wire [1:0] sg_out411;
  output [1:0] sg_out412;
  wire [1:0] sg_out412;
  output [1:0] sg_out413;
  wire [1:0] sg_out413;
  output [1:0] sg_out414;
  wire [1:0] sg_out414;
  output [1:0] sg_out417;
  wire [1:0] sg_out417;
  output [1:0] sg_out418;
  wire [1:0] sg_out418;
  output [1:0] sg_out419;
  wire [1:0] sg_out419;
  output [1:0] sg_out420;
  wire [1:0] sg_out420;
  output [1:0] sg_out421;
  wire [1:0] sg_out421;
  output [1:0] sg_out422;
  wire [1:0] sg_out422;
  output [1:0] sg_out423;
  wire [1:0] sg_out423;
  output [1:0] sg_out424;
  wire [1:0] sg_out424;
  output [1:0] sg_out425;
  wire [1:0] sg_out425;
  output [1:0] sg_out426;
  wire [1:0] sg_out426;
  output [1:0] sg_out427;
  wire [1:0] sg_out427;
  output [1:0] sg_out428;
  wire [1:0] sg_out428;
  output [1:0] sg_out429;
  wire [1:0] sg_out429;
  output [1:0] sg_out430;
  wire [1:0] sg_out430;
  output [1:0] sg_out431;
  wire [1:0] sg_out431;
  output [1:0] sg_out432;
  wire [1:0] sg_out432;
  output [1:0] sg_out433;
  wire [1:0] sg_out433;
  output [1:0] sg_out434;
  wire [1:0] sg_out434;
  output [1:0] sg_out435;
  wire [1:0] sg_out435;
  output [1:0] sg_out436;
  wire [1:0] sg_out436;
  output [1:0] sg_out437;
  wire [1:0] sg_out437;
  output [1:0] sg_out438;
  wire [1:0] sg_out438;
  output [1:0] sg_out439;
  wire [1:0] sg_out439;
  output [1:0] sg_out440;
  wire [1:0] sg_out440;
  output [1:0] sg_out441;
  wire [1:0] sg_out441;
  output [1:0] sg_out442;
  wire [1:0] sg_out442;
  output [1:0] sg_out443;
  wire [1:0] sg_out443;
  output [1:0] sg_out444;
  wire [1:0] sg_out444;
  output [1:0] sg_out445;
  wire [1:0] sg_out445;
  output [1:0] sg_out446;
  wire [1:0] sg_out446;
  output [1:0] sg_out449;
  wire [1:0] sg_out449;
  output [1:0] sg_out450;
  wire [1:0] sg_out450;
  output [1:0] sg_out451;
  wire [1:0] sg_out451;
  output [1:0] sg_out452;
  wire [1:0] sg_out452;
  output [1:0] sg_out453;
  wire [1:0] sg_out453;
  output [1:0] sg_out454;
  wire [1:0] sg_out454;
  output [1:0] sg_out455;
  wire [1:0] sg_out455;
  output [1:0] sg_out456;
  wire [1:0] sg_out456;
  output [1:0] sg_out457;
  wire [1:0] sg_out457;
  output [1:0] sg_out458;
  wire [1:0] sg_out458;
  output [1:0] sg_out459;
  wire [1:0] sg_out459;
  output [1:0] sg_out460;
  wire [1:0] sg_out460;
  output [1:0] sg_out461;
  wire [1:0] sg_out461;
  output [1:0] sg_out462;
  wire [1:0] sg_out462;
  output [1:0] sg_out463;
  wire [1:0] sg_out463;
  output [1:0] sg_out464;
  wire [1:0] sg_out464;
  output [1:0] sg_out465;
  wire [1:0] sg_out465;
  output [1:0] sg_out466;
  wire [1:0] sg_out466;
  output [1:0] sg_out467;
  wire [1:0] sg_out467;
  output [1:0] sg_out468;
  wire [1:0] sg_out468;
  output [1:0] sg_out469;
  wire [1:0] sg_out469;
  output [1:0] sg_out470;
  wire [1:0] sg_out470;
  output [1:0] sg_out471;
  wire [1:0] sg_out471;
  output [1:0] sg_out472;
  wire [1:0] sg_out472;
  output [1:0] sg_out473;
  wire [1:0] sg_out473;
  output [1:0] sg_out474;
  wire [1:0] sg_out474;
  output [1:0] sg_out475;
  wire [1:0] sg_out475;
  output [1:0] sg_out476;
  wire [1:0] sg_out476;
  output [1:0] sg_out477;
  wire [1:0] sg_out477;
  output [1:0] sg_out478;
  wire [1:0] sg_out478;
  output dig_t0;
  wire dig_t0;
  output dig_t1;
  wire dig_t1;
  output dig_t2;
  wire dig_t2;
  output dig_t3;
  wire dig_t3;
  output dig_t4;
  wire dig_t4;
  output dig_t5;
  wire dig_t5;
  output dig_t6;
  wire dig_t6;
  output dig_t7;
  wire dig_t7;
  output dig_t8;
  wire dig_t8;
  output dig_t9;
  wire dig_t9;
  output dig_t10;
  wire dig_t10;
  output dig_t11;
  wire dig_t11;
  output dig_t12;
  wire dig_t12;
  output dig_t13;
  wire dig_t13;
  output dig_t14;
  wire dig_t14;
  output dig_t15;
  wire dig_t15;
  output dig_t16;
  wire dig_t16;
  output dig_t17;
  wire dig_t17;
  output dig_t18;
  wire dig_t18;
  output dig_t19;
  wire dig_t19;
  output dig_t20;
  wire dig_t20;
  output dig_t21;
  wire dig_t21;
  output dig_t22;
  wire dig_t22;
  output dig_t23;
  wire dig_t23;
  output dig_t24;
  wire dig_t24;
  output dig_t25;
  wire dig_t25;
  output dig_t26;
  wire dig_t26;
  output dig_t27;
  wire dig_t27;
  output dig_t28;
  wire dig_t28;
  output dig_t29;
  wire dig_t29;
  output dig_t30;
  wire dig_t30;
  output dig_t31;
  wire dig_t31;
  output dig_t32;
  wire dig_t32;
  output dig_t33;
  wire dig_t33;
  output dig_t34;
  wire dig_t34;
  output dig_t35;
  wire dig_t35;
  output dig_t36;
  wire dig_t36;
  output dig_t37;
  wire dig_t37;
  output dig_t38;
  wire dig_t38;
  output dig_t39;
  wire dig_t39;
  output dig_t40;
  wire dig_t40;
  output dig_t41;
  wire dig_t41;
  output dig_t42;
  wire dig_t42;
  output dig_t43;
  wire dig_t43;
  output dig_t44;
  wire dig_t44;
  output dig_t45;
  wire dig_t45;
  output dig_t46;
  wire dig_t46;
  output dig_t47;
  wire dig_t47;
  output dig_t48;
  wire dig_t48;
  output dig_t49;
  wire dig_t49;
  output dig_t50;
  wire dig_t50;
  output dig_t51;
  wire dig_t51;
  output dig_t52;
  wire dig_t52;
  output dig_t53;
  wire dig_t53;
  output dig_t54;
  wire dig_t54;
  output dig_t55;
  wire dig_t55;
  output dig_t56;
  wire dig_t56;
  output dig_t57;
  wire dig_t57;
  output dig_t58;
  wire dig_t58;
  output dig_t59;
  wire dig_t59;
  output dig_t60;
  wire dig_t60;
  output dig_t61;
  wire dig_t61;
  output dig_t62;
  wire dig_t62;
  output dig_t63;
  wire dig_t63;
  output dig_t64;
  wire dig_t64;
  output dig_t65;
  wire dig_t65;
  output dig_t66;
  wire dig_t66;
  output dig_t67;
  wire dig_t67;
  output dig_t68;
  wire dig_t68;
  output dig_t69;
  wire dig_t69;
  output dig_t70;
  wire dig_t70;
  output dig_t71;
  wire dig_t71;
  output dig_t72;
  wire dig_t72;
  output dig_t73;
  wire dig_t73;
  output dig_t74;
  wire dig_t74;
  output dig_t75;
  wire dig_t75;
  output dig_t76;
  wire dig_t76;
  output dig_t77;
  wire dig_t77;
  output dig_t78;
  wire dig_t78;
  output dig_t79;
  wire dig_t79;
  output dig_t80;
  wire dig_t80;
  output dig_t81;
  wire dig_t81;
  output dig_t82;
  wire dig_t82;
  output dig_t83;
  wire dig_t83;
  output dig_t84;
  wire dig_t84;
  output dig_t85;
  wire dig_t85;
  output dig_t86;
  wire dig_t86;
  output dig_t87;
  wire dig_t87;
  output dig_t88;
  wire dig_t88;
  output dig_t89;
  wire dig_t89;
  output dig_t90;
  wire dig_t90;
  output dig_t91;
  wire dig_t91;
  output dig_t92;
  wire dig_t92;
  output dig_t93;
  wire dig_t93;
  output dig_t94;
  wire dig_t94;
  output dig_t95;
  wire dig_t95;
  output dig_t96;
  wire dig_t96;
  output dig_t97;
  wire dig_t97;
  output dig_t98;
  wire dig_t98;
  output dig_t99;
  wire dig_t99;
  output dig_t100;
  wire dig_t100;
  output dig_t101;
  wire dig_t101;
  output dig_t102;
  wire dig_t102;
  output dig_t103;
  wire dig_t103;
  output dig_t104;
  wire dig_t104;
  output dig_t105;
  wire dig_t105;
  output dig_t106;
  wire dig_t106;
  output dig_t107;
  wire dig_t107;
  output dig_t108;
  wire dig_t108;
  output dig_t109;
  wire dig_t109;
  output dig_t110;
  wire dig_t110;
  output dig_t111;
  wire dig_t111;
  output dig_t112;
  wire dig_t112;
  output dig_t113;
  wire dig_t113;
  output dig_t114;
  wire dig_t114;
  output dig_t115;
  wire dig_t115;
  output dig_t116;
  wire dig_t116;
  output dig_t117;
  wire dig_t117;
  output dig_t118;
  wire dig_t118;
  output dig_t119;
  wire dig_t119;
  output dig_t120;
  wire dig_t120;
  output dig_t121;
  wire dig_t121;
  output dig_t122;
  wire dig_t122;
  output dig_t123;
  wire dig_t123;
  output dig_t124;
  wire dig_t124;
  output dig_t125;
  wire dig_t125;
  output dig_t126;
  wire dig_t126;
  output dig_t127;
  wire dig_t127;
  output dig_t128;
  wire dig_t128;
  output dig_t129;
  wire dig_t129;
  output dig_t130;
  wire dig_t130;
  output dig_t131;
  wire dig_t131;
  output dig_t132;
  wire dig_t132;
  output dig_t133;
  wire dig_t133;
  output dig_t134;
  wire dig_t134;
  output dig_t135;
  wire dig_t135;
  output dig_t136;
  wire dig_t136;
  output dig_t137;
  wire dig_t137;
  output dig_t138;
  wire dig_t138;
  output dig_t139;
  wire dig_t139;
  output dig_t140;
  wire dig_t140;
  output dig_t141;
  wire dig_t141;
  output dig_t142;
  wire dig_t142;
  output dig_t143;
  wire dig_t143;
  output dig_t144;
  wire dig_t144;
  output dig_t145;
  wire dig_t145;
  output dig_t146;
  wire dig_t146;
  output dig_t147;
  wire dig_t147;
  output dig_t148;
  wire dig_t148;
  output dig_t149;
  wire dig_t149;
  output dig_t150;
  wire dig_t150;
  output dig_t151;
  wire dig_t151;
  output dig_t152;
  wire dig_t152;
  output dig_t153;
  wire dig_t153;
  output dig_t154;
  wire dig_t154;
  output dig_t155;
  wire dig_t155;
  output dig_t156;
  wire dig_t156;
  output dig_t157;
  wire dig_t157;
  output dig_t158;
  wire dig_t158;
  output dig_t159;
  wire dig_t159;
  output dig_t160;
  wire dig_t160;
  output dig_t161;
  wire dig_t161;
  output dig_t162;
  wire dig_t162;
  output dig_t163;
  wire dig_t163;
  output dig_t164;
  wire dig_t164;
  output dig_t165;
  wire dig_t165;
  output dig_t166;
  wire dig_t166;
  output dig_t167;
  wire dig_t167;
  output dig_t168;
  wire dig_t168;
  output dig_t169;
  wire dig_t169;
  output dig_t170;
  wire dig_t170;
  output dig_t171;
  wire dig_t171;
  output dig_t172;
  wire dig_t172;
  output dig_t173;
  wire dig_t173;
  output dig_t174;
  wire dig_t174;
  output dig_t175;
  wire dig_t175;
  output dig_t176;
  wire dig_t176;
  output dig_t177;
  wire dig_t177;
  output dig_t178;
  wire dig_t178;
  output dig_t179;
  wire dig_t179;
  output dig_t180;
  wire dig_t180;
  output dig_t181;
  wire dig_t181;
  output dig_t182;
  wire dig_t182;
  output dig_t183;
  wire dig_t183;
  output dig_t184;
  wire dig_t184;
  output dig_t185;
  wire dig_t185;
  output dig_t186;
  wire dig_t186;
  output dig_t187;
  wire dig_t187;
  output dig_t188;
  wire dig_t188;
  output dig_t189;
  wire dig_t189;
  output dig_t190;
  wire dig_t190;
  output dig_t191;
  wire dig_t191;
  output dig_t192;
  wire dig_t192;
  output dig_t193;
  wire dig_t193;
  output dig_t194;
  wire dig_t194;
  output dig_t195;
  wire dig_t195;
  output dig_t196;
  wire dig_t196;
  output dig_t197;
  wire dig_t197;
  output dig_t198;
  wire dig_t198;
  output dig_t199;
  wire dig_t199;
  output dig_t200;
  wire dig_t200;
  output dig_t201;
  wire dig_t201;
  output dig_t202;
  wire dig_t202;
  output dig_t203;
  wire dig_t203;
  output dig_t204;
  wire dig_t204;
  output dig_t205;
  wire dig_t205;
  output dig_t206;
  wire dig_t206;
  output dig_t207;
  wire dig_t207;
  output dig_t208;
  wire dig_t208;
  output dig_t209;
  wire dig_t209;
  input in_do;
  wire in_do;
  output out_do;
  wire out_do;
  output out_data;
  wire out_data;
  reg sig_reg;
  wire [9:0] _add_map_x_moto_org_near;
  wire [9:0] _add_map_x_moto_org_near1;
  wire [9:0] _add_map_x_moto_org_near2;
  wire [9:0] _add_map_x_moto_org_near3;
  wire [9:0] _add_map_x_moto_org;
  wire [1:0] _add_map_x_sg_up;
  wire [1:0] _add_map_x_sg_down;
  wire [1:0] _add_map_x_sg_left;
  wire [1:0] _add_map_x_sg_right;
  wire _add_map_x_wall_t_in;
  wire [9:0] _add_map_x_moto;
  wire [9:0] _add_map_x_up;
  wire [9:0] _add_map_x_right;
  wire [9:0] _add_map_x_down;
  wire [9:0] _add_map_x_left;
  wire [9:0] _add_map_x_start;
  wire [9:0] _add_map_x_goal;
  wire [9:0] _add_map_x_now;
  wire [9:0] _add_map_x_data_out;
  wire [9:0] _add_map_x_data_out_index;
  wire [9:0] _add_map_x_data_near;
  wire _add_map_x_wall_t_out;
  wire [9:0] _add_map_x_data_org;
  wire [9:0] _add_map_x_data_org_near;
  wire [1:0] _add_map_x_s_g;
  wire [1:0] _add_map_x_s_g_near;
  wire _add_map_x_add_exe;
  wire _add_map_x_p_reset;
  wire _add_map_x_m_clock;
  wire [9:0] _add_map_x_209_moto_org_near;
  wire [9:0] _add_map_x_209_moto_org_near1;
  wire [9:0] _add_map_x_209_moto_org_near2;
  wire [9:0] _add_map_x_209_moto_org_near3;
  wire [9:0] _add_map_x_209_moto_org;
  wire [1:0] _add_map_x_209_sg_up;
  wire [1:0] _add_map_x_209_sg_down;
  wire [1:0] _add_map_x_209_sg_left;
  wire [1:0] _add_map_x_209_sg_right;
  wire _add_map_x_209_wall_t_in;
  wire [9:0] _add_map_x_209_moto;
  wire [9:0] _add_map_x_209_up;
  wire [9:0] _add_map_x_209_right;
  wire [9:0] _add_map_x_209_down;
  wire [9:0] _add_map_x_209_left;
  wire [9:0] _add_map_x_209_start;
  wire [9:0] _add_map_x_209_goal;
  wire [9:0] _add_map_x_209_now;
  wire [9:0] _add_map_x_209_data_out;
  wire [9:0] _add_map_x_209_data_out_index;
  wire [9:0] _add_map_x_209_data_near;
  wire _add_map_x_209_wall_t_out;
  wire [9:0] _add_map_x_209_data_org;
  wire [9:0] _add_map_x_209_data_org_near;
  wire [1:0] _add_map_x_209_s_g;
  wire [1:0] _add_map_x_209_s_g_near;
  wire _add_map_x_209_add_exe;
  wire _add_map_x_209_p_reset;
  wire _add_map_x_209_m_clock;
  wire [9:0] _add_map_x_208_moto_org_near;
  wire [9:0] _add_map_x_208_moto_org_near1;
  wire [9:0] _add_map_x_208_moto_org_near2;
  wire [9:0] _add_map_x_208_moto_org_near3;
  wire [9:0] _add_map_x_208_moto_org;
  wire [1:0] _add_map_x_208_sg_up;
  wire [1:0] _add_map_x_208_sg_down;
  wire [1:0] _add_map_x_208_sg_left;
  wire [1:0] _add_map_x_208_sg_right;
  wire _add_map_x_208_wall_t_in;
  wire [9:0] _add_map_x_208_moto;
  wire [9:0] _add_map_x_208_up;
  wire [9:0] _add_map_x_208_right;
  wire [9:0] _add_map_x_208_down;
  wire [9:0] _add_map_x_208_left;
  wire [9:0] _add_map_x_208_start;
  wire [9:0] _add_map_x_208_goal;
  wire [9:0] _add_map_x_208_now;
  wire [9:0] _add_map_x_208_data_out;
  wire [9:0] _add_map_x_208_data_out_index;
  wire [9:0] _add_map_x_208_data_near;
  wire _add_map_x_208_wall_t_out;
  wire [9:0] _add_map_x_208_data_org;
  wire [9:0] _add_map_x_208_data_org_near;
  wire [1:0] _add_map_x_208_s_g;
  wire [1:0] _add_map_x_208_s_g_near;
  wire _add_map_x_208_add_exe;
  wire _add_map_x_208_p_reset;
  wire _add_map_x_208_m_clock;
  wire [9:0] _add_map_x_207_moto_org_near;
  wire [9:0] _add_map_x_207_moto_org_near1;
  wire [9:0] _add_map_x_207_moto_org_near2;
  wire [9:0] _add_map_x_207_moto_org_near3;
  wire [9:0] _add_map_x_207_moto_org;
  wire [1:0] _add_map_x_207_sg_up;
  wire [1:0] _add_map_x_207_sg_down;
  wire [1:0] _add_map_x_207_sg_left;
  wire [1:0] _add_map_x_207_sg_right;
  wire _add_map_x_207_wall_t_in;
  wire [9:0] _add_map_x_207_moto;
  wire [9:0] _add_map_x_207_up;
  wire [9:0] _add_map_x_207_right;
  wire [9:0] _add_map_x_207_down;
  wire [9:0] _add_map_x_207_left;
  wire [9:0] _add_map_x_207_start;
  wire [9:0] _add_map_x_207_goal;
  wire [9:0] _add_map_x_207_now;
  wire [9:0] _add_map_x_207_data_out;
  wire [9:0] _add_map_x_207_data_out_index;
  wire [9:0] _add_map_x_207_data_near;
  wire _add_map_x_207_wall_t_out;
  wire [9:0] _add_map_x_207_data_org;
  wire [9:0] _add_map_x_207_data_org_near;
  wire [1:0] _add_map_x_207_s_g;
  wire [1:0] _add_map_x_207_s_g_near;
  wire _add_map_x_207_add_exe;
  wire _add_map_x_207_p_reset;
  wire _add_map_x_207_m_clock;
  wire [9:0] _add_map_x_206_moto_org_near;
  wire [9:0] _add_map_x_206_moto_org_near1;
  wire [9:0] _add_map_x_206_moto_org_near2;
  wire [9:0] _add_map_x_206_moto_org_near3;
  wire [9:0] _add_map_x_206_moto_org;
  wire [1:0] _add_map_x_206_sg_up;
  wire [1:0] _add_map_x_206_sg_down;
  wire [1:0] _add_map_x_206_sg_left;
  wire [1:0] _add_map_x_206_sg_right;
  wire _add_map_x_206_wall_t_in;
  wire [9:0] _add_map_x_206_moto;
  wire [9:0] _add_map_x_206_up;
  wire [9:0] _add_map_x_206_right;
  wire [9:0] _add_map_x_206_down;
  wire [9:0] _add_map_x_206_left;
  wire [9:0] _add_map_x_206_start;
  wire [9:0] _add_map_x_206_goal;
  wire [9:0] _add_map_x_206_now;
  wire [9:0] _add_map_x_206_data_out;
  wire [9:0] _add_map_x_206_data_out_index;
  wire [9:0] _add_map_x_206_data_near;
  wire _add_map_x_206_wall_t_out;
  wire [9:0] _add_map_x_206_data_org;
  wire [9:0] _add_map_x_206_data_org_near;
  wire [1:0] _add_map_x_206_s_g;
  wire [1:0] _add_map_x_206_s_g_near;
  wire _add_map_x_206_add_exe;
  wire _add_map_x_206_p_reset;
  wire _add_map_x_206_m_clock;
  wire [9:0] _add_map_x_205_moto_org_near;
  wire [9:0] _add_map_x_205_moto_org_near1;
  wire [9:0] _add_map_x_205_moto_org_near2;
  wire [9:0] _add_map_x_205_moto_org_near3;
  wire [9:0] _add_map_x_205_moto_org;
  wire [1:0] _add_map_x_205_sg_up;
  wire [1:0] _add_map_x_205_sg_down;
  wire [1:0] _add_map_x_205_sg_left;
  wire [1:0] _add_map_x_205_sg_right;
  wire _add_map_x_205_wall_t_in;
  wire [9:0] _add_map_x_205_moto;
  wire [9:0] _add_map_x_205_up;
  wire [9:0] _add_map_x_205_right;
  wire [9:0] _add_map_x_205_down;
  wire [9:0] _add_map_x_205_left;
  wire [9:0] _add_map_x_205_start;
  wire [9:0] _add_map_x_205_goal;
  wire [9:0] _add_map_x_205_now;
  wire [9:0] _add_map_x_205_data_out;
  wire [9:0] _add_map_x_205_data_out_index;
  wire [9:0] _add_map_x_205_data_near;
  wire _add_map_x_205_wall_t_out;
  wire [9:0] _add_map_x_205_data_org;
  wire [9:0] _add_map_x_205_data_org_near;
  wire [1:0] _add_map_x_205_s_g;
  wire [1:0] _add_map_x_205_s_g_near;
  wire _add_map_x_205_add_exe;
  wire _add_map_x_205_p_reset;
  wire _add_map_x_205_m_clock;
  wire [9:0] _add_map_x_204_moto_org_near;
  wire [9:0] _add_map_x_204_moto_org_near1;
  wire [9:0] _add_map_x_204_moto_org_near2;
  wire [9:0] _add_map_x_204_moto_org_near3;
  wire [9:0] _add_map_x_204_moto_org;
  wire [1:0] _add_map_x_204_sg_up;
  wire [1:0] _add_map_x_204_sg_down;
  wire [1:0] _add_map_x_204_sg_left;
  wire [1:0] _add_map_x_204_sg_right;
  wire _add_map_x_204_wall_t_in;
  wire [9:0] _add_map_x_204_moto;
  wire [9:0] _add_map_x_204_up;
  wire [9:0] _add_map_x_204_right;
  wire [9:0] _add_map_x_204_down;
  wire [9:0] _add_map_x_204_left;
  wire [9:0] _add_map_x_204_start;
  wire [9:0] _add_map_x_204_goal;
  wire [9:0] _add_map_x_204_now;
  wire [9:0] _add_map_x_204_data_out;
  wire [9:0] _add_map_x_204_data_out_index;
  wire [9:0] _add_map_x_204_data_near;
  wire _add_map_x_204_wall_t_out;
  wire [9:0] _add_map_x_204_data_org;
  wire [9:0] _add_map_x_204_data_org_near;
  wire [1:0] _add_map_x_204_s_g;
  wire [1:0] _add_map_x_204_s_g_near;
  wire _add_map_x_204_add_exe;
  wire _add_map_x_204_p_reset;
  wire _add_map_x_204_m_clock;
  wire [9:0] _add_map_x_203_moto_org_near;
  wire [9:0] _add_map_x_203_moto_org_near1;
  wire [9:0] _add_map_x_203_moto_org_near2;
  wire [9:0] _add_map_x_203_moto_org_near3;
  wire [9:0] _add_map_x_203_moto_org;
  wire [1:0] _add_map_x_203_sg_up;
  wire [1:0] _add_map_x_203_sg_down;
  wire [1:0] _add_map_x_203_sg_left;
  wire [1:0] _add_map_x_203_sg_right;
  wire _add_map_x_203_wall_t_in;
  wire [9:0] _add_map_x_203_moto;
  wire [9:0] _add_map_x_203_up;
  wire [9:0] _add_map_x_203_right;
  wire [9:0] _add_map_x_203_down;
  wire [9:0] _add_map_x_203_left;
  wire [9:0] _add_map_x_203_start;
  wire [9:0] _add_map_x_203_goal;
  wire [9:0] _add_map_x_203_now;
  wire [9:0] _add_map_x_203_data_out;
  wire [9:0] _add_map_x_203_data_out_index;
  wire [9:0] _add_map_x_203_data_near;
  wire _add_map_x_203_wall_t_out;
  wire [9:0] _add_map_x_203_data_org;
  wire [9:0] _add_map_x_203_data_org_near;
  wire [1:0] _add_map_x_203_s_g;
  wire [1:0] _add_map_x_203_s_g_near;
  wire _add_map_x_203_add_exe;
  wire _add_map_x_203_p_reset;
  wire _add_map_x_203_m_clock;
  wire [9:0] _add_map_x_202_moto_org_near;
  wire [9:0] _add_map_x_202_moto_org_near1;
  wire [9:0] _add_map_x_202_moto_org_near2;
  wire [9:0] _add_map_x_202_moto_org_near3;
  wire [9:0] _add_map_x_202_moto_org;
  wire [1:0] _add_map_x_202_sg_up;
  wire [1:0] _add_map_x_202_sg_down;
  wire [1:0] _add_map_x_202_sg_left;
  wire [1:0] _add_map_x_202_sg_right;
  wire _add_map_x_202_wall_t_in;
  wire [9:0] _add_map_x_202_moto;
  wire [9:0] _add_map_x_202_up;
  wire [9:0] _add_map_x_202_right;
  wire [9:0] _add_map_x_202_down;
  wire [9:0] _add_map_x_202_left;
  wire [9:0] _add_map_x_202_start;
  wire [9:0] _add_map_x_202_goal;
  wire [9:0] _add_map_x_202_now;
  wire [9:0] _add_map_x_202_data_out;
  wire [9:0] _add_map_x_202_data_out_index;
  wire [9:0] _add_map_x_202_data_near;
  wire _add_map_x_202_wall_t_out;
  wire [9:0] _add_map_x_202_data_org;
  wire [9:0] _add_map_x_202_data_org_near;
  wire [1:0] _add_map_x_202_s_g;
  wire [1:0] _add_map_x_202_s_g_near;
  wire _add_map_x_202_add_exe;
  wire _add_map_x_202_p_reset;
  wire _add_map_x_202_m_clock;
  wire [9:0] _add_map_x_201_moto_org_near;
  wire [9:0] _add_map_x_201_moto_org_near1;
  wire [9:0] _add_map_x_201_moto_org_near2;
  wire [9:0] _add_map_x_201_moto_org_near3;
  wire [9:0] _add_map_x_201_moto_org;
  wire [1:0] _add_map_x_201_sg_up;
  wire [1:0] _add_map_x_201_sg_down;
  wire [1:0] _add_map_x_201_sg_left;
  wire [1:0] _add_map_x_201_sg_right;
  wire _add_map_x_201_wall_t_in;
  wire [9:0] _add_map_x_201_moto;
  wire [9:0] _add_map_x_201_up;
  wire [9:0] _add_map_x_201_right;
  wire [9:0] _add_map_x_201_down;
  wire [9:0] _add_map_x_201_left;
  wire [9:0] _add_map_x_201_start;
  wire [9:0] _add_map_x_201_goal;
  wire [9:0] _add_map_x_201_now;
  wire [9:0] _add_map_x_201_data_out;
  wire [9:0] _add_map_x_201_data_out_index;
  wire [9:0] _add_map_x_201_data_near;
  wire _add_map_x_201_wall_t_out;
  wire [9:0] _add_map_x_201_data_org;
  wire [9:0] _add_map_x_201_data_org_near;
  wire [1:0] _add_map_x_201_s_g;
  wire [1:0] _add_map_x_201_s_g_near;
  wire _add_map_x_201_add_exe;
  wire _add_map_x_201_p_reset;
  wire _add_map_x_201_m_clock;
  wire [9:0] _add_map_x_200_moto_org_near;
  wire [9:0] _add_map_x_200_moto_org_near1;
  wire [9:0] _add_map_x_200_moto_org_near2;
  wire [9:0] _add_map_x_200_moto_org_near3;
  wire [9:0] _add_map_x_200_moto_org;
  wire [1:0] _add_map_x_200_sg_up;
  wire [1:0] _add_map_x_200_sg_down;
  wire [1:0] _add_map_x_200_sg_left;
  wire [1:0] _add_map_x_200_sg_right;
  wire _add_map_x_200_wall_t_in;
  wire [9:0] _add_map_x_200_moto;
  wire [9:0] _add_map_x_200_up;
  wire [9:0] _add_map_x_200_right;
  wire [9:0] _add_map_x_200_down;
  wire [9:0] _add_map_x_200_left;
  wire [9:0] _add_map_x_200_start;
  wire [9:0] _add_map_x_200_goal;
  wire [9:0] _add_map_x_200_now;
  wire [9:0] _add_map_x_200_data_out;
  wire [9:0] _add_map_x_200_data_out_index;
  wire [9:0] _add_map_x_200_data_near;
  wire _add_map_x_200_wall_t_out;
  wire [9:0] _add_map_x_200_data_org;
  wire [9:0] _add_map_x_200_data_org_near;
  wire [1:0] _add_map_x_200_s_g;
  wire [1:0] _add_map_x_200_s_g_near;
  wire _add_map_x_200_add_exe;
  wire _add_map_x_200_p_reset;
  wire _add_map_x_200_m_clock;
  wire [9:0] _add_map_x_199_moto_org_near;
  wire [9:0] _add_map_x_199_moto_org_near1;
  wire [9:0] _add_map_x_199_moto_org_near2;
  wire [9:0] _add_map_x_199_moto_org_near3;
  wire [9:0] _add_map_x_199_moto_org;
  wire [1:0] _add_map_x_199_sg_up;
  wire [1:0] _add_map_x_199_sg_down;
  wire [1:0] _add_map_x_199_sg_left;
  wire [1:0] _add_map_x_199_sg_right;
  wire _add_map_x_199_wall_t_in;
  wire [9:0] _add_map_x_199_moto;
  wire [9:0] _add_map_x_199_up;
  wire [9:0] _add_map_x_199_right;
  wire [9:0] _add_map_x_199_down;
  wire [9:0] _add_map_x_199_left;
  wire [9:0] _add_map_x_199_start;
  wire [9:0] _add_map_x_199_goal;
  wire [9:0] _add_map_x_199_now;
  wire [9:0] _add_map_x_199_data_out;
  wire [9:0] _add_map_x_199_data_out_index;
  wire [9:0] _add_map_x_199_data_near;
  wire _add_map_x_199_wall_t_out;
  wire [9:0] _add_map_x_199_data_org;
  wire [9:0] _add_map_x_199_data_org_near;
  wire [1:0] _add_map_x_199_s_g;
  wire [1:0] _add_map_x_199_s_g_near;
  wire _add_map_x_199_add_exe;
  wire _add_map_x_199_p_reset;
  wire _add_map_x_199_m_clock;
  wire [9:0] _add_map_x_198_moto_org_near;
  wire [9:0] _add_map_x_198_moto_org_near1;
  wire [9:0] _add_map_x_198_moto_org_near2;
  wire [9:0] _add_map_x_198_moto_org_near3;
  wire [9:0] _add_map_x_198_moto_org;
  wire [1:0] _add_map_x_198_sg_up;
  wire [1:0] _add_map_x_198_sg_down;
  wire [1:0] _add_map_x_198_sg_left;
  wire [1:0] _add_map_x_198_sg_right;
  wire _add_map_x_198_wall_t_in;
  wire [9:0] _add_map_x_198_moto;
  wire [9:0] _add_map_x_198_up;
  wire [9:0] _add_map_x_198_right;
  wire [9:0] _add_map_x_198_down;
  wire [9:0] _add_map_x_198_left;
  wire [9:0] _add_map_x_198_start;
  wire [9:0] _add_map_x_198_goal;
  wire [9:0] _add_map_x_198_now;
  wire [9:0] _add_map_x_198_data_out;
  wire [9:0] _add_map_x_198_data_out_index;
  wire [9:0] _add_map_x_198_data_near;
  wire _add_map_x_198_wall_t_out;
  wire [9:0] _add_map_x_198_data_org;
  wire [9:0] _add_map_x_198_data_org_near;
  wire [1:0] _add_map_x_198_s_g;
  wire [1:0] _add_map_x_198_s_g_near;
  wire _add_map_x_198_add_exe;
  wire _add_map_x_198_p_reset;
  wire _add_map_x_198_m_clock;
  wire [9:0] _add_map_x_197_moto_org_near;
  wire [9:0] _add_map_x_197_moto_org_near1;
  wire [9:0] _add_map_x_197_moto_org_near2;
  wire [9:0] _add_map_x_197_moto_org_near3;
  wire [9:0] _add_map_x_197_moto_org;
  wire [1:0] _add_map_x_197_sg_up;
  wire [1:0] _add_map_x_197_sg_down;
  wire [1:0] _add_map_x_197_sg_left;
  wire [1:0] _add_map_x_197_sg_right;
  wire _add_map_x_197_wall_t_in;
  wire [9:0] _add_map_x_197_moto;
  wire [9:0] _add_map_x_197_up;
  wire [9:0] _add_map_x_197_right;
  wire [9:0] _add_map_x_197_down;
  wire [9:0] _add_map_x_197_left;
  wire [9:0] _add_map_x_197_start;
  wire [9:0] _add_map_x_197_goal;
  wire [9:0] _add_map_x_197_now;
  wire [9:0] _add_map_x_197_data_out;
  wire [9:0] _add_map_x_197_data_out_index;
  wire [9:0] _add_map_x_197_data_near;
  wire _add_map_x_197_wall_t_out;
  wire [9:0] _add_map_x_197_data_org;
  wire [9:0] _add_map_x_197_data_org_near;
  wire [1:0] _add_map_x_197_s_g;
  wire [1:0] _add_map_x_197_s_g_near;
  wire _add_map_x_197_add_exe;
  wire _add_map_x_197_p_reset;
  wire _add_map_x_197_m_clock;
  wire [9:0] _add_map_x_196_moto_org_near;
  wire [9:0] _add_map_x_196_moto_org_near1;
  wire [9:0] _add_map_x_196_moto_org_near2;
  wire [9:0] _add_map_x_196_moto_org_near3;
  wire [9:0] _add_map_x_196_moto_org;
  wire [1:0] _add_map_x_196_sg_up;
  wire [1:0] _add_map_x_196_sg_down;
  wire [1:0] _add_map_x_196_sg_left;
  wire [1:0] _add_map_x_196_sg_right;
  wire _add_map_x_196_wall_t_in;
  wire [9:0] _add_map_x_196_moto;
  wire [9:0] _add_map_x_196_up;
  wire [9:0] _add_map_x_196_right;
  wire [9:0] _add_map_x_196_down;
  wire [9:0] _add_map_x_196_left;
  wire [9:0] _add_map_x_196_start;
  wire [9:0] _add_map_x_196_goal;
  wire [9:0] _add_map_x_196_now;
  wire [9:0] _add_map_x_196_data_out;
  wire [9:0] _add_map_x_196_data_out_index;
  wire [9:0] _add_map_x_196_data_near;
  wire _add_map_x_196_wall_t_out;
  wire [9:0] _add_map_x_196_data_org;
  wire [9:0] _add_map_x_196_data_org_near;
  wire [1:0] _add_map_x_196_s_g;
  wire [1:0] _add_map_x_196_s_g_near;
  wire _add_map_x_196_add_exe;
  wire _add_map_x_196_p_reset;
  wire _add_map_x_196_m_clock;
  wire [9:0] _add_map_x_195_moto_org_near;
  wire [9:0] _add_map_x_195_moto_org_near1;
  wire [9:0] _add_map_x_195_moto_org_near2;
  wire [9:0] _add_map_x_195_moto_org_near3;
  wire [9:0] _add_map_x_195_moto_org;
  wire [1:0] _add_map_x_195_sg_up;
  wire [1:0] _add_map_x_195_sg_down;
  wire [1:0] _add_map_x_195_sg_left;
  wire [1:0] _add_map_x_195_sg_right;
  wire _add_map_x_195_wall_t_in;
  wire [9:0] _add_map_x_195_moto;
  wire [9:0] _add_map_x_195_up;
  wire [9:0] _add_map_x_195_right;
  wire [9:0] _add_map_x_195_down;
  wire [9:0] _add_map_x_195_left;
  wire [9:0] _add_map_x_195_start;
  wire [9:0] _add_map_x_195_goal;
  wire [9:0] _add_map_x_195_now;
  wire [9:0] _add_map_x_195_data_out;
  wire [9:0] _add_map_x_195_data_out_index;
  wire [9:0] _add_map_x_195_data_near;
  wire _add_map_x_195_wall_t_out;
  wire [9:0] _add_map_x_195_data_org;
  wire [9:0] _add_map_x_195_data_org_near;
  wire [1:0] _add_map_x_195_s_g;
  wire [1:0] _add_map_x_195_s_g_near;
  wire _add_map_x_195_add_exe;
  wire _add_map_x_195_p_reset;
  wire _add_map_x_195_m_clock;
  wire [9:0] _add_map_x_194_moto_org_near;
  wire [9:0] _add_map_x_194_moto_org_near1;
  wire [9:0] _add_map_x_194_moto_org_near2;
  wire [9:0] _add_map_x_194_moto_org_near3;
  wire [9:0] _add_map_x_194_moto_org;
  wire [1:0] _add_map_x_194_sg_up;
  wire [1:0] _add_map_x_194_sg_down;
  wire [1:0] _add_map_x_194_sg_left;
  wire [1:0] _add_map_x_194_sg_right;
  wire _add_map_x_194_wall_t_in;
  wire [9:0] _add_map_x_194_moto;
  wire [9:0] _add_map_x_194_up;
  wire [9:0] _add_map_x_194_right;
  wire [9:0] _add_map_x_194_down;
  wire [9:0] _add_map_x_194_left;
  wire [9:0] _add_map_x_194_start;
  wire [9:0] _add_map_x_194_goal;
  wire [9:0] _add_map_x_194_now;
  wire [9:0] _add_map_x_194_data_out;
  wire [9:0] _add_map_x_194_data_out_index;
  wire [9:0] _add_map_x_194_data_near;
  wire _add_map_x_194_wall_t_out;
  wire [9:0] _add_map_x_194_data_org;
  wire [9:0] _add_map_x_194_data_org_near;
  wire [1:0] _add_map_x_194_s_g;
  wire [1:0] _add_map_x_194_s_g_near;
  wire _add_map_x_194_add_exe;
  wire _add_map_x_194_p_reset;
  wire _add_map_x_194_m_clock;
  wire [9:0] _add_map_x_193_moto_org_near;
  wire [9:0] _add_map_x_193_moto_org_near1;
  wire [9:0] _add_map_x_193_moto_org_near2;
  wire [9:0] _add_map_x_193_moto_org_near3;
  wire [9:0] _add_map_x_193_moto_org;
  wire [1:0] _add_map_x_193_sg_up;
  wire [1:0] _add_map_x_193_sg_down;
  wire [1:0] _add_map_x_193_sg_left;
  wire [1:0] _add_map_x_193_sg_right;
  wire _add_map_x_193_wall_t_in;
  wire [9:0] _add_map_x_193_moto;
  wire [9:0] _add_map_x_193_up;
  wire [9:0] _add_map_x_193_right;
  wire [9:0] _add_map_x_193_down;
  wire [9:0] _add_map_x_193_left;
  wire [9:0] _add_map_x_193_start;
  wire [9:0] _add_map_x_193_goal;
  wire [9:0] _add_map_x_193_now;
  wire [9:0] _add_map_x_193_data_out;
  wire [9:0] _add_map_x_193_data_out_index;
  wire [9:0] _add_map_x_193_data_near;
  wire _add_map_x_193_wall_t_out;
  wire [9:0] _add_map_x_193_data_org;
  wire [9:0] _add_map_x_193_data_org_near;
  wire [1:0] _add_map_x_193_s_g;
  wire [1:0] _add_map_x_193_s_g_near;
  wire _add_map_x_193_add_exe;
  wire _add_map_x_193_p_reset;
  wire _add_map_x_193_m_clock;
  wire [9:0] _add_map_x_192_moto_org_near;
  wire [9:0] _add_map_x_192_moto_org_near1;
  wire [9:0] _add_map_x_192_moto_org_near2;
  wire [9:0] _add_map_x_192_moto_org_near3;
  wire [9:0] _add_map_x_192_moto_org;
  wire [1:0] _add_map_x_192_sg_up;
  wire [1:0] _add_map_x_192_sg_down;
  wire [1:0] _add_map_x_192_sg_left;
  wire [1:0] _add_map_x_192_sg_right;
  wire _add_map_x_192_wall_t_in;
  wire [9:0] _add_map_x_192_moto;
  wire [9:0] _add_map_x_192_up;
  wire [9:0] _add_map_x_192_right;
  wire [9:0] _add_map_x_192_down;
  wire [9:0] _add_map_x_192_left;
  wire [9:0] _add_map_x_192_start;
  wire [9:0] _add_map_x_192_goal;
  wire [9:0] _add_map_x_192_now;
  wire [9:0] _add_map_x_192_data_out;
  wire [9:0] _add_map_x_192_data_out_index;
  wire [9:0] _add_map_x_192_data_near;
  wire _add_map_x_192_wall_t_out;
  wire [9:0] _add_map_x_192_data_org;
  wire [9:0] _add_map_x_192_data_org_near;
  wire [1:0] _add_map_x_192_s_g;
  wire [1:0] _add_map_x_192_s_g_near;
  wire _add_map_x_192_add_exe;
  wire _add_map_x_192_p_reset;
  wire _add_map_x_192_m_clock;
  wire [9:0] _add_map_x_191_moto_org_near;
  wire [9:0] _add_map_x_191_moto_org_near1;
  wire [9:0] _add_map_x_191_moto_org_near2;
  wire [9:0] _add_map_x_191_moto_org_near3;
  wire [9:0] _add_map_x_191_moto_org;
  wire [1:0] _add_map_x_191_sg_up;
  wire [1:0] _add_map_x_191_sg_down;
  wire [1:0] _add_map_x_191_sg_left;
  wire [1:0] _add_map_x_191_sg_right;
  wire _add_map_x_191_wall_t_in;
  wire [9:0] _add_map_x_191_moto;
  wire [9:0] _add_map_x_191_up;
  wire [9:0] _add_map_x_191_right;
  wire [9:0] _add_map_x_191_down;
  wire [9:0] _add_map_x_191_left;
  wire [9:0] _add_map_x_191_start;
  wire [9:0] _add_map_x_191_goal;
  wire [9:0] _add_map_x_191_now;
  wire [9:0] _add_map_x_191_data_out;
  wire [9:0] _add_map_x_191_data_out_index;
  wire [9:0] _add_map_x_191_data_near;
  wire _add_map_x_191_wall_t_out;
  wire [9:0] _add_map_x_191_data_org;
  wire [9:0] _add_map_x_191_data_org_near;
  wire [1:0] _add_map_x_191_s_g;
  wire [1:0] _add_map_x_191_s_g_near;
  wire _add_map_x_191_add_exe;
  wire _add_map_x_191_p_reset;
  wire _add_map_x_191_m_clock;
  wire [9:0] _add_map_x_190_moto_org_near;
  wire [9:0] _add_map_x_190_moto_org_near1;
  wire [9:0] _add_map_x_190_moto_org_near2;
  wire [9:0] _add_map_x_190_moto_org_near3;
  wire [9:0] _add_map_x_190_moto_org;
  wire [1:0] _add_map_x_190_sg_up;
  wire [1:0] _add_map_x_190_sg_down;
  wire [1:0] _add_map_x_190_sg_left;
  wire [1:0] _add_map_x_190_sg_right;
  wire _add_map_x_190_wall_t_in;
  wire [9:0] _add_map_x_190_moto;
  wire [9:0] _add_map_x_190_up;
  wire [9:0] _add_map_x_190_right;
  wire [9:0] _add_map_x_190_down;
  wire [9:0] _add_map_x_190_left;
  wire [9:0] _add_map_x_190_start;
  wire [9:0] _add_map_x_190_goal;
  wire [9:0] _add_map_x_190_now;
  wire [9:0] _add_map_x_190_data_out;
  wire [9:0] _add_map_x_190_data_out_index;
  wire [9:0] _add_map_x_190_data_near;
  wire _add_map_x_190_wall_t_out;
  wire [9:0] _add_map_x_190_data_org;
  wire [9:0] _add_map_x_190_data_org_near;
  wire [1:0] _add_map_x_190_s_g;
  wire [1:0] _add_map_x_190_s_g_near;
  wire _add_map_x_190_add_exe;
  wire _add_map_x_190_p_reset;
  wire _add_map_x_190_m_clock;
  wire [9:0] _add_map_x_189_moto_org_near;
  wire [9:0] _add_map_x_189_moto_org_near1;
  wire [9:0] _add_map_x_189_moto_org_near2;
  wire [9:0] _add_map_x_189_moto_org_near3;
  wire [9:0] _add_map_x_189_moto_org;
  wire [1:0] _add_map_x_189_sg_up;
  wire [1:0] _add_map_x_189_sg_down;
  wire [1:0] _add_map_x_189_sg_left;
  wire [1:0] _add_map_x_189_sg_right;
  wire _add_map_x_189_wall_t_in;
  wire [9:0] _add_map_x_189_moto;
  wire [9:0] _add_map_x_189_up;
  wire [9:0] _add_map_x_189_right;
  wire [9:0] _add_map_x_189_down;
  wire [9:0] _add_map_x_189_left;
  wire [9:0] _add_map_x_189_start;
  wire [9:0] _add_map_x_189_goal;
  wire [9:0] _add_map_x_189_now;
  wire [9:0] _add_map_x_189_data_out;
  wire [9:0] _add_map_x_189_data_out_index;
  wire [9:0] _add_map_x_189_data_near;
  wire _add_map_x_189_wall_t_out;
  wire [9:0] _add_map_x_189_data_org;
  wire [9:0] _add_map_x_189_data_org_near;
  wire [1:0] _add_map_x_189_s_g;
  wire [1:0] _add_map_x_189_s_g_near;
  wire _add_map_x_189_add_exe;
  wire _add_map_x_189_p_reset;
  wire _add_map_x_189_m_clock;
  wire [9:0] _add_map_x_188_moto_org_near;
  wire [9:0] _add_map_x_188_moto_org_near1;
  wire [9:0] _add_map_x_188_moto_org_near2;
  wire [9:0] _add_map_x_188_moto_org_near3;
  wire [9:0] _add_map_x_188_moto_org;
  wire [1:0] _add_map_x_188_sg_up;
  wire [1:0] _add_map_x_188_sg_down;
  wire [1:0] _add_map_x_188_sg_left;
  wire [1:0] _add_map_x_188_sg_right;
  wire _add_map_x_188_wall_t_in;
  wire [9:0] _add_map_x_188_moto;
  wire [9:0] _add_map_x_188_up;
  wire [9:0] _add_map_x_188_right;
  wire [9:0] _add_map_x_188_down;
  wire [9:0] _add_map_x_188_left;
  wire [9:0] _add_map_x_188_start;
  wire [9:0] _add_map_x_188_goal;
  wire [9:0] _add_map_x_188_now;
  wire [9:0] _add_map_x_188_data_out;
  wire [9:0] _add_map_x_188_data_out_index;
  wire [9:0] _add_map_x_188_data_near;
  wire _add_map_x_188_wall_t_out;
  wire [9:0] _add_map_x_188_data_org;
  wire [9:0] _add_map_x_188_data_org_near;
  wire [1:0] _add_map_x_188_s_g;
  wire [1:0] _add_map_x_188_s_g_near;
  wire _add_map_x_188_add_exe;
  wire _add_map_x_188_p_reset;
  wire _add_map_x_188_m_clock;
  wire [9:0] _add_map_x_187_moto_org_near;
  wire [9:0] _add_map_x_187_moto_org_near1;
  wire [9:0] _add_map_x_187_moto_org_near2;
  wire [9:0] _add_map_x_187_moto_org_near3;
  wire [9:0] _add_map_x_187_moto_org;
  wire [1:0] _add_map_x_187_sg_up;
  wire [1:0] _add_map_x_187_sg_down;
  wire [1:0] _add_map_x_187_sg_left;
  wire [1:0] _add_map_x_187_sg_right;
  wire _add_map_x_187_wall_t_in;
  wire [9:0] _add_map_x_187_moto;
  wire [9:0] _add_map_x_187_up;
  wire [9:0] _add_map_x_187_right;
  wire [9:0] _add_map_x_187_down;
  wire [9:0] _add_map_x_187_left;
  wire [9:0] _add_map_x_187_start;
  wire [9:0] _add_map_x_187_goal;
  wire [9:0] _add_map_x_187_now;
  wire [9:0] _add_map_x_187_data_out;
  wire [9:0] _add_map_x_187_data_out_index;
  wire [9:0] _add_map_x_187_data_near;
  wire _add_map_x_187_wall_t_out;
  wire [9:0] _add_map_x_187_data_org;
  wire [9:0] _add_map_x_187_data_org_near;
  wire [1:0] _add_map_x_187_s_g;
  wire [1:0] _add_map_x_187_s_g_near;
  wire _add_map_x_187_add_exe;
  wire _add_map_x_187_p_reset;
  wire _add_map_x_187_m_clock;
  wire [9:0] _add_map_x_186_moto_org_near;
  wire [9:0] _add_map_x_186_moto_org_near1;
  wire [9:0] _add_map_x_186_moto_org_near2;
  wire [9:0] _add_map_x_186_moto_org_near3;
  wire [9:0] _add_map_x_186_moto_org;
  wire [1:0] _add_map_x_186_sg_up;
  wire [1:0] _add_map_x_186_sg_down;
  wire [1:0] _add_map_x_186_sg_left;
  wire [1:0] _add_map_x_186_sg_right;
  wire _add_map_x_186_wall_t_in;
  wire [9:0] _add_map_x_186_moto;
  wire [9:0] _add_map_x_186_up;
  wire [9:0] _add_map_x_186_right;
  wire [9:0] _add_map_x_186_down;
  wire [9:0] _add_map_x_186_left;
  wire [9:0] _add_map_x_186_start;
  wire [9:0] _add_map_x_186_goal;
  wire [9:0] _add_map_x_186_now;
  wire [9:0] _add_map_x_186_data_out;
  wire [9:0] _add_map_x_186_data_out_index;
  wire [9:0] _add_map_x_186_data_near;
  wire _add_map_x_186_wall_t_out;
  wire [9:0] _add_map_x_186_data_org;
  wire [9:0] _add_map_x_186_data_org_near;
  wire [1:0] _add_map_x_186_s_g;
  wire [1:0] _add_map_x_186_s_g_near;
  wire _add_map_x_186_add_exe;
  wire _add_map_x_186_p_reset;
  wire _add_map_x_186_m_clock;
  wire [9:0] _add_map_x_185_moto_org_near;
  wire [9:0] _add_map_x_185_moto_org_near1;
  wire [9:0] _add_map_x_185_moto_org_near2;
  wire [9:0] _add_map_x_185_moto_org_near3;
  wire [9:0] _add_map_x_185_moto_org;
  wire [1:0] _add_map_x_185_sg_up;
  wire [1:0] _add_map_x_185_sg_down;
  wire [1:0] _add_map_x_185_sg_left;
  wire [1:0] _add_map_x_185_sg_right;
  wire _add_map_x_185_wall_t_in;
  wire [9:0] _add_map_x_185_moto;
  wire [9:0] _add_map_x_185_up;
  wire [9:0] _add_map_x_185_right;
  wire [9:0] _add_map_x_185_down;
  wire [9:0] _add_map_x_185_left;
  wire [9:0] _add_map_x_185_start;
  wire [9:0] _add_map_x_185_goal;
  wire [9:0] _add_map_x_185_now;
  wire [9:0] _add_map_x_185_data_out;
  wire [9:0] _add_map_x_185_data_out_index;
  wire [9:0] _add_map_x_185_data_near;
  wire _add_map_x_185_wall_t_out;
  wire [9:0] _add_map_x_185_data_org;
  wire [9:0] _add_map_x_185_data_org_near;
  wire [1:0] _add_map_x_185_s_g;
  wire [1:0] _add_map_x_185_s_g_near;
  wire _add_map_x_185_add_exe;
  wire _add_map_x_185_p_reset;
  wire _add_map_x_185_m_clock;
  wire [9:0] _add_map_x_184_moto_org_near;
  wire [9:0] _add_map_x_184_moto_org_near1;
  wire [9:0] _add_map_x_184_moto_org_near2;
  wire [9:0] _add_map_x_184_moto_org_near3;
  wire [9:0] _add_map_x_184_moto_org;
  wire [1:0] _add_map_x_184_sg_up;
  wire [1:0] _add_map_x_184_sg_down;
  wire [1:0] _add_map_x_184_sg_left;
  wire [1:0] _add_map_x_184_sg_right;
  wire _add_map_x_184_wall_t_in;
  wire [9:0] _add_map_x_184_moto;
  wire [9:0] _add_map_x_184_up;
  wire [9:0] _add_map_x_184_right;
  wire [9:0] _add_map_x_184_down;
  wire [9:0] _add_map_x_184_left;
  wire [9:0] _add_map_x_184_start;
  wire [9:0] _add_map_x_184_goal;
  wire [9:0] _add_map_x_184_now;
  wire [9:0] _add_map_x_184_data_out;
  wire [9:0] _add_map_x_184_data_out_index;
  wire [9:0] _add_map_x_184_data_near;
  wire _add_map_x_184_wall_t_out;
  wire [9:0] _add_map_x_184_data_org;
  wire [9:0] _add_map_x_184_data_org_near;
  wire [1:0] _add_map_x_184_s_g;
  wire [1:0] _add_map_x_184_s_g_near;
  wire _add_map_x_184_add_exe;
  wire _add_map_x_184_p_reset;
  wire _add_map_x_184_m_clock;
  wire [9:0] _add_map_x_183_moto_org_near;
  wire [9:0] _add_map_x_183_moto_org_near1;
  wire [9:0] _add_map_x_183_moto_org_near2;
  wire [9:0] _add_map_x_183_moto_org_near3;
  wire [9:0] _add_map_x_183_moto_org;
  wire [1:0] _add_map_x_183_sg_up;
  wire [1:0] _add_map_x_183_sg_down;
  wire [1:0] _add_map_x_183_sg_left;
  wire [1:0] _add_map_x_183_sg_right;
  wire _add_map_x_183_wall_t_in;
  wire [9:0] _add_map_x_183_moto;
  wire [9:0] _add_map_x_183_up;
  wire [9:0] _add_map_x_183_right;
  wire [9:0] _add_map_x_183_down;
  wire [9:0] _add_map_x_183_left;
  wire [9:0] _add_map_x_183_start;
  wire [9:0] _add_map_x_183_goal;
  wire [9:0] _add_map_x_183_now;
  wire [9:0] _add_map_x_183_data_out;
  wire [9:0] _add_map_x_183_data_out_index;
  wire [9:0] _add_map_x_183_data_near;
  wire _add_map_x_183_wall_t_out;
  wire [9:0] _add_map_x_183_data_org;
  wire [9:0] _add_map_x_183_data_org_near;
  wire [1:0] _add_map_x_183_s_g;
  wire [1:0] _add_map_x_183_s_g_near;
  wire _add_map_x_183_add_exe;
  wire _add_map_x_183_p_reset;
  wire _add_map_x_183_m_clock;
  wire [9:0] _add_map_x_182_moto_org_near;
  wire [9:0] _add_map_x_182_moto_org_near1;
  wire [9:0] _add_map_x_182_moto_org_near2;
  wire [9:0] _add_map_x_182_moto_org_near3;
  wire [9:0] _add_map_x_182_moto_org;
  wire [1:0] _add_map_x_182_sg_up;
  wire [1:0] _add_map_x_182_sg_down;
  wire [1:0] _add_map_x_182_sg_left;
  wire [1:0] _add_map_x_182_sg_right;
  wire _add_map_x_182_wall_t_in;
  wire [9:0] _add_map_x_182_moto;
  wire [9:0] _add_map_x_182_up;
  wire [9:0] _add_map_x_182_right;
  wire [9:0] _add_map_x_182_down;
  wire [9:0] _add_map_x_182_left;
  wire [9:0] _add_map_x_182_start;
  wire [9:0] _add_map_x_182_goal;
  wire [9:0] _add_map_x_182_now;
  wire [9:0] _add_map_x_182_data_out;
  wire [9:0] _add_map_x_182_data_out_index;
  wire [9:0] _add_map_x_182_data_near;
  wire _add_map_x_182_wall_t_out;
  wire [9:0] _add_map_x_182_data_org;
  wire [9:0] _add_map_x_182_data_org_near;
  wire [1:0] _add_map_x_182_s_g;
  wire [1:0] _add_map_x_182_s_g_near;
  wire _add_map_x_182_add_exe;
  wire _add_map_x_182_p_reset;
  wire _add_map_x_182_m_clock;
  wire [9:0] _add_map_x_181_moto_org_near;
  wire [9:0] _add_map_x_181_moto_org_near1;
  wire [9:0] _add_map_x_181_moto_org_near2;
  wire [9:0] _add_map_x_181_moto_org_near3;
  wire [9:0] _add_map_x_181_moto_org;
  wire [1:0] _add_map_x_181_sg_up;
  wire [1:0] _add_map_x_181_sg_down;
  wire [1:0] _add_map_x_181_sg_left;
  wire [1:0] _add_map_x_181_sg_right;
  wire _add_map_x_181_wall_t_in;
  wire [9:0] _add_map_x_181_moto;
  wire [9:0] _add_map_x_181_up;
  wire [9:0] _add_map_x_181_right;
  wire [9:0] _add_map_x_181_down;
  wire [9:0] _add_map_x_181_left;
  wire [9:0] _add_map_x_181_start;
  wire [9:0] _add_map_x_181_goal;
  wire [9:0] _add_map_x_181_now;
  wire [9:0] _add_map_x_181_data_out;
  wire [9:0] _add_map_x_181_data_out_index;
  wire [9:0] _add_map_x_181_data_near;
  wire _add_map_x_181_wall_t_out;
  wire [9:0] _add_map_x_181_data_org;
  wire [9:0] _add_map_x_181_data_org_near;
  wire [1:0] _add_map_x_181_s_g;
  wire [1:0] _add_map_x_181_s_g_near;
  wire _add_map_x_181_add_exe;
  wire _add_map_x_181_p_reset;
  wire _add_map_x_181_m_clock;
  wire [9:0] _add_map_x_180_moto_org_near;
  wire [9:0] _add_map_x_180_moto_org_near1;
  wire [9:0] _add_map_x_180_moto_org_near2;
  wire [9:0] _add_map_x_180_moto_org_near3;
  wire [9:0] _add_map_x_180_moto_org;
  wire [1:0] _add_map_x_180_sg_up;
  wire [1:0] _add_map_x_180_sg_down;
  wire [1:0] _add_map_x_180_sg_left;
  wire [1:0] _add_map_x_180_sg_right;
  wire _add_map_x_180_wall_t_in;
  wire [9:0] _add_map_x_180_moto;
  wire [9:0] _add_map_x_180_up;
  wire [9:0] _add_map_x_180_right;
  wire [9:0] _add_map_x_180_down;
  wire [9:0] _add_map_x_180_left;
  wire [9:0] _add_map_x_180_start;
  wire [9:0] _add_map_x_180_goal;
  wire [9:0] _add_map_x_180_now;
  wire [9:0] _add_map_x_180_data_out;
  wire [9:0] _add_map_x_180_data_out_index;
  wire [9:0] _add_map_x_180_data_near;
  wire _add_map_x_180_wall_t_out;
  wire [9:0] _add_map_x_180_data_org;
  wire [9:0] _add_map_x_180_data_org_near;
  wire [1:0] _add_map_x_180_s_g;
  wire [1:0] _add_map_x_180_s_g_near;
  wire _add_map_x_180_add_exe;
  wire _add_map_x_180_p_reset;
  wire _add_map_x_180_m_clock;
  wire [9:0] _add_map_x_179_moto_org_near;
  wire [9:0] _add_map_x_179_moto_org_near1;
  wire [9:0] _add_map_x_179_moto_org_near2;
  wire [9:0] _add_map_x_179_moto_org_near3;
  wire [9:0] _add_map_x_179_moto_org;
  wire [1:0] _add_map_x_179_sg_up;
  wire [1:0] _add_map_x_179_sg_down;
  wire [1:0] _add_map_x_179_sg_left;
  wire [1:0] _add_map_x_179_sg_right;
  wire _add_map_x_179_wall_t_in;
  wire [9:0] _add_map_x_179_moto;
  wire [9:0] _add_map_x_179_up;
  wire [9:0] _add_map_x_179_right;
  wire [9:0] _add_map_x_179_down;
  wire [9:0] _add_map_x_179_left;
  wire [9:0] _add_map_x_179_start;
  wire [9:0] _add_map_x_179_goal;
  wire [9:0] _add_map_x_179_now;
  wire [9:0] _add_map_x_179_data_out;
  wire [9:0] _add_map_x_179_data_out_index;
  wire [9:0] _add_map_x_179_data_near;
  wire _add_map_x_179_wall_t_out;
  wire [9:0] _add_map_x_179_data_org;
  wire [9:0] _add_map_x_179_data_org_near;
  wire [1:0] _add_map_x_179_s_g;
  wire [1:0] _add_map_x_179_s_g_near;
  wire _add_map_x_179_add_exe;
  wire _add_map_x_179_p_reset;
  wire _add_map_x_179_m_clock;
  wire [9:0] _add_map_x_178_moto_org_near;
  wire [9:0] _add_map_x_178_moto_org_near1;
  wire [9:0] _add_map_x_178_moto_org_near2;
  wire [9:0] _add_map_x_178_moto_org_near3;
  wire [9:0] _add_map_x_178_moto_org;
  wire [1:0] _add_map_x_178_sg_up;
  wire [1:0] _add_map_x_178_sg_down;
  wire [1:0] _add_map_x_178_sg_left;
  wire [1:0] _add_map_x_178_sg_right;
  wire _add_map_x_178_wall_t_in;
  wire [9:0] _add_map_x_178_moto;
  wire [9:0] _add_map_x_178_up;
  wire [9:0] _add_map_x_178_right;
  wire [9:0] _add_map_x_178_down;
  wire [9:0] _add_map_x_178_left;
  wire [9:0] _add_map_x_178_start;
  wire [9:0] _add_map_x_178_goal;
  wire [9:0] _add_map_x_178_now;
  wire [9:0] _add_map_x_178_data_out;
  wire [9:0] _add_map_x_178_data_out_index;
  wire [9:0] _add_map_x_178_data_near;
  wire _add_map_x_178_wall_t_out;
  wire [9:0] _add_map_x_178_data_org;
  wire [9:0] _add_map_x_178_data_org_near;
  wire [1:0] _add_map_x_178_s_g;
  wire [1:0] _add_map_x_178_s_g_near;
  wire _add_map_x_178_add_exe;
  wire _add_map_x_178_p_reset;
  wire _add_map_x_178_m_clock;
  wire [9:0] _add_map_x_177_moto_org_near;
  wire [9:0] _add_map_x_177_moto_org_near1;
  wire [9:0] _add_map_x_177_moto_org_near2;
  wire [9:0] _add_map_x_177_moto_org_near3;
  wire [9:0] _add_map_x_177_moto_org;
  wire [1:0] _add_map_x_177_sg_up;
  wire [1:0] _add_map_x_177_sg_down;
  wire [1:0] _add_map_x_177_sg_left;
  wire [1:0] _add_map_x_177_sg_right;
  wire _add_map_x_177_wall_t_in;
  wire [9:0] _add_map_x_177_moto;
  wire [9:0] _add_map_x_177_up;
  wire [9:0] _add_map_x_177_right;
  wire [9:0] _add_map_x_177_down;
  wire [9:0] _add_map_x_177_left;
  wire [9:0] _add_map_x_177_start;
  wire [9:0] _add_map_x_177_goal;
  wire [9:0] _add_map_x_177_now;
  wire [9:0] _add_map_x_177_data_out;
  wire [9:0] _add_map_x_177_data_out_index;
  wire [9:0] _add_map_x_177_data_near;
  wire _add_map_x_177_wall_t_out;
  wire [9:0] _add_map_x_177_data_org;
  wire [9:0] _add_map_x_177_data_org_near;
  wire [1:0] _add_map_x_177_s_g;
  wire [1:0] _add_map_x_177_s_g_near;
  wire _add_map_x_177_add_exe;
  wire _add_map_x_177_p_reset;
  wire _add_map_x_177_m_clock;
  wire [9:0] _add_map_x_176_moto_org_near;
  wire [9:0] _add_map_x_176_moto_org_near1;
  wire [9:0] _add_map_x_176_moto_org_near2;
  wire [9:0] _add_map_x_176_moto_org_near3;
  wire [9:0] _add_map_x_176_moto_org;
  wire [1:0] _add_map_x_176_sg_up;
  wire [1:0] _add_map_x_176_sg_down;
  wire [1:0] _add_map_x_176_sg_left;
  wire [1:0] _add_map_x_176_sg_right;
  wire _add_map_x_176_wall_t_in;
  wire [9:0] _add_map_x_176_moto;
  wire [9:0] _add_map_x_176_up;
  wire [9:0] _add_map_x_176_right;
  wire [9:0] _add_map_x_176_down;
  wire [9:0] _add_map_x_176_left;
  wire [9:0] _add_map_x_176_start;
  wire [9:0] _add_map_x_176_goal;
  wire [9:0] _add_map_x_176_now;
  wire [9:0] _add_map_x_176_data_out;
  wire [9:0] _add_map_x_176_data_out_index;
  wire [9:0] _add_map_x_176_data_near;
  wire _add_map_x_176_wall_t_out;
  wire [9:0] _add_map_x_176_data_org;
  wire [9:0] _add_map_x_176_data_org_near;
  wire [1:0] _add_map_x_176_s_g;
  wire [1:0] _add_map_x_176_s_g_near;
  wire _add_map_x_176_add_exe;
  wire _add_map_x_176_p_reset;
  wire _add_map_x_176_m_clock;
  wire [9:0] _add_map_x_175_moto_org_near;
  wire [9:0] _add_map_x_175_moto_org_near1;
  wire [9:0] _add_map_x_175_moto_org_near2;
  wire [9:0] _add_map_x_175_moto_org_near3;
  wire [9:0] _add_map_x_175_moto_org;
  wire [1:0] _add_map_x_175_sg_up;
  wire [1:0] _add_map_x_175_sg_down;
  wire [1:0] _add_map_x_175_sg_left;
  wire [1:0] _add_map_x_175_sg_right;
  wire _add_map_x_175_wall_t_in;
  wire [9:0] _add_map_x_175_moto;
  wire [9:0] _add_map_x_175_up;
  wire [9:0] _add_map_x_175_right;
  wire [9:0] _add_map_x_175_down;
  wire [9:0] _add_map_x_175_left;
  wire [9:0] _add_map_x_175_start;
  wire [9:0] _add_map_x_175_goal;
  wire [9:0] _add_map_x_175_now;
  wire [9:0] _add_map_x_175_data_out;
  wire [9:0] _add_map_x_175_data_out_index;
  wire [9:0] _add_map_x_175_data_near;
  wire _add_map_x_175_wall_t_out;
  wire [9:0] _add_map_x_175_data_org;
  wire [9:0] _add_map_x_175_data_org_near;
  wire [1:0] _add_map_x_175_s_g;
  wire [1:0] _add_map_x_175_s_g_near;
  wire _add_map_x_175_add_exe;
  wire _add_map_x_175_p_reset;
  wire _add_map_x_175_m_clock;
  wire [9:0] _add_map_x_174_moto_org_near;
  wire [9:0] _add_map_x_174_moto_org_near1;
  wire [9:0] _add_map_x_174_moto_org_near2;
  wire [9:0] _add_map_x_174_moto_org_near3;
  wire [9:0] _add_map_x_174_moto_org;
  wire [1:0] _add_map_x_174_sg_up;
  wire [1:0] _add_map_x_174_sg_down;
  wire [1:0] _add_map_x_174_sg_left;
  wire [1:0] _add_map_x_174_sg_right;
  wire _add_map_x_174_wall_t_in;
  wire [9:0] _add_map_x_174_moto;
  wire [9:0] _add_map_x_174_up;
  wire [9:0] _add_map_x_174_right;
  wire [9:0] _add_map_x_174_down;
  wire [9:0] _add_map_x_174_left;
  wire [9:0] _add_map_x_174_start;
  wire [9:0] _add_map_x_174_goal;
  wire [9:0] _add_map_x_174_now;
  wire [9:0] _add_map_x_174_data_out;
  wire [9:0] _add_map_x_174_data_out_index;
  wire [9:0] _add_map_x_174_data_near;
  wire _add_map_x_174_wall_t_out;
  wire [9:0] _add_map_x_174_data_org;
  wire [9:0] _add_map_x_174_data_org_near;
  wire [1:0] _add_map_x_174_s_g;
  wire [1:0] _add_map_x_174_s_g_near;
  wire _add_map_x_174_add_exe;
  wire _add_map_x_174_p_reset;
  wire _add_map_x_174_m_clock;
  wire [9:0] _add_map_x_173_moto_org_near;
  wire [9:0] _add_map_x_173_moto_org_near1;
  wire [9:0] _add_map_x_173_moto_org_near2;
  wire [9:0] _add_map_x_173_moto_org_near3;
  wire [9:0] _add_map_x_173_moto_org;
  wire [1:0] _add_map_x_173_sg_up;
  wire [1:0] _add_map_x_173_sg_down;
  wire [1:0] _add_map_x_173_sg_left;
  wire [1:0] _add_map_x_173_sg_right;
  wire _add_map_x_173_wall_t_in;
  wire [9:0] _add_map_x_173_moto;
  wire [9:0] _add_map_x_173_up;
  wire [9:0] _add_map_x_173_right;
  wire [9:0] _add_map_x_173_down;
  wire [9:0] _add_map_x_173_left;
  wire [9:0] _add_map_x_173_start;
  wire [9:0] _add_map_x_173_goal;
  wire [9:0] _add_map_x_173_now;
  wire [9:0] _add_map_x_173_data_out;
  wire [9:0] _add_map_x_173_data_out_index;
  wire [9:0] _add_map_x_173_data_near;
  wire _add_map_x_173_wall_t_out;
  wire [9:0] _add_map_x_173_data_org;
  wire [9:0] _add_map_x_173_data_org_near;
  wire [1:0] _add_map_x_173_s_g;
  wire [1:0] _add_map_x_173_s_g_near;
  wire _add_map_x_173_add_exe;
  wire _add_map_x_173_p_reset;
  wire _add_map_x_173_m_clock;
  wire [9:0] _add_map_x_172_moto_org_near;
  wire [9:0] _add_map_x_172_moto_org_near1;
  wire [9:0] _add_map_x_172_moto_org_near2;
  wire [9:0] _add_map_x_172_moto_org_near3;
  wire [9:0] _add_map_x_172_moto_org;
  wire [1:0] _add_map_x_172_sg_up;
  wire [1:0] _add_map_x_172_sg_down;
  wire [1:0] _add_map_x_172_sg_left;
  wire [1:0] _add_map_x_172_sg_right;
  wire _add_map_x_172_wall_t_in;
  wire [9:0] _add_map_x_172_moto;
  wire [9:0] _add_map_x_172_up;
  wire [9:0] _add_map_x_172_right;
  wire [9:0] _add_map_x_172_down;
  wire [9:0] _add_map_x_172_left;
  wire [9:0] _add_map_x_172_start;
  wire [9:0] _add_map_x_172_goal;
  wire [9:0] _add_map_x_172_now;
  wire [9:0] _add_map_x_172_data_out;
  wire [9:0] _add_map_x_172_data_out_index;
  wire [9:0] _add_map_x_172_data_near;
  wire _add_map_x_172_wall_t_out;
  wire [9:0] _add_map_x_172_data_org;
  wire [9:0] _add_map_x_172_data_org_near;
  wire [1:0] _add_map_x_172_s_g;
  wire [1:0] _add_map_x_172_s_g_near;
  wire _add_map_x_172_add_exe;
  wire _add_map_x_172_p_reset;
  wire _add_map_x_172_m_clock;
  wire [9:0] _add_map_x_171_moto_org_near;
  wire [9:0] _add_map_x_171_moto_org_near1;
  wire [9:0] _add_map_x_171_moto_org_near2;
  wire [9:0] _add_map_x_171_moto_org_near3;
  wire [9:0] _add_map_x_171_moto_org;
  wire [1:0] _add_map_x_171_sg_up;
  wire [1:0] _add_map_x_171_sg_down;
  wire [1:0] _add_map_x_171_sg_left;
  wire [1:0] _add_map_x_171_sg_right;
  wire _add_map_x_171_wall_t_in;
  wire [9:0] _add_map_x_171_moto;
  wire [9:0] _add_map_x_171_up;
  wire [9:0] _add_map_x_171_right;
  wire [9:0] _add_map_x_171_down;
  wire [9:0] _add_map_x_171_left;
  wire [9:0] _add_map_x_171_start;
  wire [9:0] _add_map_x_171_goal;
  wire [9:0] _add_map_x_171_now;
  wire [9:0] _add_map_x_171_data_out;
  wire [9:0] _add_map_x_171_data_out_index;
  wire [9:0] _add_map_x_171_data_near;
  wire _add_map_x_171_wall_t_out;
  wire [9:0] _add_map_x_171_data_org;
  wire [9:0] _add_map_x_171_data_org_near;
  wire [1:0] _add_map_x_171_s_g;
  wire [1:0] _add_map_x_171_s_g_near;
  wire _add_map_x_171_add_exe;
  wire _add_map_x_171_p_reset;
  wire _add_map_x_171_m_clock;
  wire [9:0] _add_map_x_170_moto_org_near;
  wire [9:0] _add_map_x_170_moto_org_near1;
  wire [9:0] _add_map_x_170_moto_org_near2;
  wire [9:0] _add_map_x_170_moto_org_near3;
  wire [9:0] _add_map_x_170_moto_org;
  wire [1:0] _add_map_x_170_sg_up;
  wire [1:0] _add_map_x_170_sg_down;
  wire [1:0] _add_map_x_170_sg_left;
  wire [1:0] _add_map_x_170_sg_right;
  wire _add_map_x_170_wall_t_in;
  wire [9:0] _add_map_x_170_moto;
  wire [9:0] _add_map_x_170_up;
  wire [9:0] _add_map_x_170_right;
  wire [9:0] _add_map_x_170_down;
  wire [9:0] _add_map_x_170_left;
  wire [9:0] _add_map_x_170_start;
  wire [9:0] _add_map_x_170_goal;
  wire [9:0] _add_map_x_170_now;
  wire [9:0] _add_map_x_170_data_out;
  wire [9:0] _add_map_x_170_data_out_index;
  wire [9:0] _add_map_x_170_data_near;
  wire _add_map_x_170_wall_t_out;
  wire [9:0] _add_map_x_170_data_org;
  wire [9:0] _add_map_x_170_data_org_near;
  wire [1:0] _add_map_x_170_s_g;
  wire [1:0] _add_map_x_170_s_g_near;
  wire _add_map_x_170_add_exe;
  wire _add_map_x_170_p_reset;
  wire _add_map_x_170_m_clock;
  wire [9:0] _add_map_x_169_moto_org_near;
  wire [9:0] _add_map_x_169_moto_org_near1;
  wire [9:0] _add_map_x_169_moto_org_near2;
  wire [9:0] _add_map_x_169_moto_org_near3;
  wire [9:0] _add_map_x_169_moto_org;
  wire [1:0] _add_map_x_169_sg_up;
  wire [1:0] _add_map_x_169_sg_down;
  wire [1:0] _add_map_x_169_sg_left;
  wire [1:0] _add_map_x_169_sg_right;
  wire _add_map_x_169_wall_t_in;
  wire [9:0] _add_map_x_169_moto;
  wire [9:0] _add_map_x_169_up;
  wire [9:0] _add_map_x_169_right;
  wire [9:0] _add_map_x_169_down;
  wire [9:0] _add_map_x_169_left;
  wire [9:0] _add_map_x_169_start;
  wire [9:0] _add_map_x_169_goal;
  wire [9:0] _add_map_x_169_now;
  wire [9:0] _add_map_x_169_data_out;
  wire [9:0] _add_map_x_169_data_out_index;
  wire [9:0] _add_map_x_169_data_near;
  wire _add_map_x_169_wall_t_out;
  wire [9:0] _add_map_x_169_data_org;
  wire [9:0] _add_map_x_169_data_org_near;
  wire [1:0] _add_map_x_169_s_g;
  wire [1:0] _add_map_x_169_s_g_near;
  wire _add_map_x_169_add_exe;
  wire _add_map_x_169_p_reset;
  wire _add_map_x_169_m_clock;
  wire [9:0] _add_map_x_168_moto_org_near;
  wire [9:0] _add_map_x_168_moto_org_near1;
  wire [9:0] _add_map_x_168_moto_org_near2;
  wire [9:0] _add_map_x_168_moto_org_near3;
  wire [9:0] _add_map_x_168_moto_org;
  wire [1:0] _add_map_x_168_sg_up;
  wire [1:0] _add_map_x_168_sg_down;
  wire [1:0] _add_map_x_168_sg_left;
  wire [1:0] _add_map_x_168_sg_right;
  wire _add_map_x_168_wall_t_in;
  wire [9:0] _add_map_x_168_moto;
  wire [9:0] _add_map_x_168_up;
  wire [9:0] _add_map_x_168_right;
  wire [9:0] _add_map_x_168_down;
  wire [9:0] _add_map_x_168_left;
  wire [9:0] _add_map_x_168_start;
  wire [9:0] _add_map_x_168_goal;
  wire [9:0] _add_map_x_168_now;
  wire [9:0] _add_map_x_168_data_out;
  wire [9:0] _add_map_x_168_data_out_index;
  wire [9:0] _add_map_x_168_data_near;
  wire _add_map_x_168_wall_t_out;
  wire [9:0] _add_map_x_168_data_org;
  wire [9:0] _add_map_x_168_data_org_near;
  wire [1:0] _add_map_x_168_s_g;
  wire [1:0] _add_map_x_168_s_g_near;
  wire _add_map_x_168_add_exe;
  wire _add_map_x_168_p_reset;
  wire _add_map_x_168_m_clock;
  wire [9:0] _add_map_x_167_moto_org_near;
  wire [9:0] _add_map_x_167_moto_org_near1;
  wire [9:0] _add_map_x_167_moto_org_near2;
  wire [9:0] _add_map_x_167_moto_org_near3;
  wire [9:0] _add_map_x_167_moto_org;
  wire [1:0] _add_map_x_167_sg_up;
  wire [1:0] _add_map_x_167_sg_down;
  wire [1:0] _add_map_x_167_sg_left;
  wire [1:0] _add_map_x_167_sg_right;
  wire _add_map_x_167_wall_t_in;
  wire [9:0] _add_map_x_167_moto;
  wire [9:0] _add_map_x_167_up;
  wire [9:0] _add_map_x_167_right;
  wire [9:0] _add_map_x_167_down;
  wire [9:0] _add_map_x_167_left;
  wire [9:0] _add_map_x_167_start;
  wire [9:0] _add_map_x_167_goal;
  wire [9:0] _add_map_x_167_now;
  wire [9:0] _add_map_x_167_data_out;
  wire [9:0] _add_map_x_167_data_out_index;
  wire [9:0] _add_map_x_167_data_near;
  wire _add_map_x_167_wall_t_out;
  wire [9:0] _add_map_x_167_data_org;
  wire [9:0] _add_map_x_167_data_org_near;
  wire [1:0] _add_map_x_167_s_g;
  wire [1:0] _add_map_x_167_s_g_near;
  wire _add_map_x_167_add_exe;
  wire _add_map_x_167_p_reset;
  wire _add_map_x_167_m_clock;
  wire [9:0] _add_map_x_166_moto_org_near;
  wire [9:0] _add_map_x_166_moto_org_near1;
  wire [9:0] _add_map_x_166_moto_org_near2;
  wire [9:0] _add_map_x_166_moto_org_near3;
  wire [9:0] _add_map_x_166_moto_org;
  wire [1:0] _add_map_x_166_sg_up;
  wire [1:0] _add_map_x_166_sg_down;
  wire [1:0] _add_map_x_166_sg_left;
  wire [1:0] _add_map_x_166_sg_right;
  wire _add_map_x_166_wall_t_in;
  wire [9:0] _add_map_x_166_moto;
  wire [9:0] _add_map_x_166_up;
  wire [9:0] _add_map_x_166_right;
  wire [9:0] _add_map_x_166_down;
  wire [9:0] _add_map_x_166_left;
  wire [9:0] _add_map_x_166_start;
  wire [9:0] _add_map_x_166_goal;
  wire [9:0] _add_map_x_166_now;
  wire [9:0] _add_map_x_166_data_out;
  wire [9:0] _add_map_x_166_data_out_index;
  wire [9:0] _add_map_x_166_data_near;
  wire _add_map_x_166_wall_t_out;
  wire [9:0] _add_map_x_166_data_org;
  wire [9:0] _add_map_x_166_data_org_near;
  wire [1:0] _add_map_x_166_s_g;
  wire [1:0] _add_map_x_166_s_g_near;
  wire _add_map_x_166_add_exe;
  wire _add_map_x_166_p_reset;
  wire _add_map_x_166_m_clock;
  wire [9:0] _add_map_x_165_moto_org_near;
  wire [9:0] _add_map_x_165_moto_org_near1;
  wire [9:0] _add_map_x_165_moto_org_near2;
  wire [9:0] _add_map_x_165_moto_org_near3;
  wire [9:0] _add_map_x_165_moto_org;
  wire [1:0] _add_map_x_165_sg_up;
  wire [1:0] _add_map_x_165_sg_down;
  wire [1:0] _add_map_x_165_sg_left;
  wire [1:0] _add_map_x_165_sg_right;
  wire _add_map_x_165_wall_t_in;
  wire [9:0] _add_map_x_165_moto;
  wire [9:0] _add_map_x_165_up;
  wire [9:0] _add_map_x_165_right;
  wire [9:0] _add_map_x_165_down;
  wire [9:0] _add_map_x_165_left;
  wire [9:0] _add_map_x_165_start;
  wire [9:0] _add_map_x_165_goal;
  wire [9:0] _add_map_x_165_now;
  wire [9:0] _add_map_x_165_data_out;
  wire [9:0] _add_map_x_165_data_out_index;
  wire [9:0] _add_map_x_165_data_near;
  wire _add_map_x_165_wall_t_out;
  wire [9:0] _add_map_x_165_data_org;
  wire [9:0] _add_map_x_165_data_org_near;
  wire [1:0] _add_map_x_165_s_g;
  wire [1:0] _add_map_x_165_s_g_near;
  wire _add_map_x_165_add_exe;
  wire _add_map_x_165_p_reset;
  wire _add_map_x_165_m_clock;
  wire [9:0] _add_map_x_164_moto_org_near;
  wire [9:0] _add_map_x_164_moto_org_near1;
  wire [9:0] _add_map_x_164_moto_org_near2;
  wire [9:0] _add_map_x_164_moto_org_near3;
  wire [9:0] _add_map_x_164_moto_org;
  wire [1:0] _add_map_x_164_sg_up;
  wire [1:0] _add_map_x_164_sg_down;
  wire [1:0] _add_map_x_164_sg_left;
  wire [1:0] _add_map_x_164_sg_right;
  wire _add_map_x_164_wall_t_in;
  wire [9:0] _add_map_x_164_moto;
  wire [9:0] _add_map_x_164_up;
  wire [9:0] _add_map_x_164_right;
  wire [9:0] _add_map_x_164_down;
  wire [9:0] _add_map_x_164_left;
  wire [9:0] _add_map_x_164_start;
  wire [9:0] _add_map_x_164_goal;
  wire [9:0] _add_map_x_164_now;
  wire [9:0] _add_map_x_164_data_out;
  wire [9:0] _add_map_x_164_data_out_index;
  wire [9:0] _add_map_x_164_data_near;
  wire _add_map_x_164_wall_t_out;
  wire [9:0] _add_map_x_164_data_org;
  wire [9:0] _add_map_x_164_data_org_near;
  wire [1:0] _add_map_x_164_s_g;
  wire [1:0] _add_map_x_164_s_g_near;
  wire _add_map_x_164_add_exe;
  wire _add_map_x_164_p_reset;
  wire _add_map_x_164_m_clock;
  wire [9:0] _add_map_x_163_moto_org_near;
  wire [9:0] _add_map_x_163_moto_org_near1;
  wire [9:0] _add_map_x_163_moto_org_near2;
  wire [9:0] _add_map_x_163_moto_org_near3;
  wire [9:0] _add_map_x_163_moto_org;
  wire [1:0] _add_map_x_163_sg_up;
  wire [1:0] _add_map_x_163_sg_down;
  wire [1:0] _add_map_x_163_sg_left;
  wire [1:0] _add_map_x_163_sg_right;
  wire _add_map_x_163_wall_t_in;
  wire [9:0] _add_map_x_163_moto;
  wire [9:0] _add_map_x_163_up;
  wire [9:0] _add_map_x_163_right;
  wire [9:0] _add_map_x_163_down;
  wire [9:0] _add_map_x_163_left;
  wire [9:0] _add_map_x_163_start;
  wire [9:0] _add_map_x_163_goal;
  wire [9:0] _add_map_x_163_now;
  wire [9:0] _add_map_x_163_data_out;
  wire [9:0] _add_map_x_163_data_out_index;
  wire [9:0] _add_map_x_163_data_near;
  wire _add_map_x_163_wall_t_out;
  wire [9:0] _add_map_x_163_data_org;
  wire [9:0] _add_map_x_163_data_org_near;
  wire [1:0] _add_map_x_163_s_g;
  wire [1:0] _add_map_x_163_s_g_near;
  wire _add_map_x_163_add_exe;
  wire _add_map_x_163_p_reset;
  wire _add_map_x_163_m_clock;
  wire [9:0] _add_map_x_162_moto_org_near;
  wire [9:0] _add_map_x_162_moto_org_near1;
  wire [9:0] _add_map_x_162_moto_org_near2;
  wire [9:0] _add_map_x_162_moto_org_near3;
  wire [9:0] _add_map_x_162_moto_org;
  wire [1:0] _add_map_x_162_sg_up;
  wire [1:0] _add_map_x_162_sg_down;
  wire [1:0] _add_map_x_162_sg_left;
  wire [1:0] _add_map_x_162_sg_right;
  wire _add_map_x_162_wall_t_in;
  wire [9:0] _add_map_x_162_moto;
  wire [9:0] _add_map_x_162_up;
  wire [9:0] _add_map_x_162_right;
  wire [9:0] _add_map_x_162_down;
  wire [9:0] _add_map_x_162_left;
  wire [9:0] _add_map_x_162_start;
  wire [9:0] _add_map_x_162_goal;
  wire [9:0] _add_map_x_162_now;
  wire [9:0] _add_map_x_162_data_out;
  wire [9:0] _add_map_x_162_data_out_index;
  wire [9:0] _add_map_x_162_data_near;
  wire _add_map_x_162_wall_t_out;
  wire [9:0] _add_map_x_162_data_org;
  wire [9:0] _add_map_x_162_data_org_near;
  wire [1:0] _add_map_x_162_s_g;
  wire [1:0] _add_map_x_162_s_g_near;
  wire _add_map_x_162_add_exe;
  wire _add_map_x_162_p_reset;
  wire _add_map_x_162_m_clock;
  wire [9:0] _add_map_x_161_moto_org_near;
  wire [9:0] _add_map_x_161_moto_org_near1;
  wire [9:0] _add_map_x_161_moto_org_near2;
  wire [9:0] _add_map_x_161_moto_org_near3;
  wire [9:0] _add_map_x_161_moto_org;
  wire [1:0] _add_map_x_161_sg_up;
  wire [1:0] _add_map_x_161_sg_down;
  wire [1:0] _add_map_x_161_sg_left;
  wire [1:0] _add_map_x_161_sg_right;
  wire _add_map_x_161_wall_t_in;
  wire [9:0] _add_map_x_161_moto;
  wire [9:0] _add_map_x_161_up;
  wire [9:0] _add_map_x_161_right;
  wire [9:0] _add_map_x_161_down;
  wire [9:0] _add_map_x_161_left;
  wire [9:0] _add_map_x_161_start;
  wire [9:0] _add_map_x_161_goal;
  wire [9:0] _add_map_x_161_now;
  wire [9:0] _add_map_x_161_data_out;
  wire [9:0] _add_map_x_161_data_out_index;
  wire [9:0] _add_map_x_161_data_near;
  wire _add_map_x_161_wall_t_out;
  wire [9:0] _add_map_x_161_data_org;
  wire [9:0] _add_map_x_161_data_org_near;
  wire [1:0] _add_map_x_161_s_g;
  wire [1:0] _add_map_x_161_s_g_near;
  wire _add_map_x_161_add_exe;
  wire _add_map_x_161_p_reset;
  wire _add_map_x_161_m_clock;
  wire [9:0] _add_map_x_160_moto_org_near;
  wire [9:0] _add_map_x_160_moto_org_near1;
  wire [9:0] _add_map_x_160_moto_org_near2;
  wire [9:0] _add_map_x_160_moto_org_near3;
  wire [9:0] _add_map_x_160_moto_org;
  wire [1:0] _add_map_x_160_sg_up;
  wire [1:0] _add_map_x_160_sg_down;
  wire [1:0] _add_map_x_160_sg_left;
  wire [1:0] _add_map_x_160_sg_right;
  wire _add_map_x_160_wall_t_in;
  wire [9:0] _add_map_x_160_moto;
  wire [9:0] _add_map_x_160_up;
  wire [9:0] _add_map_x_160_right;
  wire [9:0] _add_map_x_160_down;
  wire [9:0] _add_map_x_160_left;
  wire [9:0] _add_map_x_160_start;
  wire [9:0] _add_map_x_160_goal;
  wire [9:0] _add_map_x_160_now;
  wire [9:0] _add_map_x_160_data_out;
  wire [9:0] _add_map_x_160_data_out_index;
  wire [9:0] _add_map_x_160_data_near;
  wire _add_map_x_160_wall_t_out;
  wire [9:0] _add_map_x_160_data_org;
  wire [9:0] _add_map_x_160_data_org_near;
  wire [1:0] _add_map_x_160_s_g;
  wire [1:0] _add_map_x_160_s_g_near;
  wire _add_map_x_160_add_exe;
  wire _add_map_x_160_p_reset;
  wire _add_map_x_160_m_clock;
  wire [9:0] _add_map_x_159_moto_org_near;
  wire [9:0] _add_map_x_159_moto_org_near1;
  wire [9:0] _add_map_x_159_moto_org_near2;
  wire [9:0] _add_map_x_159_moto_org_near3;
  wire [9:0] _add_map_x_159_moto_org;
  wire [1:0] _add_map_x_159_sg_up;
  wire [1:0] _add_map_x_159_sg_down;
  wire [1:0] _add_map_x_159_sg_left;
  wire [1:0] _add_map_x_159_sg_right;
  wire _add_map_x_159_wall_t_in;
  wire [9:0] _add_map_x_159_moto;
  wire [9:0] _add_map_x_159_up;
  wire [9:0] _add_map_x_159_right;
  wire [9:0] _add_map_x_159_down;
  wire [9:0] _add_map_x_159_left;
  wire [9:0] _add_map_x_159_start;
  wire [9:0] _add_map_x_159_goal;
  wire [9:0] _add_map_x_159_now;
  wire [9:0] _add_map_x_159_data_out;
  wire [9:0] _add_map_x_159_data_out_index;
  wire [9:0] _add_map_x_159_data_near;
  wire _add_map_x_159_wall_t_out;
  wire [9:0] _add_map_x_159_data_org;
  wire [9:0] _add_map_x_159_data_org_near;
  wire [1:0] _add_map_x_159_s_g;
  wire [1:0] _add_map_x_159_s_g_near;
  wire _add_map_x_159_add_exe;
  wire _add_map_x_159_p_reset;
  wire _add_map_x_159_m_clock;
  wire [9:0] _add_map_x_158_moto_org_near;
  wire [9:0] _add_map_x_158_moto_org_near1;
  wire [9:0] _add_map_x_158_moto_org_near2;
  wire [9:0] _add_map_x_158_moto_org_near3;
  wire [9:0] _add_map_x_158_moto_org;
  wire [1:0] _add_map_x_158_sg_up;
  wire [1:0] _add_map_x_158_sg_down;
  wire [1:0] _add_map_x_158_sg_left;
  wire [1:0] _add_map_x_158_sg_right;
  wire _add_map_x_158_wall_t_in;
  wire [9:0] _add_map_x_158_moto;
  wire [9:0] _add_map_x_158_up;
  wire [9:0] _add_map_x_158_right;
  wire [9:0] _add_map_x_158_down;
  wire [9:0] _add_map_x_158_left;
  wire [9:0] _add_map_x_158_start;
  wire [9:0] _add_map_x_158_goal;
  wire [9:0] _add_map_x_158_now;
  wire [9:0] _add_map_x_158_data_out;
  wire [9:0] _add_map_x_158_data_out_index;
  wire [9:0] _add_map_x_158_data_near;
  wire _add_map_x_158_wall_t_out;
  wire [9:0] _add_map_x_158_data_org;
  wire [9:0] _add_map_x_158_data_org_near;
  wire [1:0] _add_map_x_158_s_g;
  wire [1:0] _add_map_x_158_s_g_near;
  wire _add_map_x_158_add_exe;
  wire _add_map_x_158_p_reset;
  wire _add_map_x_158_m_clock;
  wire [9:0] _add_map_x_157_moto_org_near;
  wire [9:0] _add_map_x_157_moto_org_near1;
  wire [9:0] _add_map_x_157_moto_org_near2;
  wire [9:0] _add_map_x_157_moto_org_near3;
  wire [9:0] _add_map_x_157_moto_org;
  wire [1:0] _add_map_x_157_sg_up;
  wire [1:0] _add_map_x_157_sg_down;
  wire [1:0] _add_map_x_157_sg_left;
  wire [1:0] _add_map_x_157_sg_right;
  wire _add_map_x_157_wall_t_in;
  wire [9:0] _add_map_x_157_moto;
  wire [9:0] _add_map_x_157_up;
  wire [9:0] _add_map_x_157_right;
  wire [9:0] _add_map_x_157_down;
  wire [9:0] _add_map_x_157_left;
  wire [9:0] _add_map_x_157_start;
  wire [9:0] _add_map_x_157_goal;
  wire [9:0] _add_map_x_157_now;
  wire [9:0] _add_map_x_157_data_out;
  wire [9:0] _add_map_x_157_data_out_index;
  wire [9:0] _add_map_x_157_data_near;
  wire _add_map_x_157_wall_t_out;
  wire [9:0] _add_map_x_157_data_org;
  wire [9:0] _add_map_x_157_data_org_near;
  wire [1:0] _add_map_x_157_s_g;
  wire [1:0] _add_map_x_157_s_g_near;
  wire _add_map_x_157_add_exe;
  wire _add_map_x_157_p_reset;
  wire _add_map_x_157_m_clock;
  wire [9:0] _add_map_x_156_moto_org_near;
  wire [9:0] _add_map_x_156_moto_org_near1;
  wire [9:0] _add_map_x_156_moto_org_near2;
  wire [9:0] _add_map_x_156_moto_org_near3;
  wire [9:0] _add_map_x_156_moto_org;
  wire [1:0] _add_map_x_156_sg_up;
  wire [1:0] _add_map_x_156_sg_down;
  wire [1:0] _add_map_x_156_sg_left;
  wire [1:0] _add_map_x_156_sg_right;
  wire _add_map_x_156_wall_t_in;
  wire [9:0] _add_map_x_156_moto;
  wire [9:0] _add_map_x_156_up;
  wire [9:0] _add_map_x_156_right;
  wire [9:0] _add_map_x_156_down;
  wire [9:0] _add_map_x_156_left;
  wire [9:0] _add_map_x_156_start;
  wire [9:0] _add_map_x_156_goal;
  wire [9:0] _add_map_x_156_now;
  wire [9:0] _add_map_x_156_data_out;
  wire [9:0] _add_map_x_156_data_out_index;
  wire [9:0] _add_map_x_156_data_near;
  wire _add_map_x_156_wall_t_out;
  wire [9:0] _add_map_x_156_data_org;
  wire [9:0] _add_map_x_156_data_org_near;
  wire [1:0] _add_map_x_156_s_g;
  wire [1:0] _add_map_x_156_s_g_near;
  wire _add_map_x_156_add_exe;
  wire _add_map_x_156_p_reset;
  wire _add_map_x_156_m_clock;
  wire [9:0] _add_map_x_155_moto_org_near;
  wire [9:0] _add_map_x_155_moto_org_near1;
  wire [9:0] _add_map_x_155_moto_org_near2;
  wire [9:0] _add_map_x_155_moto_org_near3;
  wire [9:0] _add_map_x_155_moto_org;
  wire [1:0] _add_map_x_155_sg_up;
  wire [1:0] _add_map_x_155_sg_down;
  wire [1:0] _add_map_x_155_sg_left;
  wire [1:0] _add_map_x_155_sg_right;
  wire _add_map_x_155_wall_t_in;
  wire [9:0] _add_map_x_155_moto;
  wire [9:0] _add_map_x_155_up;
  wire [9:0] _add_map_x_155_right;
  wire [9:0] _add_map_x_155_down;
  wire [9:0] _add_map_x_155_left;
  wire [9:0] _add_map_x_155_start;
  wire [9:0] _add_map_x_155_goal;
  wire [9:0] _add_map_x_155_now;
  wire [9:0] _add_map_x_155_data_out;
  wire [9:0] _add_map_x_155_data_out_index;
  wire [9:0] _add_map_x_155_data_near;
  wire _add_map_x_155_wall_t_out;
  wire [9:0] _add_map_x_155_data_org;
  wire [9:0] _add_map_x_155_data_org_near;
  wire [1:0] _add_map_x_155_s_g;
  wire [1:0] _add_map_x_155_s_g_near;
  wire _add_map_x_155_add_exe;
  wire _add_map_x_155_p_reset;
  wire _add_map_x_155_m_clock;
  wire [9:0] _add_map_x_154_moto_org_near;
  wire [9:0] _add_map_x_154_moto_org_near1;
  wire [9:0] _add_map_x_154_moto_org_near2;
  wire [9:0] _add_map_x_154_moto_org_near3;
  wire [9:0] _add_map_x_154_moto_org;
  wire [1:0] _add_map_x_154_sg_up;
  wire [1:0] _add_map_x_154_sg_down;
  wire [1:0] _add_map_x_154_sg_left;
  wire [1:0] _add_map_x_154_sg_right;
  wire _add_map_x_154_wall_t_in;
  wire [9:0] _add_map_x_154_moto;
  wire [9:0] _add_map_x_154_up;
  wire [9:0] _add_map_x_154_right;
  wire [9:0] _add_map_x_154_down;
  wire [9:0] _add_map_x_154_left;
  wire [9:0] _add_map_x_154_start;
  wire [9:0] _add_map_x_154_goal;
  wire [9:0] _add_map_x_154_now;
  wire [9:0] _add_map_x_154_data_out;
  wire [9:0] _add_map_x_154_data_out_index;
  wire [9:0] _add_map_x_154_data_near;
  wire _add_map_x_154_wall_t_out;
  wire [9:0] _add_map_x_154_data_org;
  wire [9:0] _add_map_x_154_data_org_near;
  wire [1:0] _add_map_x_154_s_g;
  wire [1:0] _add_map_x_154_s_g_near;
  wire _add_map_x_154_add_exe;
  wire _add_map_x_154_p_reset;
  wire _add_map_x_154_m_clock;
  wire [9:0] _add_map_x_153_moto_org_near;
  wire [9:0] _add_map_x_153_moto_org_near1;
  wire [9:0] _add_map_x_153_moto_org_near2;
  wire [9:0] _add_map_x_153_moto_org_near3;
  wire [9:0] _add_map_x_153_moto_org;
  wire [1:0] _add_map_x_153_sg_up;
  wire [1:0] _add_map_x_153_sg_down;
  wire [1:0] _add_map_x_153_sg_left;
  wire [1:0] _add_map_x_153_sg_right;
  wire _add_map_x_153_wall_t_in;
  wire [9:0] _add_map_x_153_moto;
  wire [9:0] _add_map_x_153_up;
  wire [9:0] _add_map_x_153_right;
  wire [9:0] _add_map_x_153_down;
  wire [9:0] _add_map_x_153_left;
  wire [9:0] _add_map_x_153_start;
  wire [9:0] _add_map_x_153_goal;
  wire [9:0] _add_map_x_153_now;
  wire [9:0] _add_map_x_153_data_out;
  wire [9:0] _add_map_x_153_data_out_index;
  wire [9:0] _add_map_x_153_data_near;
  wire _add_map_x_153_wall_t_out;
  wire [9:0] _add_map_x_153_data_org;
  wire [9:0] _add_map_x_153_data_org_near;
  wire [1:0] _add_map_x_153_s_g;
  wire [1:0] _add_map_x_153_s_g_near;
  wire _add_map_x_153_add_exe;
  wire _add_map_x_153_p_reset;
  wire _add_map_x_153_m_clock;
  wire [9:0] _add_map_x_152_moto_org_near;
  wire [9:0] _add_map_x_152_moto_org_near1;
  wire [9:0] _add_map_x_152_moto_org_near2;
  wire [9:0] _add_map_x_152_moto_org_near3;
  wire [9:0] _add_map_x_152_moto_org;
  wire [1:0] _add_map_x_152_sg_up;
  wire [1:0] _add_map_x_152_sg_down;
  wire [1:0] _add_map_x_152_sg_left;
  wire [1:0] _add_map_x_152_sg_right;
  wire _add_map_x_152_wall_t_in;
  wire [9:0] _add_map_x_152_moto;
  wire [9:0] _add_map_x_152_up;
  wire [9:0] _add_map_x_152_right;
  wire [9:0] _add_map_x_152_down;
  wire [9:0] _add_map_x_152_left;
  wire [9:0] _add_map_x_152_start;
  wire [9:0] _add_map_x_152_goal;
  wire [9:0] _add_map_x_152_now;
  wire [9:0] _add_map_x_152_data_out;
  wire [9:0] _add_map_x_152_data_out_index;
  wire [9:0] _add_map_x_152_data_near;
  wire _add_map_x_152_wall_t_out;
  wire [9:0] _add_map_x_152_data_org;
  wire [9:0] _add_map_x_152_data_org_near;
  wire [1:0] _add_map_x_152_s_g;
  wire [1:0] _add_map_x_152_s_g_near;
  wire _add_map_x_152_add_exe;
  wire _add_map_x_152_p_reset;
  wire _add_map_x_152_m_clock;
  wire [9:0] _add_map_x_151_moto_org_near;
  wire [9:0] _add_map_x_151_moto_org_near1;
  wire [9:0] _add_map_x_151_moto_org_near2;
  wire [9:0] _add_map_x_151_moto_org_near3;
  wire [9:0] _add_map_x_151_moto_org;
  wire [1:0] _add_map_x_151_sg_up;
  wire [1:0] _add_map_x_151_sg_down;
  wire [1:0] _add_map_x_151_sg_left;
  wire [1:0] _add_map_x_151_sg_right;
  wire _add_map_x_151_wall_t_in;
  wire [9:0] _add_map_x_151_moto;
  wire [9:0] _add_map_x_151_up;
  wire [9:0] _add_map_x_151_right;
  wire [9:0] _add_map_x_151_down;
  wire [9:0] _add_map_x_151_left;
  wire [9:0] _add_map_x_151_start;
  wire [9:0] _add_map_x_151_goal;
  wire [9:0] _add_map_x_151_now;
  wire [9:0] _add_map_x_151_data_out;
  wire [9:0] _add_map_x_151_data_out_index;
  wire [9:0] _add_map_x_151_data_near;
  wire _add_map_x_151_wall_t_out;
  wire [9:0] _add_map_x_151_data_org;
  wire [9:0] _add_map_x_151_data_org_near;
  wire [1:0] _add_map_x_151_s_g;
  wire [1:0] _add_map_x_151_s_g_near;
  wire _add_map_x_151_add_exe;
  wire _add_map_x_151_p_reset;
  wire _add_map_x_151_m_clock;
  wire [9:0] _add_map_x_150_moto_org_near;
  wire [9:0] _add_map_x_150_moto_org_near1;
  wire [9:0] _add_map_x_150_moto_org_near2;
  wire [9:0] _add_map_x_150_moto_org_near3;
  wire [9:0] _add_map_x_150_moto_org;
  wire [1:0] _add_map_x_150_sg_up;
  wire [1:0] _add_map_x_150_sg_down;
  wire [1:0] _add_map_x_150_sg_left;
  wire [1:0] _add_map_x_150_sg_right;
  wire _add_map_x_150_wall_t_in;
  wire [9:0] _add_map_x_150_moto;
  wire [9:0] _add_map_x_150_up;
  wire [9:0] _add_map_x_150_right;
  wire [9:0] _add_map_x_150_down;
  wire [9:0] _add_map_x_150_left;
  wire [9:0] _add_map_x_150_start;
  wire [9:0] _add_map_x_150_goal;
  wire [9:0] _add_map_x_150_now;
  wire [9:0] _add_map_x_150_data_out;
  wire [9:0] _add_map_x_150_data_out_index;
  wire [9:0] _add_map_x_150_data_near;
  wire _add_map_x_150_wall_t_out;
  wire [9:0] _add_map_x_150_data_org;
  wire [9:0] _add_map_x_150_data_org_near;
  wire [1:0] _add_map_x_150_s_g;
  wire [1:0] _add_map_x_150_s_g_near;
  wire _add_map_x_150_add_exe;
  wire _add_map_x_150_p_reset;
  wire _add_map_x_150_m_clock;
  wire [9:0] _add_map_x_149_moto_org_near;
  wire [9:0] _add_map_x_149_moto_org_near1;
  wire [9:0] _add_map_x_149_moto_org_near2;
  wire [9:0] _add_map_x_149_moto_org_near3;
  wire [9:0] _add_map_x_149_moto_org;
  wire [1:0] _add_map_x_149_sg_up;
  wire [1:0] _add_map_x_149_sg_down;
  wire [1:0] _add_map_x_149_sg_left;
  wire [1:0] _add_map_x_149_sg_right;
  wire _add_map_x_149_wall_t_in;
  wire [9:0] _add_map_x_149_moto;
  wire [9:0] _add_map_x_149_up;
  wire [9:0] _add_map_x_149_right;
  wire [9:0] _add_map_x_149_down;
  wire [9:0] _add_map_x_149_left;
  wire [9:0] _add_map_x_149_start;
  wire [9:0] _add_map_x_149_goal;
  wire [9:0] _add_map_x_149_now;
  wire [9:0] _add_map_x_149_data_out;
  wire [9:0] _add_map_x_149_data_out_index;
  wire [9:0] _add_map_x_149_data_near;
  wire _add_map_x_149_wall_t_out;
  wire [9:0] _add_map_x_149_data_org;
  wire [9:0] _add_map_x_149_data_org_near;
  wire [1:0] _add_map_x_149_s_g;
  wire [1:0] _add_map_x_149_s_g_near;
  wire _add_map_x_149_add_exe;
  wire _add_map_x_149_p_reset;
  wire _add_map_x_149_m_clock;
  wire [9:0] _add_map_x_148_moto_org_near;
  wire [9:0] _add_map_x_148_moto_org_near1;
  wire [9:0] _add_map_x_148_moto_org_near2;
  wire [9:0] _add_map_x_148_moto_org_near3;
  wire [9:0] _add_map_x_148_moto_org;
  wire [1:0] _add_map_x_148_sg_up;
  wire [1:0] _add_map_x_148_sg_down;
  wire [1:0] _add_map_x_148_sg_left;
  wire [1:0] _add_map_x_148_sg_right;
  wire _add_map_x_148_wall_t_in;
  wire [9:0] _add_map_x_148_moto;
  wire [9:0] _add_map_x_148_up;
  wire [9:0] _add_map_x_148_right;
  wire [9:0] _add_map_x_148_down;
  wire [9:0] _add_map_x_148_left;
  wire [9:0] _add_map_x_148_start;
  wire [9:0] _add_map_x_148_goal;
  wire [9:0] _add_map_x_148_now;
  wire [9:0] _add_map_x_148_data_out;
  wire [9:0] _add_map_x_148_data_out_index;
  wire [9:0] _add_map_x_148_data_near;
  wire _add_map_x_148_wall_t_out;
  wire [9:0] _add_map_x_148_data_org;
  wire [9:0] _add_map_x_148_data_org_near;
  wire [1:0] _add_map_x_148_s_g;
  wire [1:0] _add_map_x_148_s_g_near;
  wire _add_map_x_148_add_exe;
  wire _add_map_x_148_p_reset;
  wire _add_map_x_148_m_clock;
  wire [9:0] _add_map_x_147_moto_org_near;
  wire [9:0] _add_map_x_147_moto_org_near1;
  wire [9:0] _add_map_x_147_moto_org_near2;
  wire [9:0] _add_map_x_147_moto_org_near3;
  wire [9:0] _add_map_x_147_moto_org;
  wire [1:0] _add_map_x_147_sg_up;
  wire [1:0] _add_map_x_147_sg_down;
  wire [1:0] _add_map_x_147_sg_left;
  wire [1:0] _add_map_x_147_sg_right;
  wire _add_map_x_147_wall_t_in;
  wire [9:0] _add_map_x_147_moto;
  wire [9:0] _add_map_x_147_up;
  wire [9:0] _add_map_x_147_right;
  wire [9:0] _add_map_x_147_down;
  wire [9:0] _add_map_x_147_left;
  wire [9:0] _add_map_x_147_start;
  wire [9:0] _add_map_x_147_goal;
  wire [9:0] _add_map_x_147_now;
  wire [9:0] _add_map_x_147_data_out;
  wire [9:0] _add_map_x_147_data_out_index;
  wire [9:0] _add_map_x_147_data_near;
  wire _add_map_x_147_wall_t_out;
  wire [9:0] _add_map_x_147_data_org;
  wire [9:0] _add_map_x_147_data_org_near;
  wire [1:0] _add_map_x_147_s_g;
  wire [1:0] _add_map_x_147_s_g_near;
  wire _add_map_x_147_add_exe;
  wire _add_map_x_147_p_reset;
  wire _add_map_x_147_m_clock;
  wire [9:0] _add_map_x_146_moto_org_near;
  wire [9:0] _add_map_x_146_moto_org_near1;
  wire [9:0] _add_map_x_146_moto_org_near2;
  wire [9:0] _add_map_x_146_moto_org_near3;
  wire [9:0] _add_map_x_146_moto_org;
  wire [1:0] _add_map_x_146_sg_up;
  wire [1:0] _add_map_x_146_sg_down;
  wire [1:0] _add_map_x_146_sg_left;
  wire [1:0] _add_map_x_146_sg_right;
  wire _add_map_x_146_wall_t_in;
  wire [9:0] _add_map_x_146_moto;
  wire [9:0] _add_map_x_146_up;
  wire [9:0] _add_map_x_146_right;
  wire [9:0] _add_map_x_146_down;
  wire [9:0] _add_map_x_146_left;
  wire [9:0] _add_map_x_146_start;
  wire [9:0] _add_map_x_146_goal;
  wire [9:0] _add_map_x_146_now;
  wire [9:0] _add_map_x_146_data_out;
  wire [9:0] _add_map_x_146_data_out_index;
  wire [9:0] _add_map_x_146_data_near;
  wire _add_map_x_146_wall_t_out;
  wire [9:0] _add_map_x_146_data_org;
  wire [9:0] _add_map_x_146_data_org_near;
  wire [1:0] _add_map_x_146_s_g;
  wire [1:0] _add_map_x_146_s_g_near;
  wire _add_map_x_146_add_exe;
  wire _add_map_x_146_p_reset;
  wire _add_map_x_146_m_clock;
  wire [9:0] _add_map_x_145_moto_org_near;
  wire [9:0] _add_map_x_145_moto_org_near1;
  wire [9:0] _add_map_x_145_moto_org_near2;
  wire [9:0] _add_map_x_145_moto_org_near3;
  wire [9:0] _add_map_x_145_moto_org;
  wire [1:0] _add_map_x_145_sg_up;
  wire [1:0] _add_map_x_145_sg_down;
  wire [1:0] _add_map_x_145_sg_left;
  wire [1:0] _add_map_x_145_sg_right;
  wire _add_map_x_145_wall_t_in;
  wire [9:0] _add_map_x_145_moto;
  wire [9:0] _add_map_x_145_up;
  wire [9:0] _add_map_x_145_right;
  wire [9:0] _add_map_x_145_down;
  wire [9:0] _add_map_x_145_left;
  wire [9:0] _add_map_x_145_start;
  wire [9:0] _add_map_x_145_goal;
  wire [9:0] _add_map_x_145_now;
  wire [9:0] _add_map_x_145_data_out;
  wire [9:0] _add_map_x_145_data_out_index;
  wire [9:0] _add_map_x_145_data_near;
  wire _add_map_x_145_wall_t_out;
  wire [9:0] _add_map_x_145_data_org;
  wire [9:0] _add_map_x_145_data_org_near;
  wire [1:0] _add_map_x_145_s_g;
  wire [1:0] _add_map_x_145_s_g_near;
  wire _add_map_x_145_add_exe;
  wire _add_map_x_145_p_reset;
  wire _add_map_x_145_m_clock;
  wire [9:0] _add_map_x_144_moto_org_near;
  wire [9:0] _add_map_x_144_moto_org_near1;
  wire [9:0] _add_map_x_144_moto_org_near2;
  wire [9:0] _add_map_x_144_moto_org_near3;
  wire [9:0] _add_map_x_144_moto_org;
  wire [1:0] _add_map_x_144_sg_up;
  wire [1:0] _add_map_x_144_sg_down;
  wire [1:0] _add_map_x_144_sg_left;
  wire [1:0] _add_map_x_144_sg_right;
  wire _add_map_x_144_wall_t_in;
  wire [9:0] _add_map_x_144_moto;
  wire [9:0] _add_map_x_144_up;
  wire [9:0] _add_map_x_144_right;
  wire [9:0] _add_map_x_144_down;
  wire [9:0] _add_map_x_144_left;
  wire [9:0] _add_map_x_144_start;
  wire [9:0] _add_map_x_144_goal;
  wire [9:0] _add_map_x_144_now;
  wire [9:0] _add_map_x_144_data_out;
  wire [9:0] _add_map_x_144_data_out_index;
  wire [9:0] _add_map_x_144_data_near;
  wire _add_map_x_144_wall_t_out;
  wire [9:0] _add_map_x_144_data_org;
  wire [9:0] _add_map_x_144_data_org_near;
  wire [1:0] _add_map_x_144_s_g;
  wire [1:0] _add_map_x_144_s_g_near;
  wire _add_map_x_144_add_exe;
  wire _add_map_x_144_p_reset;
  wire _add_map_x_144_m_clock;
  wire [9:0] _add_map_x_143_moto_org_near;
  wire [9:0] _add_map_x_143_moto_org_near1;
  wire [9:0] _add_map_x_143_moto_org_near2;
  wire [9:0] _add_map_x_143_moto_org_near3;
  wire [9:0] _add_map_x_143_moto_org;
  wire [1:0] _add_map_x_143_sg_up;
  wire [1:0] _add_map_x_143_sg_down;
  wire [1:0] _add_map_x_143_sg_left;
  wire [1:0] _add_map_x_143_sg_right;
  wire _add_map_x_143_wall_t_in;
  wire [9:0] _add_map_x_143_moto;
  wire [9:0] _add_map_x_143_up;
  wire [9:0] _add_map_x_143_right;
  wire [9:0] _add_map_x_143_down;
  wire [9:0] _add_map_x_143_left;
  wire [9:0] _add_map_x_143_start;
  wire [9:0] _add_map_x_143_goal;
  wire [9:0] _add_map_x_143_now;
  wire [9:0] _add_map_x_143_data_out;
  wire [9:0] _add_map_x_143_data_out_index;
  wire [9:0] _add_map_x_143_data_near;
  wire _add_map_x_143_wall_t_out;
  wire [9:0] _add_map_x_143_data_org;
  wire [9:0] _add_map_x_143_data_org_near;
  wire [1:0] _add_map_x_143_s_g;
  wire [1:0] _add_map_x_143_s_g_near;
  wire _add_map_x_143_add_exe;
  wire _add_map_x_143_p_reset;
  wire _add_map_x_143_m_clock;
  wire [9:0] _add_map_x_142_moto_org_near;
  wire [9:0] _add_map_x_142_moto_org_near1;
  wire [9:0] _add_map_x_142_moto_org_near2;
  wire [9:0] _add_map_x_142_moto_org_near3;
  wire [9:0] _add_map_x_142_moto_org;
  wire [1:0] _add_map_x_142_sg_up;
  wire [1:0] _add_map_x_142_sg_down;
  wire [1:0] _add_map_x_142_sg_left;
  wire [1:0] _add_map_x_142_sg_right;
  wire _add_map_x_142_wall_t_in;
  wire [9:0] _add_map_x_142_moto;
  wire [9:0] _add_map_x_142_up;
  wire [9:0] _add_map_x_142_right;
  wire [9:0] _add_map_x_142_down;
  wire [9:0] _add_map_x_142_left;
  wire [9:0] _add_map_x_142_start;
  wire [9:0] _add_map_x_142_goal;
  wire [9:0] _add_map_x_142_now;
  wire [9:0] _add_map_x_142_data_out;
  wire [9:0] _add_map_x_142_data_out_index;
  wire [9:0] _add_map_x_142_data_near;
  wire _add_map_x_142_wall_t_out;
  wire [9:0] _add_map_x_142_data_org;
  wire [9:0] _add_map_x_142_data_org_near;
  wire [1:0] _add_map_x_142_s_g;
  wire [1:0] _add_map_x_142_s_g_near;
  wire _add_map_x_142_add_exe;
  wire _add_map_x_142_p_reset;
  wire _add_map_x_142_m_clock;
  wire [9:0] _add_map_x_141_moto_org_near;
  wire [9:0] _add_map_x_141_moto_org_near1;
  wire [9:0] _add_map_x_141_moto_org_near2;
  wire [9:0] _add_map_x_141_moto_org_near3;
  wire [9:0] _add_map_x_141_moto_org;
  wire [1:0] _add_map_x_141_sg_up;
  wire [1:0] _add_map_x_141_sg_down;
  wire [1:0] _add_map_x_141_sg_left;
  wire [1:0] _add_map_x_141_sg_right;
  wire _add_map_x_141_wall_t_in;
  wire [9:0] _add_map_x_141_moto;
  wire [9:0] _add_map_x_141_up;
  wire [9:0] _add_map_x_141_right;
  wire [9:0] _add_map_x_141_down;
  wire [9:0] _add_map_x_141_left;
  wire [9:0] _add_map_x_141_start;
  wire [9:0] _add_map_x_141_goal;
  wire [9:0] _add_map_x_141_now;
  wire [9:0] _add_map_x_141_data_out;
  wire [9:0] _add_map_x_141_data_out_index;
  wire [9:0] _add_map_x_141_data_near;
  wire _add_map_x_141_wall_t_out;
  wire [9:0] _add_map_x_141_data_org;
  wire [9:0] _add_map_x_141_data_org_near;
  wire [1:0] _add_map_x_141_s_g;
  wire [1:0] _add_map_x_141_s_g_near;
  wire _add_map_x_141_add_exe;
  wire _add_map_x_141_p_reset;
  wire _add_map_x_141_m_clock;
  wire [9:0] _add_map_x_140_moto_org_near;
  wire [9:0] _add_map_x_140_moto_org_near1;
  wire [9:0] _add_map_x_140_moto_org_near2;
  wire [9:0] _add_map_x_140_moto_org_near3;
  wire [9:0] _add_map_x_140_moto_org;
  wire [1:0] _add_map_x_140_sg_up;
  wire [1:0] _add_map_x_140_sg_down;
  wire [1:0] _add_map_x_140_sg_left;
  wire [1:0] _add_map_x_140_sg_right;
  wire _add_map_x_140_wall_t_in;
  wire [9:0] _add_map_x_140_moto;
  wire [9:0] _add_map_x_140_up;
  wire [9:0] _add_map_x_140_right;
  wire [9:0] _add_map_x_140_down;
  wire [9:0] _add_map_x_140_left;
  wire [9:0] _add_map_x_140_start;
  wire [9:0] _add_map_x_140_goal;
  wire [9:0] _add_map_x_140_now;
  wire [9:0] _add_map_x_140_data_out;
  wire [9:0] _add_map_x_140_data_out_index;
  wire [9:0] _add_map_x_140_data_near;
  wire _add_map_x_140_wall_t_out;
  wire [9:0] _add_map_x_140_data_org;
  wire [9:0] _add_map_x_140_data_org_near;
  wire [1:0] _add_map_x_140_s_g;
  wire [1:0] _add_map_x_140_s_g_near;
  wire _add_map_x_140_add_exe;
  wire _add_map_x_140_p_reset;
  wire _add_map_x_140_m_clock;
  wire [9:0] _add_map_x_139_moto_org_near;
  wire [9:0] _add_map_x_139_moto_org_near1;
  wire [9:0] _add_map_x_139_moto_org_near2;
  wire [9:0] _add_map_x_139_moto_org_near3;
  wire [9:0] _add_map_x_139_moto_org;
  wire [1:0] _add_map_x_139_sg_up;
  wire [1:0] _add_map_x_139_sg_down;
  wire [1:0] _add_map_x_139_sg_left;
  wire [1:0] _add_map_x_139_sg_right;
  wire _add_map_x_139_wall_t_in;
  wire [9:0] _add_map_x_139_moto;
  wire [9:0] _add_map_x_139_up;
  wire [9:0] _add_map_x_139_right;
  wire [9:0] _add_map_x_139_down;
  wire [9:0] _add_map_x_139_left;
  wire [9:0] _add_map_x_139_start;
  wire [9:0] _add_map_x_139_goal;
  wire [9:0] _add_map_x_139_now;
  wire [9:0] _add_map_x_139_data_out;
  wire [9:0] _add_map_x_139_data_out_index;
  wire [9:0] _add_map_x_139_data_near;
  wire _add_map_x_139_wall_t_out;
  wire [9:0] _add_map_x_139_data_org;
  wire [9:0] _add_map_x_139_data_org_near;
  wire [1:0] _add_map_x_139_s_g;
  wire [1:0] _add_map_x_139_s_g_near;
  wire _add_map_x_139_add_exe;
  wire _add_map_x_139_p_reset;
  wire _add_map_x_139_m_clock;
  wire [9:0] _add_map_x_138_moto_org_near;
  wire [9:0] _add_map_x_138_moto_org_near1;
  wire [9:0] _add_map_x_138_moto_org_near2;
  wire [9:0] _add_map_x_138_moto_org_near3;
  wire [9:0] _add_map_x_138_moto_org;
  wire [1:0] _add_map_x_138_sg_up;
  wire [1:0] _add_map_x_138_sg_down;
  wire [1:0] _add_map_x_138_sg_left;
  wire [1:0] _add_map_x_138_sg_right;
  wire _add_map_x_138_wall_t_in;
  wire [9:0] _add_map_x_138_moto;
  wire [9:0] _add_map_x_138_up;
  wire [9:0] _add_map_x_138_right;
  wire [9:0] _add_map_x_138_down;
  wire [9:0] _add_map_x_138_left;
  wire [9:0] _add_map_x_138_start;
  wire [9:0] _add_map_x_138_goal;
  wire [9:0] _add_map_x_138_now;
  wire [9:0] _add_map_x_138_data_out;
  wire [9:0] _add_map_x_138_data_out_index;
  wire [9:0] _add_map_x_138_data_near;
  wire _add_map_x_138_wall_t_out;
  wire [9:0] _add_map_x_138_data_org;
  wire [9:0] _add_map_x_138_data_org_near;
  wire [1:0] _add_map_x_138_s_g;
  wire [1:0] _add_map_x_138_s_g_near;
  wire _add_map_x_138_add_exe;
  wire _add_map_x_138_p_reset;
  wire _add_map_x_138_m_clock;
  wire [9:0] _add_map_x_137_moto_org_near;
  wire [9:0] _add_map_x_137_moto_org_near1;
  wire [9:0] _add_map_x_137_moto_org_near2;
  wire [9:0] _add_map_x_137_moto_org_near3;
  wire [9:0] _add_map_x_137_moto_org;
  wire [1:0] _add_map_x_137_sg_up;
  wire [1:0] _add_map_x_137_sg_down;
  wire [1:0] _add_map_x_137_sg_left;
  wire [1:0] _add_map_x_137_sg_right;
  wire _add_map_x_137_wall_t_in;
  wire [9:0] _add_map_x_137_moto;
  wire [9:0] _add_map_x_137_up;
  wire [9:0] _add_map_x_137_right;
  wire [9:0] _add_map_x_137_down;
  wire [9:0] _add_map_x_137_left;
  wire [9:0] _add_map_x_137_start;
  wire [9:0] _add_map_x_137_goal;
  wire [9:0] _add_map_x_137_now;
  wire [9:0] _add_map_x_137_data_out;
  wire [9:0] _add_map_x_137_data_out_index;
  wire [9:0] _add_map_x_137_data_near;
  wire _add_map_x_137_wall_t_out;
  wire [9:0] _add_map_x_137_data_org;
  wire [9:0] _add_map_x_137_data_org_near;
  wire [1:0] _add_map_x_137_s_g;
  wire [1:0] _add_map_x_137_s_g_near;
  wire _add_map_x_137_add_exe;
  wire _add_map_x_137_p_reset;
  wire _add_map_x_137_m_clock;
  wire [9:0] _add_map_x_136_moto_org_near;
  wire [9:0] _add_map_x_136_moto_org_near1;
  wire [9:0] _add_map_x_136_moto_org_near2;
  wire [9:0] _add_map_x_136_moto_org_near3;
  wire [9:0] _add_map_x_136_moto_org;
  wire [1:0] _add_map_x_136_sg_up;
  wire [1:0] _add_map_x_136_sg_down;
  wire [1:0] _add_map_x_136_sg_left;
  wire [1:0] _add_map_x_136_sg_right;
  wire _add_map_x_136_wall_t_in;
  wire [9:0] _add_map_x_136_moto;
  wire [9:0] _add_map_x_136_up;
  wire [9:0] _add_map_x_136_right;
  wire [9:0] _add_map_x_136_down;
  wire [9:0] _add_map_x_136_left;
  wire [9:0] _add_map_x_136_start;
  wire [9:0] _add_map_x_136_goal;
  wire [9:0] _add_map_x_136_now;
  wire [9:0] _add_map_x_136_data_out;
  wire [9:0] _add_map_x_136_data_out_index;
  wire [9:0] _add_map_x_136_data_near;
  wire _add_map_x_136_wall_t_out;
  wire [9:0] _add_map_x_136_data_org;
  wire [9:0] _add_map_x_136_data_org_near;
  wire [1:0] _add_map_x_136_s_g;
  wire [1:0] _add_map_x_136_s_g_near;
  wire _add_map_x_136_add_exe;
  wire _add_map_x_136_p_reset;
  wire _add_map_x_136_m_clock;
  wire [9:0] _add_map_x_135_moto_org_near;
  wire [9:0] _add_map_x_135_moto_org_near1;
  wire [9:0] _add_map_x_135_moto_org_near2;
  wire [9:0] _add_map_x_135_moto_org_near3;
  wire [9:0] _add_map_x_135_moto_org;
  wire [1:0] _add_map_x_135_sg_up;
  wire [1:0] _add_map_x_135_sg_down;
  wire [1:0] _add_map_x_135_sg_left;
  wire [1:0] _add_map_x_135_sg_right;
  wire _add_map_x_135_wall_t_in;
  wire [9:0] _add_map_x_135_moto;
  wire [9:0] _add_map_x_135_up;
  wire [9:0] _add_map_x_135_right;
  wire [9:0] _add_map_x_135_down;
  wire [9:0] _add_map_x_135_left;
  wire [9:0] _add_map_x_135_start;
  wire [9:0] _add_map_x_135_goal;
  wire [9:0] _add_map_x_135_now;
  wire [9:0] _add_map_x_135_data_out;
  wire [9:0] _add_map_x_135_data_out_index;
  wire [9:0] _add_map_x_135_data_near;
  wire _add_map_x_135_wall_t_out;
  wire [9:0] _add_map_x_135_data_org;
  wire [9:0] _add_map_x_135_data_org_near;
  wire [1:0] _add_map_x_135_s_g;
  wire [1:0] _add_map_x_135_s_g_near;
  wire _add_map_x_135_add_exe;
  wire _add_map_x_135_p_reset;
  wire _add_map_x_135_m_clock;
  wire [9:0] _add_map_x_134_moto_org_near;
  wire [9:0] _add_map_x_134_moto_org_near1;
  wire [9:0] _add_map_x_134_moto_org_near2;
  wire [9:0] _add_map_x_134_moto_org_near3;
  wire [9:0] _add_map_x_134_moto_org;
  wire [1:0] _add_map_x_134_sg_up;
  wire [1:0] _add_map_x_134_sg_down;
  wire [1:0] _add_map_x_134_sg_left;
  wire [1:0] _add_map_x_134_sg_right;
  wire _add_map_x_134_wall_t_in;
  wire [9:0] _add_map_x_134_moto;
  wire [9:0] _add_map_x_134_up;
  wire [9:0] _add_map_x_134_right;
  wire [9:0] _add_map_x_134_down;
  wire [9:0] _add_map_x_134_left;
  wire [9:0] _add_map_x_134_start;
  wire [9:0] _add_map_x_134_goal;
  wire [9:0] _add_map_x_134_now;
  wire [9:0] _add_map_x_134_data_out;
  wire [9:0] _add_map_x_134_data_out_index;
  wire [9:0] _add_map_x_134_data_near;
  wire _add_map_x_134_wall_t_out;
  wire [9:0] _add_map_x_134_data_org;
  wire [9:0] _add_map_x_134_data_org_near;
  wire [1:0] _add_map_x_134_s_g;
  wire [1:0] _add_map_x_134_s_g_near;
  wire _add_map_x_134_add_exe;
  wire _add_map_x_134_p_reset;
  wire _add_map_x_134_m_clock;
  wire [9:0] _add_map_x_133_moto_org_near;
  wire [9:0] _add_map_x_133_moto_org_near1;
  wire [9:0] _add_map_x_133_moto_org_near2;
  wire [9:0] _add_map_x_133_moto_org_near3;
  wire [9:0] _add_map_x_133_moto_org;
  wire [1:0] _add_map_x_133_sg_up;
  wire [1:0] _add_map_x_133_sg_down;
  wire [1:0] _add_map_x_133_sg_left;
  wire [1:0] _add_map_x_133_sg_right;
  wire _add_map_x_133_wall_t_in;
  wire [9:0] _add_map_x_133_moto;
  wire [9:0] _add_map_x_133_up;
  wire [9:0] _add_map_x_133_right;
  wire [9:0] _add_map_x_133_down;
  wire [9:0] _add_map_x_133_left;
  wire [9:0] _add_map_x_133_start;
  wire [9:0] _add_map_x_133_goal;
  wire [9:0] _add_map_x_133_now;
  wire [9:0] _add_map_x_133_data_out;
  wire [9:0] _add_map_x_133_data_out_index;
  wire [9:0] _add_map_x_133_data_near;
  wire _add_map_x_133_wall_t_out;
  wire [9:0] _add_map_x_133_data_org;
  wire [9:0] _add_map_x_133_data_org_near;
  wire [1:0] _add_map_x_133_s_g;
  wire [1:0] _add_map_x_133_s_g_near;
  wire _add_map_x_133_add_exe;
  wire _add_map_x_133_p_reset;
  wire _add_map_x_133_m_clock;
  wire [9:0] _add_map_x_132_moto_org_near;
  wire [9:0] _add_map_x_132_moto_org_near1;
  wire [9:0] _add_map_x_132_moto_org_near2;
  wire [9:0] _add_map_x_132_moto_org_near3;
  wire [9:0] _add_map_x_132_moto_org;
  wire [1:0] _add_map_x_132_sg_up;
  wire [1:0] _add_map_x_132_sg_down;
  wire [1:0] _add_map_x_132_sg_left;
  wire [1:0] _add_map_x_132_sg_right;
  wire _add_map_x_132_wall_t_in;
  wire [9:0] _add_map_x_132_moto;
  wire [9:0] _add_map_x_132_up;
  wire [9:0] _add_map_x_132_right;
  wire [9:0] _add_map_x_132_down;
  wire [9:0] _add_map_x_132_left;
  wire [9:0] _add_map_x_132_start;
  wire [9:0] _add_map_x_132_goal;
  wire [9:0] _add_map_x_132_now;
  wire [9:0] _add_map_x_132_data_out;
  wire [9:0] _add_map_x_132_data_out_index;
  wire [9:0] _add_map_x_132_data_near;
  wire _add_map_x_132_wall_t_out;
  wire [9:0] _add_map_x_132_data_org;
  wire [9:0] _add_map_x_132_data_org_near;
  wire [1:0] _add_map_x_132_s_g;
  wire [1:0] _add_map_x_132_s_g_near;
  wire _add_map_x_132_add_exe;
  wire _add_map_x_132_p_reset;
  wire _add_map_x_132_m_clock;
  wire [9:0] _add_map_x_131_moto_org_near;
  wire [9:0] _add_map_x_131_moto_org_near1;
  wire [9:0] _add_map_x_131_moto_org_near2;
  wire [9:0] _add_map_x_131_moto_org_near3;
  wire [9:0] _add_map_x_131_moto_org;
  wire [1:0] _add_map_x_131_sg_up;
  wire [1:0] _add_map_x_131_sg_down;
  wire [1:0] _add_map_x_131_sg_left;
  wire [1:0] _add_map_x_131_sg_right;
  wire _add_map_x_131_wall_t_in;
  wire [9:0] _add_map_x_131_moto;
  wire [9:0] _add_map_x_131_up;
  wire [9:0] _add_map_x_131_right;
  wire [9:0] _add_map_x_131_down;
  wire [9:0] _add_map_x_131_left;
  wire [9:0] _add_map_x_131_start;
  wire [9:0] _add_map_x_131_goal;
  wire [9:0] _add_map_x_131_now;
  wire [9:0] _add_map_x_131_data_out;
  wire [9:0] _add_map_x_131_data_out_index;
  wire [9:0] _add_map_x_131_data_near;
  wire _add_map_x_131_wall_t_out;
  wire [9:0] _add_map_x_131_data_org;
  wire [9:0] _add_map_x_131_data_org_near;
  wire [1:0] _add_map_x_131_s_g;
  wire [1:0] _add_map_x_131_s_g_near;
  wire _add_map_x_131_add_exe;
  wire _add_map_x_131_p_reset;
  wire _add_map_x_131_m_clock;
  wire [9:0] _add_map_x_130_moto_org_near;
  wire [9:0] _add_map_x_130_moto_org_near1;
  wire [9:0] _add_map_x_130_moto_org_near2;
  wire [9:0] _add_map_x_130_moto_org_near3;
  wire [9:0] _add_map_x_130_moto_org;
  wire [1:0] _add_map_x_130_sg_up;
  wire [1:0] _add_map_x_130_sg_down;
  wire [1:0] _add_map_x_130_sg_left;
  wire [1:0] _add_map_x_130_sg_right;
  wire _add_map_x_130_wall_t_in;
  wire [9:0] _add_map_x_130_moto;
  wire [9:0] _add_map_x_130_up;
  wire [9:0] _add_map_x_130_right;
  wire [9:0] _add_map_x_130_down;
  wire [9:0] _add_map_x_130_left;
  wire [9:0] _add_map_x_130_start;
  wire [9:0] _add_map_x_130_goal;
  wire [9:0] _add_map_x_130_now;
  wire [9:0] _add_map_x_130_data_out;
  wire [9:0] _add_map_x_130_data_out_index;
  wire [9:0] _add_map_x_130_data_near;
  wire _add_map_x_130_wall_t_out;
  wire [9:0] _add_map_x_130_data_org;
  wire [9:0] _add_map_x_130_data_org_near;
  wire [1:0] _add_map_x_130_s_g;
  wire [1:0] _add_map_x_130_s_g_near;
  wire _add_map_x_130_add_exe;
  wire _add_map_x_130_p_reset;
  wire _add_map_x_130_m_clock;
  wire [9:0] _add_map_x_129_moto_org_near;
  wire [9:0] _add_map_x_129_moto_org_near1;
  wire [9:0] _add_map_x_129_moto_org_near2;
  wire [9:0] _add_map_x_129_moto_org_near3;
  wire [9:0] _add_map_x_129_moto_org;
  wire [1:0] _add_map_x_129_sg_up;
  wire [1:0] _add_map_x_129_sg_down;
  wire [1:0] _add_map_x_129_sg_left;
  wire [1:0] _add_map_x_129_sg_right;
  wire _add_map_x_129_wall_t_in;
  wire [9:0] _add_map_x_129_moto;
  wire [9:0] _add_map_x_129_up;
  wire [9:0] _add_map_x_129_right;
  wire [9:0] _add_map_x_129_down;
  wire [9:0] _add_map_x_129_left;
  wire [9:0] _add_map_x_129_start;
  wire [9:0] _add_map_x_129_goal;
  wire [9:0] _add_map_x_129_now;
  wire [9:0] _add_map_x_129_data_out;
  wire [9:0] _add_map_x_129_data_out_index;
  wire [9:0] _add_map_x_129_data_near;
  wire _add_map_x_129_wall_t_out;
  wire [9:0] _add_map_x_129_data_org;
  wire [9:0] _add_map_x_129_data_org_near;
  wire [1:0] _add_map_x_129_s_g;
  wire [1:0] _add_map_x_129_s_g_near;
  wire _add_map_x_129_add_exe;
  wire _add_map_x_129_p_reset;
  wire _add_map_x_129_m_clock;
  wire [9:0] _add_map_x_128_moto_org_near;
  wire [9:0] _add_map_x_128_moto_org_near1;
  wire [9:0] _add_map_x_128_moto_org_near2;
  wire [9:0] _add_map_x_128_moto_org_near3;
  wire [9:0] _add_map_x_128_moto_org;
  wire [1:0] _add_map_x_128_sg_up;
  wire [1:0] _add_map_x_128_sg_down;
  wire [1:0] _add_map_x_128_sg_left;
  wire [1:0] _add_map_x_128_sg_right;
  wire _add_map_x_128_wall_t_in;
  wire [9:0] _add_map_x_128_moto;
  wire [9:0] _add_map_x_128_up;
  wire [9:0] _add_map_x_128_right;
  wire [9:0] _add_map_x_128_down;
  wire [9:0] _add_map_x_128_left;
  wire [9:0] _add_map_x_128_start;
  wire [9:0] _add_map_x_128_goal;
  wire [9:0] _add_map_x_128_now;
  wire [9:0] _add_map_x_128_data_out;
  wire [9:0] _add_map_x_128_data_out_index;
  wire [9:0] _add_map_x_128_data_near;
  wire _add_map_x_128_wall_t_out;
  wire [9:0] _add_map_x_128_data_org;
  wire [9:0] _add_map_x_128_data_org_near;
  wire [1:0] _add_map_x_128_s_g;
  wire [1:0] _add_map_x_128_s_g_near;
  wire _add_map_x_128_add_exe;
  wire _add_map_x_128_p_reset;
  wire _add_map_x_128_m_clock;
  wire [9:0] _add_map_x_127_moto_org_near;
  wire [9:0] _add_map_x_127_moto_org_near1;
  wire [9:0] _add_map_x_127_moto_org_near2;
  wire [9:0] _add_map_x_127_moto_org_near3;
  wire [9:0] _add_map_x_127_moto_org;
  wire [1:0] _add_map_x_127_sg_up;
  wire [1:0] _add_map_x_127_sg_down;
  wire [1:0] _add_map_x_127_sg_left;
  wire [1:0] _add_map_x_127_sg_right;
  wire _add_map_x_127_wall_t_in;
  wire [9:0] _add_map_x_127_moto;
  wire [9:0] _add_map_x_127_up;
  wire [9:0] _add_map_x_127_right;
  wire [9:0] _add_map_x_127_down;
  wire [9:0] _add_map_x_127_left;
  wire [9:0] _add_map_x_127_start;
  wire [9:0] _add_map_x_127_goal;
  wire [9:0] _add_map_x_127_now;
  wire [9:0] _add_map_x_127_data_out;
  wire [9:0] _add_map_x_127_data_out_index;
  wire [9:0] _add_map_x_127_data_near;
  wire _add_map_x_127_wall_t_out;
  wire [9:0] _add_map_x_127_data_org;
  wire [9:0] _add_map_x_127_data_org_near;
  wire [1:0] _add_map_x_127_s_g;
  wire [1:0] _add_map_x_127_s_g_near;
  wire _add_map_x_127_add_exe;
  wire _add_map_x_127_p_reset;
  wire _add_map_x_127_m_clock;
  wire [9:0] _add_map_x_126_moto_org_near;
  wire [9:0] _add_map_x_126_moto_org_near1;
  wire [9:0] _add_map_x_126_moto_org_near2;
  wire [9:0] _add_map_x_126_moto_org_near3;
  wire [9:0] _add_map_x_126_moto_org;
  wire [1:0] _add_map_x_126_sg_up;
  wire [1:0] _add_map_x_126_sg_down;
  wire [1:0] _add_map_x_126_sg_left;
  wire [1:0] _add_map_x_126_sg_right;
  wire _add_map_x_126_wall_t_in;
  wire [9:0] _add_map_x_126_moto;
  wire [9:0] _add_map_x_126_up;
  wire [9:0] _add_map_x_126_right;
  wire [9:0] _add_map_x_126_down;
  wire [9:0] _add_map_x_126_left;
  wire [9:0] _add_map_x_126_start;
  wire [9:0] _add_map_x_126_goal;
  wire [9:0] _add_map_x_126_now;
  wire [9:0] _add_map_x_126_data_out;
  wire [9:0] _add_map_x_126_data_out_index;
  wire [9:0] _add_map_x_126_data_near;
  wire _add_map_x_126_wall_t_out;
  wire [9:0] _add_map_x_126_data_org;
  wire [9:0] _add_map_x_126_data_org_near;
  wire [1:0] _add_map_x_126_s_g;
  wire [1:0] _add_map_x_126_s_g_near;
  wire _add_map_x_126_add_exe;
  wire _add_map_x_126_p_reset;
  wire _add_map_x_126_m_clock;
  wire [9:0] _add_map_x_125_moto_org_near;
  wire [9:0] _add_map_x_125_moto_org_near1;
  wire [9:0] _add_map_x_125_moto_org_near2;
  wire [9:0] _add_map_x_125_moto_org_near3;
  wire [9:0] _add_map_x_125_moto_org;
  wire [1:0] _add_map_x_125_sg_up;
  wire [1:0] _add_map_x_125_sg_down;
  wire [1:0] _add_map_x_125_sg_left;
  wire [1:0] _add_map_x_125_sg_right;
  wire _add_map_x_125_wall_t_in;
  wire [9:0] _add_map_x_125_moto;
  wire [9:0] _add_map_x_125_up;
  wire [9:0] _add_map_x_125_right;
  wire [9:0] _add_map_x_125_down;
  wire [9:0] _add_map_x_125_left;
  wire [9:0] _add_map_x_125_start;
  wire [9:0] _add_map_x_125_goal;
  wire [9:0] _add_map_x_125_now;
  wire [9:0] _add_map_x_125_data_out;
  wire [9:0] _add_map_x_125_data_out_index;
  wire [9:0] _add_map_x_125_data_near;
  wire _add_map_x_125_wall_t_out;
  wire [9:0] _add_map_x_125_data_org;
  wire [9:0] _add_map_x_125_data_org_near;
  wire [1:0] _add_map_x_125_s_g;
  wire [1:0] _add_map_x_125_s_g_near;
  wire _add_map_x_125_add_exe;
  wire _add_map_x_125_p_reset;
  wire _add_map_x_125_m_clock;
  wire [9:0] _add_map_x_124_moto_org_near;
  wire [9:0] _add_map_x_124_moto_org_near1;
  wire [9:0] _add_map_x_124_moto_org_near2;
  wire [9:0] _add_map_x_124_moto_org_near3;
  wire [9:0] _add_map_x_124_moto_org;
  wire [1:0] _add_map_x_124_sg_up;
  wire [1:0] _add_map_x_124_sg_down;
  wire [1:0] _add_map_x_124_sg_left;
  wire [1:0] _add_map_x_124_sg_right;
  wire _add_map_x_124_wall_t_in;
  wire [9:0] _add_map_x_124_moto;
  wire [9:0] _add_map_x_124_up;
  wire [9:0] _add_map_x_124_right;
  wire [9:0] _add_map_x_124_down;
  wire [9:0] _add_map_x_124_left;
  wire [9:0] _add_map_x_124_start;
  wire [9:0] _add_map_x_124_goal;
  wire [9:0] _add_map_x_124_now;
  wire [9:0] _add_map_x_124_data_out;
  wire [9:0] _add_map_x_124_data_out_index;
  wire [9:0] _add_map_x_124_data_near;
  wire _add_map_x_124_wall_t_out;
  wire [9:0] _add_map_x_124_data_org;
  wire [9:0] _add_map_x_124_data_org_near;
  wire [1:0] _add_map_x_124_s_g;
  wire [1:0] _add_map_x_124_s_g_near;
  wire _add_map_x_124_add_exe;
  wire _add_map_x_124_p_reset;
  wire _add_map_x_124_m_clock;
  wire [9:0] _add_map_x_123_moto_org_near;
  wire [9:0] _add_map_x_123_moto_org_near1;
  wire [9:0] _add_map_x_123_moto_org_near2;
  wire [9:0] _add_map_x_123_moto_org_near3;
  wire [9:0] _add_map_x_123_moto_org;
  wire [1:0] _add_map_x_123_sg_up;
  wire [1:0] _add_map_x_123_sg_down;
  wire [1:0] _add_map_x_123_sg_left;
  wire [1:0] _add_map_x_123_sg_right;
  wire _add_map_x_123_wall_t_in;
  wire [9:0] _add_map_x_123_moto;
  wire [9:0] _add_map_x_123_up;
  wire [9:0] _add_map_x_123_right;
  wire [9:0] _add_map_x_123_down;
  wire [9:0] _add_map_x_123_left;
  wire [9:0] _add_map_x_123_start;
  wire [9:0] _add_map_x_123_goal;
  wire [9:0] _add_map_x_123_now;
  wire [9:0] _add_map_x_123_data_out;
  wire [9:0] _add_map_x_123_data_out_index;
  wire [9:0] _add_map_x_123_data_near;
  wire _add_map_x_123_wall_t_out;
  wire [9:0] _add_map_x_123_data_org;
  wire [9:0] _add_map_x_123_data_org_near;
  wire [1:0] _add_map_x_123_s_g;
  wire [1:0] _add_map_x_123_s_g_near;
  wire _add_map_x_123_add_exe;
  wire _add_map_x_123_p_reset;
  wire _add_map_x_123_m_clock;
  wire [9:0] _add_map_x_122_moto_org_near;
  wire [9:0] _add_map_x_122_moto_org_near1;
  wire [9:0] _add_map_x_122_moto_org_near2;
  wire [9:0] _add_map_x_122_moto_org_near3;
  wire [9:0] _add_map_x_122_moto_org;
  wire [1:0] _add_map_x_122_sg_up;
  wire [1:0] _add_map_x_122_sg_down;
  wire [1:0] _add_map_x_122_sg_left;
  wire [1:0] _add_map_x_122_sg_right;
  wire _add_map_x_122_wall_t_in;
  wire [9:0] _add_map_x_122_moto;
  wire [9:0] _add_map_x_122_up;
  wire [9:0] _add_map_x_122_right;
  wire [9:0] _add_map_x_122_down;
  wire [9:0] _add_map_x_122_left;
  wire [9:0] _add_map_x_122_start;
  wire [9:0] _add_map_x_122_goal;
  wire [9:0] _add_map_x_122_now;
  wire [9:0] _add_map_x_122_data_out;
  wire [9:0] _add_map_x_122_data_out_index;
  wire [9:0] _add_map_x_122_data_near;
  wire _add_map_x_122_wall_t_out;
  wire [9:0] _add_map_x_122_data_org;
  wire [9:0] _add_map_x_122_data_org_near;
  wire [1:0] _add_map_x_122_s_g;
  wire [1:0] _add_map_x_122_s_g_near;
  wire _add_map_x_122_add_exe;
  wire _add_map_x_122_p_reset;
  wire _add_map_x_122_m_clock;
  wire [9:0] _add_map_x_121_moto_org_near;
  wire [9:0] _add_map_x_121_moto_org_near1;
  wire [9:0] _add_map_x_121_moto_org_near2;
  wire [9:0] _add_map_x_121_moto_org_near3;
  wire [9:0] _add_map_x_121_moto_org;
  wire [1:0] _add_map_x_121_sg_up;
  wire [1:0] _add_map_x_121_sg_down;
  wire [1:0] _add_map_x_121_sg_left;
  wire [1:0] _add_map_x_121_sg_right;
  wire _add_map_x_121_wall_t_in;
  wire [9:0] _add_map_x_121_moto;
  wire [9:0] _add_map_x_121_up;
  wire [9:0] _add_map_x_121_right;
  wire [9:0] _add_map_x_121_down;
  wire [9:0] _add_map_x_121_left;
  wire [9:0] _add_map_x_121_start;
  wire [9:0] _add_map_x_121_goal;
  wire [9:0] _add_map_x_121_now;
  wire [9:0] _add_map_x_121_data_out;
  wire [9:0] _add_map_x_121_data_out_index;
  wire [9:0] _add_map_x_121_data_near;
  wire _add_map_x_121_wall_t_out;
  wire [9:0] _add_map_x_121_data_org;
  wire [9:0] _add_map_x_121_data_org_near;
  wire [1:0] _add_map_x_121_s_g;
  wire [1:0] _add_map_x_121_s_g_near;
  wire _add_map_x_121_add_exe;
  wire _add_map_x_121_p_reset;
  wire _add_map_x_121_m_clock;
  wire [9:0] _add_map_x_120_moto_org_near;
  wire [9:0] _add_map_x_120_moto_org_near1;
  wire [9:0] _add_map_x_120_moto_org_near2;
  wire [9:0] _add_map_x_120_moto_org_near3;
  wire [9:0] _add_map_x_120_moto_org;
  wire [1:0] _add_map_x_120_sg_up;
  wire [1:0] _add_map_x_120_sg_down;
  wire [1:0] _add_map_x_120_sg_left;
  wire [1:0] _add_map_x_120_sg_right;
  wire _add_map_x_120_wall_t_in;
  wire [9:0] _add_map_x_120_moto;
  wire [9:0] _add_map_x_120_up;
  wire [9:0] _add_map_x_120_right;
  wire [9:0] _add_map_x_120_down;
  wire [9:0] _add_map_x_120_left;
  wire [9:0] _add_map_x_120_start;
  wire [9:0] _add_map_x_120_goal;
  wire [9:0] _add_map_x_120_now;
  wire [9:0] _add_map_x_120_data_out;
  wire [9:0] _add_map_x_120_data_out_index;
  wire [9:0] _add_map_x_120_data_near;
  wire _add_map_x_120_wall_t_out;
  wire [9:0] _add_map_x_120_data_org;
  wire [9:0] _add_map_x_120_data_org_near;
  wire [1:0] _add_map_x_120_s_g;
  wire [1:0] _add_map_x_120_s_g_near;
  wire _add_map_x_120_add_exe;
  wire _add_map_x_120_p_reset;
  wire _add_map_x_120_m_clock;
  wire [9:0] _add_map_x_119_moto_org_near;
  wire [9:0] _add_map_x_119_moto_org_near1;
  wire [9:0] _add_map_x_119_moto_org_near2;
  wire [9:0] _add_map_x_119_moto_org_near3;
  wire [9:0] _add_map_x_119_moto_org;
  wire [1:0] _add_map_x_119_sg_up;
  wire [1:0] _add_map_x_119_sg_down;
  wire [1:0] _add_map_x_119_sg_left;
  wire [1:0] _add_map_x_119_sg_right;
  wire _add_map_x_119_wall_t_in;
  wire [9:0] _add_map_x_119_moto;
  wire [9:0] _add_map_x_119_up;
  wire [9:0] _add_map_x_119_right;
  wire [9:0] _add_map_x_119_down;
  wire [9:0] _add_map_x_119_left;
  wire [9:0] _add_map_x_119_start;
  wire [9:0] _add_map_x_119_goal;
  wire [9:0] _add_map_x_119_now;
  wire [9:0] _add_map_x_119_data_out;
  wire [9:0] _add_map_x_119_data_out_index;
  wire [9:0] _add_map_x_119_data_near;
  wire _add_map_x_119_wall_t_out;
  wire [9:0] _add_map_x_119_data_org;
  wire [9:0] _add_map_x_119_data_org_near;
  wire [1:0] _add_map_x_119_s_g;
  wire [1:0] _add_map_x_119_s_g_near;
  wire _add_map_x_119_add_exe;
  wire _add_map_x_119_p_reset;
  wire _add_map_x_119_m_clock;
  wire [9:0] _add_map_x_118_moto_org_near;
  wire [9:0] _add_map_x_118_moto_org_near1;
  wire [9:0] _add_map_x_118_moto_org_near2;
  wire [9:0] _add_map_x_118_moto_org_near3;
  wire [9:0] _add_map_x_118_moto_org;
  wire [1:0] _add_map_x_118_sg_up;
  wire [1:0] _add_map_x_118_sg_down;
  wire [1:0] _add_map_x_118_sg_left;
  wire [1:0] _add_map_x_118_sg_right;
  wire _add_map_x_118_wall_t_in;
  wire [9:0] _add_map_x_118_moto;
  wire [9:0] _add_map_x_118_up;
  wire [9:0] _add_map_x_118_right;
  wire [9:0] _add_map_x_118_down;
  wire [9:0] _add_map_x_118_left;
  wire [9:0] _add_map_x_118_start;
  wire [9:0] _add_map_x_118_goal;
  wire [9:0] _add_map_x_118_now;
  wire [9:0] _add_map_x_118_data_out;
  wire [9:0] _add_map_x_118_data_out_index;
  wire [9:0] _add_map_x_118_data_near;
  wire _add_map_x_118_wall_t_out;
  wire [9:0] _add_map_x_118_data_org;
  wire [9:0] _add_map_x_118_data_org_near;
  wire [1:0] _add_map_x_118_s_g;
  wire [1:0] _add_map_x_118_s_g_near;
  wire _add_map_x_118_add_exe;
  wire _add_map_x_118_p_reset;
  wire _add_map_x_118_m_clock;
  wire [9:0] _add_map_x_117_moto_org_near;
  wire [9:0] _add_map_x_117_moto_org_near1;
  wire [9:0] _add_map_x_117_moto_org_near2;
  wire [9:0] _add_map_x_117_moto_org_near3;
  wire [9:0] _add_map_x_117_moto_org;
  wire [1:0] _add_map_x_117_sg_up;
  wire [1:0] _add_map_x_117_sg_down;
  wire [1:0] _add_map_x_117_sg_left;
  wire [1:0] _add_map_x_117_sg_right;
  wire _add_map_x_117_wall_t_in;
  wire [9:0] _add_map_x_117_moto;
  wire [9:0] _add_map_x_117_up;
  wire [9:0] _add_map_x_117_right;
  wire [9:0] _add_map_x_117_down;
  wire [9:0] _add_map_x_117_left;
  wire [9:0] _add_map_x_117_start;
  wire [9:0] _add_map_x_117_goal;
  wire [9:0] _add_map_x_117_now;
  wire [9:0] _add_map_x_117_data_out;
  wire [9:0] _add_map_x_117_data_out_index;
  wire [9:0] _add_map_x_117_data_near;
  wire _add_map_x_117_wall_t_out;
  wire [9:0] _add_map_x_117_data_org;
  wire [9:0] _add_map_x_117_data_org_near;
  wire [1:0] _add_map_x_117_s_g;
  wire [1:0] _add_map_x_117_s_g_near;
  wire _add_map_x_117_add_exe;
  wire _add_map_x_117_p_reset;
  wire _add_map_x_117_m_clock;
  wire [9:0] _add_map_x_116_moto_org_near;
  wire [9:0] _add_map_x_116_moto_org_near1;
  wire [9:0] _add_map_x_116_moto_org_near2;
  wire [9:0] _add_map_x_116_moto_org_near3;
  wire [9:0] _add_map_x_116_moto_org;
  wire [1:0] _add_map_x_116_sg_up;
  wire [1:0] _add_map_x_116_sg_down;
  wire [1:0] _add_map_x_116_sg_left;
  wire [1:0] _add_map_x_116_sg_right;
  wire _add_map_x_116_wall_t_in;
  wire [9:0] _add_map_x_116_moto;
  wire [9:0] _add_map_x_116_up;
  wire [9:0] _add_map_x_116_right;
  wire [9:0] _add_map_x_116_down;
  wire [9:0] _add_map_x_116_left;
  wire [9:0] _add_map_x_116_start;
  wire [9:0] _add_map_x_116_goal;
  wire [9:0] _add_map_x_116_now;
  wire [9:0] _add_map_x_116_data_out;
  wire [9:0] _add_map_x_116_data_out_index;
  wire [9:0] _add_map_x_116_data_near;
  wire _add_map_x_116_wall_t_out;
  wire [9:0] _add_map_x_116_data_org;
  wire [9:0] _add_map_x_116_data_org_near;
  wire [1:0] _add_map_x_116_s_g;
  wire [1:0] _add_map_x_116_s_g_near;
  wire _add_map_x_116_add_exe;
  wire _add_map_x_116_p_reset;
  wire _add_map_x_116_m_clock;
  wire [9:0] _add_map_x_115_moto_org_near;
  wire [9:0] _add_map_x_115_moto_org_near1;
  wire [9:0] _add_map_x_115_moto_org_near2;
  wire [9:0] _add_map_x_115_moto_org_near3;
  wire [9:0] _add_map_x_115_moto_org;
  wire [1:0] _add_map_x_115_sg_up;
  wire [1:0] _add_map_x_115_sg_down;
  wire [1:0] _add_map_x_115_sg_left;
  wire [1:0] _add_map_x_115_sg_right;
  wire _add_map_x_115_wall_t_in;
  wire [9:0] _add_map_x_115_moto;
  wire [9:0] _add_map_x_115_up;
  wire [9:0] _add_map_x_115_right;
  wire [9:0] _add_map_x_115_down;
  wire [9:0] _add_map_x_115_left;
  wire [9:0] _add_map_x_115_start;
  wire [9:0] _add_map_x_115_goal;
  wire [9:0] _add_map_x_115_now;
  wire [9:0] _add_map_x_115_data_out;
  wire [9:0] _add_map_x_115_data_out_index;
  wire [9:0] _add_map_x_115_data_near;
  wire _add_map_x_115_wall_t_out;
  wire [9:0] _add_map_x_115_data_org;
  wire [9:0] _add_map_x_115_data_org_near;
  wire [1:0] _add_map_x_115_s_g;
  wire [1:0] _add_map_x_115_s_g_near;
  wire _add_map_x_115_add_exe;
  wire _add_map_x_115_p_reset;
  wire _add_map_x_115_m_clock;
  wire [9:0] _add_map_x_114_moto_org_near;
  wire [9:0] _add_map_x_114_moto_org_near1;
  wire [9:0] _add_map_x_114_moto_org_near2;
  wire [9:0] _add_map_x_114_moto_org_near3;
  wire [9:0] _add_map_x_114_moto_org;
  wire [1:0] _add_map_x_114_sg_up;
  wire [1:0] _add_map_x_114_sg_down;
  wire [1:0] _add_map_x_114_sg_left;
  wire [1:0] _add_map_x_114_sg_right;
  wire _add_map_x_114_wall_t_in;
  wire [9:0] _add_map_x_114_moto;
  wire [9:0] _add_map_x_114_up;
  wire [9:0] _add_map_x_114_right;
  wire [9:0] _add_map_x_114_down;
  wire [9:0] _add_map_x_114_left;
  wire [9:0] _add_map_x_114_start;
  wire [9:0] _add_map_x_114_goal;
  wire [9:0] _add_map_x_114_now;
  wire [9:0] _add_map_x_114_data_out;
  wire [9:0] _add_map_x_114_data_out_index;
  wire [9:0] _add_map_x_114_data_near;
  wire _add_map_x_114_wall_t_out;
  wire [9:0] _add_map_x_114_data_org;
  wire [9:0] _add_map_x_114_data_org_near;
  wire [1:0] _add_map_x_114_s_g;
  wire [1:0] _add_map_x_114_s_g_near;
  wire _add_map_x_114_add_exe;
  wire _add_map_x_114_p_reset;
  wire _add_map_x_114_m_clock;
  wire [9:0] _add_map_x_113_moto_org_near;
  wire [9:0] _add_map_x_113_moto_org_near1;
  wire [9:0] _add_map_x_113_moto_org_near2;
  wire [9:0] _add_map_x_113_moto_org_near3;
  wire [9:0] _add_map_x_113_moto_org;
  wire [1:0] _add_map_x_113_sg_up;
  wire [1:0] _add_map_x_113_sg_down;
  wire [1:0] _add_map_x_113_sg_left;
  wire [1:0] _add_map_x_113_sg_right;
  wire _add_map_x_113_wall_t_in;
  wire [9:0] _add_map_x_113_moto;
  wire [9:0] _add_map_x_113_up;
  wire [9:0] _add_map_x_113_right;
  wire [9:0] _add_map_x_113_down;
  wire [9:0] _add_map_x_113_left;
  wire [9:0] _add_map_x_113_start;
  wire [9:0] _add_map_x_113_goal;
  wire [9:0] _add_map_x_113_now;
  wire [9:0] _add_map_x_113_data_out;
  wire [9:0] _add_map_x_113_data_out_index;
  wire [9:0] _add_map_x_113_data_near;
  wire _add_map_x_113_wall_t_out;
  wire [9:0] _add_map_x_113_data_org;
  wire [9:0] _add_map_x_113_data_org_near;
  wire [1:0] _add_map_x_113_s_g;
  wire [1:0] _add_map_x_113_s_g_near;
  wire _add_map_x_113_add_exe;
  wire _add_map_x_113_p_reset;
  wire _add_map_x_113_m_clock;
  wire [9:0] _add_map_x_112_moto_org_near;
  wire [9:0] _add_map_x_112_moto_org_near1;
  wire [9:0] _add_map_x_112_moto_org_near2;
  wire [9:0] _add_map_x_112_moto_org_near3;
  wire [9:0] _add_map_x_112_moto_org;
  wire [1:0] _add_map_x_112_sg_up;
  wire [1:0] _add_map_x_112_sg_down;
  wire [1:0] _add_map_x_112_sg_left;
  wire [1:0] _add_map_x_112_sg_right;
  wire _add_map_x_112_wall_t_in;
  wire [9:0] _add_map_x_112_moto;
  wire [9:0] _add_map_x_112_up;
  wire [9:0] _add_map_x_112_right;
  wire [9:0] _add_map_x_112_down;
  wire [9:0] _add_map_x_112_left;
  wire [9:0] _add_map_x_112_start;
  wire [9:0] _add_map_x_112_goal;
  wire [9:0] _add_map_x_112_now;
  wire [9:0] _add_map_x_112_data_out;
  wire [9:0] _add_map_x_112_data_out_index;
  wire [9:0] _add_map_x_112_data_near;
  wire _add_map_x_112_wall_t_out;
  wire [9:0] _add_map_x_112_data_org;
  wire [9:0] _add_map_x_112_data_org_near;
  wire [1:0] _add_map_x_112_s_g;
  wire [1:0] _add_map_x_112_s_g_near;
  wire _add_map_x_112_add_exe;
  wire _add_map_x_112_p_reset;
  wire _add_map_x_112_m_clock;
  wire [9:0] _add_map_x_111_moto_org_near;
  wire [9:0] _add_map_x_111_moto_org_near1;
  wire [9:0] _add_map_x_111_moto_org_near2;
  wire [9:0] _add_map_x_111_moto_org_near3;
  wire [9:0] _add_map_x_111_moto_org;
  wire [1:0] _add_map_x_111_sg_up;
  wire [1:0] _add_map_x_111_sg_down;
  wire [1:0] _add_map_x_111_sg_left;
  wire [1:0] _add_map_x_111_sg_right;
  wire _add_map_x_111_wall_t_in;
  wire [9:0] _add_map_x_111_moto;
  wire [9:0] _add_map_x_111_up;
  wire [9:0] _add_map_x_111_right;
  wire [9:0] _add_map_x_111_down;
  wire [9:0] _add_map_x_111_left;
  wire [9:0] _add_map_x_111_start;
  wire [9:0] _add_map_x_111_goal;
  wire [9:0] _add_map_x_111_now;
  wire [9:0] _add_map_x_111_data_out;
  wire [9:0] _add_map_x_111_data_out_index;
  wire [9:0] _add_map_x_111_data_near;
  wire _add_map_x_111_wall_t_out;
  wire [9:0] _add_map_x_111_data_org;
  wire [9:0] _add_map_x_111_data_org_near;
  wire [1:0] _add_map_x_111_s_g;
  wire [1:0] _add_map_x_111_s_g_near;
  wire _add_map_x_111_add_exe;
  wire _add_map_x_111_p_reset;
  wire _add_map_x_111_m_clock;
  wire [9:0] _add_map_x_110_moto_org_near;
  wire [9:0] _add_map_x_110_moto_org_near1;
  wire [9:0] _add_map_x_110_moto_org_near2;
  wire [9:0] _add_map_x_110_moto_org_near3;
  wire [9:0] _add_map_x_110_moto_org;
  wire [1:0] _add_map_x_110_sg_up;
  wire [1:0] _add_map_x_110_sg_down;
  wire [1:0] _add_map_x_110_sg_left;
  wire [1:0] _add_map_x_110_sg_right;
  wire _add_map_x_110_wall_t_in;
  wire [9:0] _add_map_x_110_moto;
  wire [9:0] _add_map_x_110_up;
  wire [9:0] _add_map_x_110_right;
  wire [9:0] _add_map_x_110_down;
  wire [9:0] _add_map_x_110_left;
  wire [9:0] _add_map_x_110_start;
  wire [9:0] _add_map_x_110_goal;
  wire [9:0] _add_map_x_110_now;
  wire [9:0] _add_map_x_110_data_out;
  wire [9:0] _add_map_x_110_data_out_index;
  wire [9:0] _add_map_x_110_data_near;
  wire _add_map_x_110_wall_t_out;
  wire [9:0] _add_map_x_110_data_org;
  wire [9:0] _add_map_x_110_data_org_near;
  wire [1:0] _add_map_x_110_s_g;
  wire [1:0] _add_map_x_110_s_g_near;
  wire _add_map_x_110_add_exe;
  wire _add_map_x_110_p_reset;
  wire _add_map_x_110_m_clock;
  wire [9:0] _add_map_x_109_moto_org_near;
  wire [9:0] _add_map_x_109_moto_org_near1;
  wire [9:0] _add_map_x_109_moto_org_near2;
  wire [9:0] _add_map_x_109_moto_org_near3;
  wire [9:0] _add_map_x_109_moto_org;
  wire [1:0] _add_map_x_109_sg_up;
  wire [1:0] _add_map_x_109_sg_down;
  wire [1:0] _add_map_x_109_sg_left;
  wire [1:0] _add_map_x_109_sg_right;
  wire _add_map_x_109_wall_t_in;
  wire [9:0] _add_map_x_109_moto;
  wire [9:0] _add_map_x_109_up;
  wire [9:0] _add_map_x_109_right;
  wire [9:0] _add_map_x_109_down;
  wire [9:0] _add_map_x_109_left;
  wire [9:0] _add_map_x_109_start;
  wire [9:0] _add_map_x_109_goal;
  wire [9:0] _add_map_x_109_now;
  wire [9:0] _add_map_x_109_data_out;
  wire [9:0] _add_map_x_109_data_out_index;
  wire [9:0] _add_map_x_109_data_near;
  wire _add_map_x_109_wall_t_out;
  wire [9:0] _add_map_x_109_data_org;
  wire [9:0] _add_map_x_109_data_org_near;
  wire [1:0] _add_map_x_109_s_g;
  wire [1:0] _add_map_x_109_s_g_near;
  wire _add_map_x_109_add_exe;
  wire _add_map_x_109_p_reset;
  wire _add_map_x_109_m_clock;
  wire [9:0] _add_map_x_108_moto_org_near;
  wire [9:0] _add_map_x_108_moto_org_near1;
  wire [9:0] _add_map_x_108_moto_org_near2;
  wire [9:0] _add_map_x_108_moto_org_near3;
  wire [9:0] _add_map_x_108_moto_org;
  wire [1:0] _add_map_x_108_sg_up;
  wire [1:0] _add_map_x_108_sg_down;
  wire [1:0] _add_map_x_108_sg_left;
  wire [1:0] _add_map_x_108_sg_right;
  wire _add_map_x_108_wall_t_in;
  wire [9:0] _add_map_x_108_moto;
  wire [9:0] _add_map_x_108_up;
  wire [9:0] _add_map_x_108_right;
  wire [9:0] _add_map_x_108_down;
  wire [9:0] _add_map_x_108_left;
  wire [9:0] _add_map_x_108_start;
  wire [9:0] _add_map_x_108_goal;
  wire [9:0] _add_map_x_108_now;
  wire [9:0] _add_map_x_108_data_out;
  wire [9:0] _add_map_x_108_data_out_index;
  wire [9:0] _add_map_x_108_data_near;
  wire _add_map_x_108_wall_t_out;
  wire [9:0] _add_map_x_108_data_org;
  wire [9:0] _add_map_x_108_data_org_near;
  wire [1:0] _add_map_x_108_s_g;
  wire [1:0] _add_map_x_108_s_g_near;
  wire _add_map_x_108_add_exe;
  wire _add_map_x_108_p_reset;
  wire _add_map_x_108_m_clock;
  wire [9:0] _add_map_x_107_moto_org_near;
  wire [9:0] _add_map_x_107_moto_org_near1;
  wire [9:0] _add_map_x_107_moto_org_near2;
  wire [9:0] _add_map_x_107_moto_org_near3;
  wire [9:0] _add_map_x_107_moto_org;
  wire [1:0] _add_map_x_107_sg_up;
  wire [1:0] _add_map_x_107_sg_down;
  wire [1:0] _add_map_x_107_sg_left;
  wire [1:0] _add_map_x_107_sg_right;
  wire _add_map_x_107_wall_t_in;
  wire [9:0] _add_map_x_107_moto;
  wire [9:0] _add_map_x_107_up;
  wire [9:0] _add_map_x_107_right;
  wire [9:0] _add_map_x_107_down;
  wire [9:0] _add_map_x_107_left;
  wire [9:0] _add_map_x_107_start;
  wire [9:0] _add_map_x_107_goal;
  wire [9:0] _add_map_x_107_now;
  wire [9:0] _add_map_x_107_data_out;
  wire [9:0] _add_map_x_107_data_out_index;
  wire [9:0] _add_map_x_107_data_near;
  wire _add_map_x_107_wall_t_out;
  wire [9:0] _add_map_x_107_data_org;
  wire [9:0] _add_map_x_107_data_org_near;
  wire [1:0] _add_map_x_107_s_g;
  wire [1:0] _add_map_x_107_s_g_near;
  wire _add_map_x_107_add_exe;
  wire _add_map_x_107_p_reset;
  wire _add_map_x_107_m_clock;
  wire [9:0] _add_map_x_106_moto_org_near;
  wire [9:0] _add_map_x_106_moto_org_near1;
  wire [9:0] _add_map_x_106_moto_org_near2;
  wire [9:0] _add_map_x_106_moto_org_near3;
  wire [9:0] _add_map_x_106_moto_org;
  wire [1:0] _add_map_x_106_sg_up;
  wire [1:0] _add_map_x_106_sg_down;
  wire [1:0] _add_map_x_106_sg_left;
  wire [1:0] _add_map_x_106_sg_right;
  wire _add_map_x_106_wall_t_in;
  wire [9:0] _add_map_x_106_moto;
  wire [9:0] _add_map_x_106_up;
  wire [9:0] _add_map_x_106_right;
  wire [9:0] _add_map_x_106_down;
  wire [9:0] _add_map_x_106_left;
  wire [9:0] _add_map_x_106_start;
  wire [9:0] _add_map_x_106_goal;
  wire [9:0] _add_map_x_106_now;
  wire [9:0] _add_map_x_106_data_out;
  wire [9:0] _add_map_x_106_data_out_index;
  wire [9:0] _add_map_x_106_data_near;
  wire _add_map_x_106_wall_t_out;
  wire [9:0] _add_map_x_106_data_org;
  wire [9:0] _add_map_x_106_data_org_near;
  wire [1:0] _add_map_x_106_s_g;
  wire [1:0] _add_map_x_106_s_g_near;
  wire _add_map_x_106_add_exe;
  wire _add_map_x_106_p_reset;
  wire _add_map_x_106_m_clock;
  wire [9:0] _add_map_x_105_moto_org_near;
  wire [9:0] _add_map_x_105_moto_org_near1;
  wire [9:0] _add_map_x_105_moto_org_near2;
  wire [9:0] _add_map_x_105_moto_org_near3;
  wire [9:0] _add_map_x_105_moto_org;
  wire [1:0] _add_map_x_105_sg_up;
  wire [1:0] _add_map_x_105_sg_down;
  wire [1:0] _add_map_x_105_sg_left;
  wire [1:0] _add_map_x_105_sg_right;
  wire _add_map_x_105_wall_t_in;
  wire [9:0] _add_map_x_105_moto;
  wire [9:0] _add_map_x_105_up;
  wire [9:0] _add_map_x_105_right;
  wire [9:0] _add_map_x_105_down;
  wire [9:0] _add_map_x_105_left;
  wire [9:0] _add_map_x_105_start;
  wire [9:0] _add_map_x_105_goal;
  wire [9:0] _add_map_x_105_now;
  wire [9:0] _add_map_x_105_data_out;
  wire [9:0] _add_map_x_105_data_out_index;
  wire [9:0] _add_map_x_105_data_near;
  wire _add_map_x_105_wall_t_out;
  wire [9:0] _add_map_x_105_data_org;
  wire [9:0] _add_map_x_105_data_org_near;
  wire [1:0] _add_map_x_105_s_g;
  wire [1:0] _add_map_x_105_s_g_near;
  wire _add_map_x_105_add_exe;
  wire _add_map_x_105_p_reset;
  wire _add_map_x_105_m_clock;
  wire [9:0] _add_map_x_104_moto_org_near;
  wire [9:0] _add_map_x_104_moto_org_near1;
  wire [9:0] _add_map_x_104_moto_org_near2;
  wire [9:0] _add_map_x_104_moto_org_near3;
  wire [9:0] _add_map_x_104_moto_org;
  wire [1:0] _add_map_x_104_sg_up;
  wire [1:0] _add_map_x_104_sg_down;
  wire [1:0] _add_map_x_104_sg_left;
  wire [1:0] _add_map_x_104_sg_right;
  wire _add_map_x_104_wall_t_in;
  wire [9:0] _add_map_x_104_moto;
  wire [9:0] _add_map_x_104_up;
  wire [9:0] _add_map_x_104_right;
  wire [9:0] _add_map_x_104_down;
  wire [9:0] _add_map_x_104_left;
  wire [9:0] _add_map_x_104_start;
  wire [9:0] _add_map_x_104_goal;
  wire [9:0] _add_map_x_104_now;
  wire [9:0] _add_map_x_104_data_out;
  wire [9:0] _add_map_x_104_data_out_index;
  wire [9:0] _add_map_x_104_data_near;
  wire _add_map_x_104_wall_t_out;
  wire [9:0] _add_map_x_104_data_org;
  wire [9:0] _add_map_x_104_data_org_near;
  wire [1:0] _add_map_x_104_s_g;
  wire [1:0] _add_map_x_104_s_g_near;
  wire _add_map_x_104_add_exe;
  wire _add_map_x_104_p_reset;
  wire _add_map_x_104_m_clock;
  wire [9:0] _add_map_x_103_moto_org_near;
  wire [9:0] _add_map_x_103_moto_org_near1;
  wire [9:0] _add_map_x_103_moto_org_near2;
  wire [9:0] _add_map_x_103_moto_org_near3;
  wire [9:0] _add_map_x_103_moto_org;
  wire [1:0] _add_map_x_103_sg_up;
  wire [1:0] _add_map_x_103_sg_down;
  wire [1:0] _add_map_x_103_sg_left;
  wire [1:0] _add_map_x_103_sg_right;
  wire _add_map_x_103_wall_t_in;
  wire [9:0] _add_map_x_103_moto;
  wire [9:0] _add_map_x_103_up;
  wire [9:0] _add_map_x_103_right;
  wire [9:0] _add_map_x_103_down;
  wire [9:0] _add_map_x_103_left;
  wire [9:0] _add_map_x_103_start;
  wire [9:0] _add_map_x_103_goal;
  wire [9:0] _add_map_x_103_now;
  wire [9:0] _add_map_x_103_data_out;
  wire [9:0] _add_map_x_103_data_out_index;
  wire [9:0] _add_map_x_103_data_near;
  wire _add_map_x_103_wall_t_out;
  wire [9:0] _add_map_x_103_data_org;
  wire [9:0] _add_map_x_103_data_org_near;
  wire [1:0] _add_map_x_103_s_g;
  wire [1:0] _add_map_x_103_s_g_near;
  wire _add_map_x_103_add_exe;
  wire _add_map_x_103_p_reset;
  wire _add_map_x_103_m_clock;
  wire [9:0] _add_map_x_102_moto_org_near;
  wire [9:0] _add_map_x_102_moto_org_near1;
  wire [9:0] _add_map_x_102_moto_org_near2;
  wire [9:0] _add_map_x_102_moto_org_near3;
  wire [9:0] _add_map_x_102_moto_org;
  wire [1:0] _add_map_x_102_sg_up;
  wire [1:0] _add_map_x_102_sg_down;
  wire [1:0] _add_map_x_102_sg_left;
  wire [1:0] _add_map_x_102_sg_right;
  wire _add_map_x_102_wall_t_in;
  wire [9:0] _add_map_x_102_moto;
  wire [9:0] _add_map_x_102_up;
  wire [9:0] _add_map_x_102_right;
  wire [9:0] _add_map_x_102_down;
  wire [9:0] _add_map_x_102_left;
  wire [9:0] _add_map_x_102_start;
  wire [9:0] _add_map_x_102_goal;
  wire [9:0] _add_map_x_102_now;
  wire [9:0] _add_map_x_102_data_out;
  wire [9:0] _add_map_x_102_data_out_index;
  wire [9:0] _add_map_x_102_data_near;
  wire _add_map_x_102_wall_t_out;
  wire [9:0] _add_map_x_102_data_org;
  wire [9:0] _add_map_x_102_data_org_near;
  wire [1:0] _add_map_x_102_s_g;
  wire [1:0] _add_map_x_102_s_g_near;
  wire _add_map_x_102_add_exe;
  wire _add_map_x_102_p_reset;
  wire _add_map_x_102_m_clock;
  wire [9:0] _add_map_x_101_moto_org_near;
  wire [9:0] _add_map_x_101_moto_org_near1;
  wire [9:0] _add_map_x_101_moto_org_near2;
  wire [9:0] _add_map_x_101_moto_org_near3;
  wire [9:0] _add_map_x_101_moto_org;
  wire [1:0] _add_map_x_101_sg_up;
  wire [1:0] _add_map_x_101_sg_down;
  wire [1:0] _add_map_x_101_sg_left;
  wire [1:0] _add_map_x_101_sg_right;
  wire _add_map_x_101_wall_t_in;
  wire [9:0] _add_map_x_101_moto;
  wire [9:0] _add_map_x_101_up;
  wire [9:0] _add_map_x_101_right;
  wire [9:0] _add_map_x_101_down;
  wire [9:0] _add_map_x_101_left;
  wire [9:0] _add_map_x_101_start;
  wire [9:0] _add_map_x_101_goal;
  wire [9:0] _add_map_x_101_now;
  wire [9:0] _add_map_x_101_data_out;
  wire [9:0] _add_map_x_101_data_out_index;
  wire [9:0] _add_map_x_101_data_near;
  wire _add_map_x_101_wall_t_out;
  wire [9:0] _add_map_x_101_data_org;
  wire [9:0] _add_map_x_101_data_org_near;
  wire [1:0] _add_map_x_101_s_g;
  wire [1:0] _add_map_x_101_s_g_near;
  wire _add_map_x_101_add_exe;
  wire _add_map_x_101_p_reset;
  wire _add_map_x_101_m_clock;
  wire [9:0] _add_map_x_100_moto_org_near;
  wire [9:0] _add_map_x_100_moto_org_near1;
  wire [9:0] _add_map_x_100_moto_org_near2;
  wire [9:0] _add_map_x_100_moto_org_near3;
  wire [9:0] _add_map_x_100_moto_org;
  wire [1:0] _add_map_x_100_sg_up;
  wire [1:0] _add_map_x_100_sg_down;
  wire [1:0] _add_map_x_100_sg_left;
  wire [1:0] _add_map_x_100_sg_right;
  wire _add_map_x_100_wall_t_in;
  wire [9:0] _add_map_x_100_moto;
  wire [9:0] _add_map_x_100_up;
  wire [9:0] _add_map_x_100_right;
  wire [9:0] _add_map_x_100_down;
  wire [9:0] _add_map_x_100_left;
  wire [9:0] _add_map_x_100_start;
  wire [9:0] _add_map_x_100_goal;
  wire [9:0] _add_map_x_100_now;
  wire [9:0] _add_map_x_100_data_out;
  wire [9:0] _add_map_x_100_data_out_index;
  wire [9:0] _add_map_x_100_data_near;
  wire _add_map_x_100_wall_t_out;
  wire [9:0] _add_map_x_100_data_org;
  wire [9:0] _add_map_x_100_data_org_near;
  wire [1:0] _add_map_x_100_s_g;
  wire [1:0] _add_map_x_100_s_g_near;
  wire _add_map_x_100_add_exe;
  wire _add_map_x_100_p_reset;
  wire _add_map_x_100_m_clock;
  wire [9:0] _add_map_x_99_moto_org_near;
  wire [9:0] _add_map_x_99_moto_org_near1;
  wire [9:0] _add_map_x_99_moto_org_near2;
  wire [9:0] _add_map_x_99_moto_org_near3;
  wire [9:0] _add_map_x_99_moto_org;
  wire [1:0] _add_map_x_99_sg_up;
  wire [1:0] _add_map_x_99_sg_down;
  wire [1:0] _add_map_x_99_sg_left;
  wire [1:0] _add_map_x_99_sg_right;
  wire _add_map_x_99_wall_t_in;
  wire [9:0] _add_map_x_99_moto;
  wire [9:0] _add_map_x_99_up;
  wire [9:0] _add_map_x_99_right;
  wire [9:0] _add_map_x_99_down;
  wire [9:0] _add_map_x_99_left;
  wire [9:0] _add_map_x_99_start;
  wire [9:0] _add_map_x_99_goal;
  wire [9:0] _add_map_x_99_now;
  wire [9:0] _add_map_x_99_data_out;
  wire [9:0] _add_map_x_99_data_out_index;
  wire [9:0] _add_map_x_99_data_near;
  wire _add_map_x_99_wall_t_out;
  wire [9:0] _add_map_x_99_data_org;
  wire [9:0] _add_map_x_99_data_org_near;
  wire [1:0] _add_map_x_99_s_g;
  wire [1:0] _add_map_x_99_s_g_near;
  wire _add_map_x_99_add_exe;
  wire _add_map_x_99_p_reset;
  wire _add_map_x_99_m_clock;
  wire [9:0] _add_map_x_98_moto_org_near;
  wire [9:0] _add_map_x_98_moto_org_near1;
  wire [9:0] _add_map_x_98_moto_org_near2;
  wire [9:0] _add_map_x_98_moto_org_near3;
  wire [9:0] _add_map_x_98_moto_org;
  wire [1:0] _add_map_x_98_sg_up;
  wire [1:0] _add_map_x_98_sg_down;
  wire [1:0] _add_map_x_98_sg_left;
  wire [1:0] _add_map_x_98_sg_right;
  wire _add_map_x_98_wall_t_in;
  wire [9:0] _add_map_x_98_moto;
  wire [9:0] _add_map_x_98_up;
  wire [9:0] _add_map_x_98_right;
  wire [9:0] _add_map_x_98_down;
  wire [9:0] _add_map_x_98_left;
  wire [9:0] _add_map_x_98_start;
  wire [9:0] _add_map_x_98_goal;
  wire [9:0] _add_map_x_98_now;
  wire [9:0] _add_map_x_98_data_out;
  wire [9:0] _add_map_x_98_data_out_index;
  wire [9:0] _add_map_x_98_data_near;
  wire _add_map_x_98_wall_t_out;
  wire [9:0] _add_map_x_98_data_org;
  wire [9:0] _add_map_x_98_data_org_near;
  wire [1:0] _add_map_x_98_s_g;
  wire [1:0] _add_map_x_98_s_g_near;
  wire _add_map_x_98_add_exe;
  wire _add_map_x_98_p_reset;
  wire _add_map_x_98_m_clock;
  wire [9:0] _add_map_x_97_moto_org_near;
  wire [9:0] _add_map_x_97_moto_org_near1;
  wire [9:0] _add_map_x_97_moto_org_near2;
  wire [9:0] _add_map_x_97_moto_org_near3;
  wire [9:0] _add_map_x_97_moto_org;
  wire [1:0] _add_map_x_97_sg_up;
  wire [1:0] _add_map_x_97_sg_down;
  wire [1:0] _add_map_x_97_sg_left;
  wire [1:0] _add_map_x_97_sg_right;
  wire _add_map_x_97_wall_t_in;
  wire [9:0] _add_map_x_97_moto;
  wire [9:0] _add_map_x_97_up;
  wire [9:0] _add_map_x_97_right;
  wire [9:0] _add_map_x_97_down;
  wire [9:0] _add_map_x_97_left;
  wire [9:0] _add_map_x_97_start;
  wire [9:0] _add_map_x_97_goal;
  wire [9:0] _add_map_x_97_now;
  wire [9:0] _add_map_x_97_data_out;
  wire [9:0] _add_map_x_97_data_out_index;
  wire [9:0] _add_map_x_97_data_near;
  wire _add_map_x_97_wall_t_out;
  wire [9:0] _add_map_x_97_data_org;
  wire [9:0] _add_map_x_97_data_org_near;
  wire [1:0] _add_map_x_97_s_g;
  wire [1:0] _add_map_x_97_s_g_near;
  wire _add_map_x_97_add_exe;
  wire _add_map_x_97_p_reset;
  wire _add_map_x_97_m_clock;
  wire [9:0] _add_map_x_96_moto_org_near;
  wire [9:0] _add_map_x_96_moto_org_near1;
  wire [9:0] _add_map_x_96_moto_org_near2;
  wire [9:0] _add_map_x_96_moto_org_near3;
  wire [9:0] _add_map_x_96_moto_org;
  wire [1:0] _add_map_x_96_sg_up;
  wire [1:0] _add_map_x_96_sg_down;
  wire [1:0] _add_map_x_96_sg_left;
  wire [1:0] _add_map_x_96_sg_right;
  wire _add_map_x_96_wall_t_in;
  wire [9:0] _add_map_x_96_moto;
  wire [9:0] _add_map_x_96_up;
  wire [9:0] _add_map_x_96_right;
  wire [9:0] _add_map_x_96_down;
  wire [9:0] _add_map_x_96_left;
  wire [9:0] _add_map_x_96_start;
  wire [9:0] _add_map_x_96_goal;
  wire [9:0] _add_map_x_96_now;
  wire [9:0] _add_map_x_96_data_out;
  wire [9:0] _add_map_x_96_data_out_index;
  wire [9:0] _add_map_x_96_data_near;
  wire _add_map_x_96_wall_t_out;
  wire [9:0] _add_map_x_96_data_org;
  wire [9:0] _add_map_x_96_data_org_near;
  wire [1:0] _add_map_x_96_s_g;
  wire [1:0] _add_map_x_96_s_g_near;
  wire _add_map_x_96_add_exe;
  wire _add_map_x_96_p_reset;
  wire _add_map_x_96_m_clock;
  wire [9:0] _add_map_x_95_moto_org_near;
  wire [9:0] _add_map_x_95_moto_org_near1;
  wire [9:0] _add_map_x_95_moto_org_near2;
  wire [9:0] _add_map_x_95_moto_org_near3;
  wire [9:0] _add_map_x_95_moto_org;
  wire [1:0] _add_map_x_95_sg_up;
  wire [1:0] _add_map_x_95_sg_down;
  wire [1:0] _add_map_x_95_sg_left;
  wire [1:0] _add_map_x_95_sg_right;
  wire _add_map_x_95_wall_t_in;
  wire [9:0] _add_map_x_95_moto;
  wire [9:0] _add_map_x_95_up;
  wire [9:0] _add_map_x_95_right;
  wire [9:0] _add_map_x_95_down;
  wire [9:0] _add_map_x_95_left;
  wire [9:0] _add_map_x_95_start;
  wire [9:0] _add_map_x_95_goal;
  wire [9:0] _add_map_x_95_now;
  wire [9:0] _add_map_x_95_data_out;
  wire [9:0] _add_map_x_95_data_out_index;
  wire [9:0] _add_map_x_95_data_near;
  wire _add_map_x_95_wall_t_out;
  wire [9:0] _add_map_x_95_data_org;
  wire [9:0] _add_map_x_95_data_org_near;
  wire [1:0] _add_map_x_95_s_g;
  wire [1:0] _add_map_x_95_s_g_near;
  wire _add_map_x_95_add_exe;
  wire _add_map_x_95_p_reset;
  wire _add_map_x_95_m_clock;
  wire [9:0] _add_map_x_94_moto_org_near;
  wire [9:0] _add_map_x_94_moto_org_near1;
  wire [9:0] _add_map_x_94_moto_org_near2;
  wire [9:0] _add_map_x_94_moto_org_near3;
  wire [9:0] _add_map_x_94_moto_org;
  wire [1:0] _add_map_x_94_sg_up;
  wire [1:0] _add_map_x_94_sg_down;
  wire [1:0] _add_map_x_94_sg_left;
  wire [1:0] _add_map_x_94_sg_right;
  wire _add_map_x_94_wall_t_in;
  wire [9:0] _add_map_x_94_moto;
  wire [9:0] _add_map_x_94_up;
  wire [9:0] _add_map_x_94_right;
  wire [9:0] _add_map_x_94_down;
  wire [9:0] _add_map_x_94_left;
  wire [9:0] _add_map_x_94_start;
  wire [9:0] _add_map_x_94_goal;
  wire [9:0] _add_map_x_94_now;
  wire [9:0] _add_map_x_94_data_out;
  wire [9:0] _add_map_x_94_data_out_index;
  wire [9:0] _add_map_x_94_data_near;
  wire _add_map_x_94_wall_t_out;
  wire [9:0] _add_map_x_94_data_org;
  wire [9:0] _add_map_x_94_data_org_near;
  wire [1:0] _add_map_x_94_s_g;
  wire [1:0] _add_map_x_94_s_g_near;
  wire _add_map_x_94_add_exe;
  wire _add_map_x_94_p_reset;
  wire _add_map_x_94_m_clock;
  wire [9:0] _add_map_x_93_moto_org_near;
  wire [9:0] _add_map_x_93_moto_org_near1;
  wire [9:0] _add_map_x_93_moto_org_near2;
  wire [9:0] _add_map_x_93_moto_org_near3;
  wire [9:0] _add_map_x_93_moto_org;
  wire [1:0] _add_map_x_93_sg_up;
  wire [1:0] _add_map_x_93_sg_down;
  wire [1:0] _add_map_x_93_sg_left;
  wire [1:0] _add_map_x_93_sg_right;
  wire _add_map_x_93_wall_t_in;
  wire [9:0] _add_map_x_93_moto;
  wire [9:0] _add_map_x_93_up;
  wire [9:0] _add_map_x_93_right;
  wire [9:0] _add_map_x_93_down;
  wire [9:0] _add_map_x_93_left;
  wire [9:0] _add_map_x_93_start;
  wire [9:0] _add_map_x_93_goal;
  wire [9:0] _add_map_x_93_now;
  wire [9:0] _add_map_x_93_data_out;
  wire [9:0] _add_map_x_93_data_out_index;
  wire [9:0] _add_map_x_93_data_near;
  wire _add_map_x_93_wall_t_out;
  wire [9:0] _add_map_x_93_data_org;
  wire [9:0] _add_map_x_93_data_org_near;
  wire [1:0] _add_map_x_93_s_g;
  wire [1:0] _add_map_x_93_s_g_near;
  wire _add_map_x_93_add_exe;
  wire _add_map_x_93_p_reset;
  wire _add_map_x_93_m_clock;
  wire [9:0] _add_map_x_92_moto_org_near;
  wire [9:0] _add_map_x_92_moto_org_near1;
  wire [9:0] _add_map_x_92_moto_org_near2;
  wire [9:0] _add_map_x_92_moto_org_near3;
  wire [9:0] _add_map_x_92_moto_org;
  wire [1:0] _add_map_x_92_sg_up;
  wire [1:0] _add_map_x_92_sg_down;
  wire [1:0] _add_map_x_92_sg_left;
  wire [1:0] _add_map_x_92_sg_right;
  wire _add_map_x_92_wall_t_in;
  wire [9:0] _add_map_x_92_moto;
  wire [9:0] _add_map_x_92_up;
  wire [9:0] _add_map_x_92_right;
  wire [9:0] _add_map_x_92_down;
  wire [9:0] _add_map_x_92_left;
  wire [9:0] _add_map_x_92_start;
  wire [9:0] _add_map_x_92_goal;
  wire [9:0] _add_map_x_92_now;
  wire [9:0] _add_map_x_92_data_out;
  wire [9:0] _add_map_x_92_data_out_index;
  wire [9:0] _add_map_x_92_data_near;
  wire _add_map_x_92_wall_t_out;
  wire [9:0] _add_map_x_92_data_org;
  wire [9:0] _add_map_x_92_data_org_near;
  wire [1:0] _add_map_x_92_s_g;
  wire [1:0] _add_map_x_92_s_g_near;
  wire _add_map_x_92_add_exe;
  wire _add_map_x_92_p_reset;
  wire _add_map_x_92_m_clock;
  wire [9:0] _add_map_x_91_moto_org_near;
  wire [9:0] _add_map_x_91_moto_org_near1;
  wire [9:0] _add_map_x_91_moto_org_near2;
  wire [9:0] _add_map_x_91_moto_org_near3;
  wire [9:0] _add_map_x_91_moto_org;
  wire [1:0] _add_map_x_91_sg_up;
  wire [1:0] _add_map_x_91_sg_down;
  wire [1:0] _add_map_x_91_sg_left;
  wire [1:0] _add_map_x_91_sg_right;
  wire _add_map_x_91_wall_t_in;
  wire [9:0] _add_map_x_91_moto;
  wire [9:0] _add_map_x_91_up;
  wire [9:0] _add_map_x_91_right;
  wire [9:0] _add_map_x_91_down;
  wire [9:0] _add_map_x_91_left;
  wire [9:0] _add_map_x_91_start;
  wire [9:0] _add_map_x_91_goal;
  wire [9:0] _add_map_x_91_now;
  wire [9:0] _add_map_x_91_data_out;
  wire [9:0] _add_map_x_91_data_out_index;
  wire [9:0] _add_map_x_91_data_near;
  wire _add_map_x_91_wall_t_out;
  wire [9:0] _add_map_x_91_data_org;
  wire [9:0] _add_map_x_91_data_org_near;
  wire [1:0] _add_map_x_91_s_g;
  wire [1:0] _add_map_x_91_s_g_near;
  wire _add_map_x_91_add_exe;
  wire _add_map_x_91_p_reset;
  wire _add_map_x_91_m_clock;
  wire [9:0] _add_map_x_90_moto_org_near;
  wire [9:0] _add_map_x_90_moto_org_near1;
  wire [9:0] _add_map_x_90_moto_org_near2;
  wire [9:0] _add_map_x_90_moto_org_near3;
  wire [9:0] _add_map_x_90_moto_org;
  wire [1:0] _add_map_x_90_sg_up;
  wire [1:0] _add_map_x_90_sg_down;
  wire [1:0] _add_map_x_90_sg_left;
  wire [1:0] _add_map_x_90_sg_right;
  wire _add_map_x_90_wall_t_in;
  wire [9:0] _add_map_x_90_moto;
  wire [9:0] _add_map_x_90_up;
  wire [9:0] _add_map_x_90_right;
  wire [9:0] _add_map_x_90_down;
  wire [9:0] _add_map_x_90_left;
  wire [9:0] _add_map_x_90_start;
  wire [9:0] _add_map_x_90_goal;
  wire [9:0] _add_map_x_90_now;
  wire [9:0] _add_map_x_90_data_out;
  wire [9:0] _add_map_x_90_data_out_index;
  wire [9:0] _add_map_x_90_data_near;
  wire _add_map_x_90_wall_t_out;
  wire [9:0] _add_map_x_90_data_org;
  wire [9:0] _add_map_x_90_data_org_near;
  wire [1:0] _add_map_x_90_s_g;
  wire [1:0] _add_map_x_90_s_g_near;
  wire _add_map_x_90_add_exe;
  wire _add_map_x_90_p_reset;
  wire _add_map_x_90_m_clock;
  wire [9:0] _add_map_x_89_moto_org_near;
  wire [9:0] _add_map_x_89_moto_org_near1;
  wire [9:0] _add_map_x_89_moto_org_near2;
  wire [9:0] _add_map_x_89_moto_org_near3;
  wire [9:0] _add_map_x_89_moto_org;
  wire [1:0] _add_map_x_89_sg_up;
  wire [1:0] _add_map_x_89_sg_down;
  wire [1:0] _add_map_x_89_sg_left;
  wire [1:0] _add_map_x_89_sg_right;
  wire _add_map_x_89_wall_t_in;
  wire [9:0] _add_map_x_89_moto;
  wire [9:0] _add_map_x_89_up;
  wire [9:0] _add_map_x_89_right;
  wire [9:0] _add_map_x_89_down;
  wire [9:0] _add_map_x_89_left;
  wire [9:0] _add_map_x_89_start;
  wire [9:0] _add_map_x_89_goal;
  wire [9:0] _add_map_x_89_now;
  wire [9:0] _add_map_x_89_data_out;
  wire [9:0] _add_map_x_89_data_out_index;
  wire [9:0] _add_map_x_89_data_near;
  wire _add_map_x_89_wall_t_out;
  wire [9:0] _add_map_x_89_data_org;
  wire [9:0] _add_map_x_89_data_org_near;
  wire [1:0] _add_map_x_89_s_g;
  wire [1:0] _add_map_x_89_s_g_near;
  wire _add_map_x_89_add_exe;
  wire _add_map_x_89_p_reset;
  wire _add_map_x_89_m_clock;
  wire [9:0] _add_map_x_88_moto_org_near;
  wire [9:0] _add_map_x_88_moto_org_near1;
  wire [9:0] _add_map_x_88_moto_org_near2;
  wire [9:0] _add_map_x_88_moto_org_near3;
  wire [9:0] _add_map_x_88_moto_org;
  wire [1:0] _add_map_x_88_sg_up;
  wire [1:0] _add_map_x_88_sg_down;
  wire [1:0] _add_map_x_88_sg_left;
  wire [1:0] _add_map_x_88_sg_right;
  wire _add_map_x_88_wall_t_in;
  wire [9:0] _add_map_x_88_moto;
  wire [9:0] _add_map_x_88_up;
  wire [9:0] _add_map_x_88_right;
  wire [9:0] _add_map_x_88_down;
  wire [9:0] _add_map_x_88_left;
  wire [9:0] _add_map_x_88_start;
  wire [9:0] _add_map_x_88_goal;
  wire [9:0] _add_map_x_88_now;
  wire [9:0] _add_map_x_88_data_out;
  wire [9:0] _add_map_x_88_data_out_index;
  wire [9:0] _add_map_x_88_data_near;
  wire _add_map_x_88_wall_t_out;
  wire [9:0] _add_map_x_88_data_org;
  wire [9:0] _add_map_x_88_data_org_near;
  wire [1:0] _add_map_x_88_s_g;
  wire [1:0] _add_map_x_88_s_g_near;
  wire _add_map_x_88_add_exe;
  wire _add_map_x_88_p_reset;
  wire _add_map_x_88_m_clock;
  wire [9:0] _add_map_x_87_moto_org_near;
  wire [9:0] _add_map_x_87_moto_org_near1;
  wire [9:0] _add_map_x_87_moto_org_near2;
  wire [9:0] _add_map_x_87_moto_org_near3;
  wire [9:0] _add_map_x_87_moto_org;
  wire [1:0] _add_map_x_87_sg_up;
  wire [1:0] _add_map_x_87_sg_down;
  wire [1:0] _add_map_x_87_sg_left;
  wire [1:0] _add_map_x_87_sg_right;
  wire _add_map_x_87_wall_t_in;
  wire [9:0] _add_map_x_87_moto;
  wire [9:0] _add_map_x_87_up;
  wire [9:0] _add_map_x_87_right;
  wire [9:0] _add_map_x_87_down;
  wire [9:0] _add_map_x_87_left;
  wire [9:0] _add_map_x_87_start;
  wire [9:0] _add_map_x_87_goal;
  wire [9:0] _add_map_x_87_now;
  wire [9:0] _add_map_x_87_data_out;
  wire [9:0] _add_map_x_87_data_out_index;
  wire [9:0] _add_map_x_87_data_near;
  wire _add_map_x_87_wall_t_out;
  wire [9:0] _add_map_x_87_data_org;
  wire [9:0] _add_map_x_87_data_org_near;
  wire [1:0] _add_map_x_87_s_g;
  wire [1:0] _add_map_x_87_s_g_near;
  wire _add_map_x_87_add_exe;
  wire _add_map_x_87_p_reset;
  wire _add_map_x_87_m_clock;
  wire [9:0] _add_map_x_86_moto_org_near;
  wire [9:0] _add_map_x_86_moto_org_near1;
  wire [9:0] _add_map_x_86_moto_org_near2;
  wire [9:0] _add_map_x_86_moto_org_near3;
  wire [9:0] _add_map_x_86_moto_org;
  wire [1:0] _add_map_x_86_sg_up;
  wire [1:0] _add_map_x_86_sg_down;
  wire [1:0] _add_map_x_86_sg_left;
  wire [1:0] _add_map_x_86_sg_right;
  wire _add_map_x_86_wall_t_in;
  wire [9:0] _add_map_x_86_moto;
  wire [9:0] _add_map_x_86_up;
  wire [9:0] _add_map_x_86_right;
  wire [9:0] _add_map_x_86_down;
  wire [9:0] _add_map_x_86_left;
  wire [9:0] _add_map_x_86_start;
  wire [9:0] _add_map_x_86_goal;
  wire [9:0] _add_map_x_86_now;
  wire [9:0] _add_map_x_86_data_out;
  wire [9:0] _add_map_x_86_data_out_index;
  wire [9:0] _add_map_x_86_data_near;
  wire _add_map_x_86_wall_t_out;
  wire [9:0] _add_map_x_86_data_org;
  wire [9:0] _add_map_x_86_data_org_near;
  wire [1:0] _add_map_x_86_s_g;
  wire [1:0] _add_map_x_86_s_g_near;
  wire _add_map_x_86_add_exe;
  wire _add_map_x_86_p_reset;
  wire _add_map_x_86_m_clock;
  wire [9:0] _add_map_x_85_moto_org_near;
  wire [9:0] _add_map_x_85_moto_org_near1;
  wire [9:0] _add_map_x_85_moto_org_near2;
  wire [9:0] _add_map_x_85_moto_org_near3;
  wire [9:0] _add_map_x_85_moto_org;
  wire [1:0] _add_map_x_85_sg_up;
  wire [1:0] _add_map_x_85_sg_down;
  wire [1:0] _add_map_x_85_sg_left;
  wire [1:0] _add_map_x_85_sg_right;
  wire _add_map_x_85_wall_t_in;
  wire [9:0] _add_map_x_85_moto;
  wire [9:0] _add_map_x_85_up;
  wire [9:0] _add_map_x_85_right;
  wire [9:0] _add_map_x_85_down;
  wire [9:0] _add_map_x_85_left;
  wire [9:0] _add_map_x_85_start;
  wire [9:0] _add_map_x_85_goal;
  wire [9:0] _add_map_x_85_now;
  wire [9:0] _add_map_x_85_data_out;
  wire [9:0] _add_map_x_85_data_out_index;
  wire [9:0] _add_map_x_85_data_near;
  wire _add_map_x_85_wall_t_out;
  wire [9:0] _add_map_x_85_data_org;
  wire [9:0] _add_map_x_85_data_org_near;
  wire [1:0] _add_map_x_85_s_g;
  wire [1:0] _add_map_x_85_s_g_near;
  wire _add_map_x_85_add_exe;
  wire _add_map_x_85_p_reset;
  wire _add_map_x_85_m_clock;
  wire [9:0] _add_map_x_84_moto_org_near;
  wire [9:0] _add_map_x_84_moto_org_near1;
  wire [9:0] _add_map_x_84_moto_org_near2;
  wire [9:0] _add_map_x_84_moto_org_near3;
  wire [9:0] _add_map_x_84_moto_org;
  wire [1:0] _add_map_x_84_sg_up;
  wire [1:0] _add_map_x_84_sg_down;
  wire [1:0] _add_map_x_84_sg_left;
  wire [1:0] _add_map_x_84_sg_right;
  wire _add_map_x_84_wall_t_in;
  wire [9:0] _add_map_x_84_moto;
  wire [9:0] _add_map_x_84_up;
  wire [9:0] _add_map_x_84_right;
  wire [9:0] _add_map_x_84_down;
  wire [9:0] _add_map_x_84_left;
  wire [9:0] _add_map_x_84_start;
  wire [9:0] _add_map_x_84_goal;
  wire [9:0] _add_map_x_84_now;
  wire [9:0] _add_map_x_84_data_out;
  wire [9:0] _add_map_x_84_data_out_index;
  wire [9:0] _add_map_x_84_data_near;
  wire _add_map_x_84_wall_t_out;
  wire [9:0] _add_map_x_84_data_org;
  wire [9:0] _add_map_x_84_data_org_near;
  wire [1:0] _add_map_x_84_s_g;
  wire [1:0] _add_map_x_84_s_g_near;
  wire _add_map_x_84_add_exe;
  wire _add_map_x_84_p_reset;
  wire _add_map_x_84_m_clock;
  wire [9:0] _add_map_x_83_moto_org_near;
  wire [9:0] _add_map_x_83_moto_org_near1;
  wire [9:0] _add_map_x_83_moto_org_near2;
  wire [9:0] _add_map_x_83_moto_org_near3;
  wire [9:0] _add_map_x_83_moto_org;
  wire [1:0] _add_map_x_83_sg_up;
  wire [1:0] _add_map_x_83_sg_down;
  wire [1:0] _add_map_x_83_sg_left;
  wire [1:0] _add_map_x_83_sg_right;
  wire _add_map_x_83_wall_t_in;
  wire [9:0] _add_map_x_83_moto;
  wire [9:0] _add_map_x_83_up;
  wire [9:0] _add_map_x_83_right;
  wire [9:0] _add_map_x_83_down;
  wire [9:0] _add_map_x_83_left;
  wire [9:0] _add_map_x_83_start;
  wire [9:0] _add_map_x_83_goal;
  wire [9:0] _add_map_x_83_now;
  wire [9:0] _add_map_x_83_data_out;
  wire [9:0] _add_map_x_83_data_out_index;
  wire [9:0] _add_map_x_83_data_near;
  wire _add_map_x_83_wall_t_out;
  wire [9:0] _add_map_x_83_data_org;
  wire [9:0] _add_map_x_83_data_org_near;
  wire [1:0] _add_map_x_83_s_g;
  wire [1:0] _add_map_x_83_s_g_near;
  wire _add_map_x_83_add_exe;
  wire _add_map_x_83_p_reset;
  wire _add_map_x_83_m_clock;
  wire [9:0] _add_map_x_82_moto_org_near;
  wire [9:0] _add_map_x_82_moto_org_near1;
  wire [9:0] _add_map_x_82_moto_org_near2;
  wire [9:0] _add_map_x_82_moto_org_near3;
  wire [9:0] _add_map_x_82_moto_org;
  wire [1:0] _add_map_x_82_sg_up;
  wire [1:0] _add_map_x_82_sg_down;
  wire [1:0] _add_map_x_82_sg_left;
  wire [1:0] _add_map_x_82_sg_right;
  wire _add_map_x_82_wall_t_in;
  wire [9:0] _add_map_x_82_moto;
  wire [9:0] _add_map_x_82_up;
  wire [9:0] _add_map_x_82_right;
  wire [9:0] _add_map_x_82_down;
  wire [9:0] _add_map_x_82_left;
  wire [9:0] _add_map_x_82_start;
  wire [9:0] _add_map_x_82_goal;
  wire [9:0] _add_map_x_82_now;
  wire [9:0] _add_map_x_82_data_out;
  wire [9:0] _add_map_x_82_data_out_index;
  wire [9:0] _add_map_x_82_data_near;
  wire _add_map_x_82_wall_t_out;
  wire [9:0] _add_map_x_82_data_org;
  wire [9:0] _add_map_x_82_data_org_near;
  wire [1:0] _add_map_x_82_s_g;
  wire [1:0] _add_map_x_82_s_g_near;
  wire _add_map_x_82_add_exe;
  wire _add_map_x_82_p_reset;
  wire _add_map_x_82_m_clock;
  wire [9:0] _add_map_x_81_moto_org_near;
  wire [9:0] _add_map_x_81_moto_org_near1;
  wire [9:0] _add_map_x_81_moto_org_near2;
  wire [9:0] _add_map_x_81_moto_org_near3;
  wire [9:0] _add_map_x_81_moto_org;
  wire [1:0] _add_map_x_81_sg_up;
  wire [1:0] _add_map_x_81_sg_down;
  wire [1:0] _add_map_x_81_sg_left;
  wire [1:0] _add_map_x_81_sg_right;
  wire _add_map_x_81_wall_t_in;
  wire [9:0] _add_map_x_81_moto;
  wire [9:0] _add_map_x_81_up;
  wire [9:0] _add_map_x_81_right;
  wire [9:0] _add_map_x_81_down;
  wire [9:0] _add_map_x_81_left;
  wire [9:0] _add_map_x_81_start;
  wire [9:0] _add_map_x_81_goal;
  wire [9:0] _add_map_x_81_now;
  wire [9:0] _add_map_x_81_data_out;
  wire [9:0] _add_map_x_81_data_out_index;
  wire [9:0] _add_map_x_81_data_near;
  wire _add_map_x_81_wall_t_out;
  wire [9:0] _add_map_x_81_data_org;
  wire [9:0] _add_map_x_81_data_org_near;
  wire [1:0] _add_map_x_81_s_g;
  wire [1:0] _add_map_x_81_s_g_near;
  wire _add_map_x_81_add_exe;
  wire _add_map_x_81_p_reset;
  wire _add_map_x_81_m_clock;
  wire [9:0] _add_map_x_80_moto_org_near;
  wire [9:0] _add_map_x_80_moto_org_near1;
  wire [9:0] _add_map_x_80_moto_org_near2;
  wire [9:0] _add_map_x_80_moto_org_near3;
  wire [9:0] _add_map_x_80_moto_org;
  wire [1:0] _add_map_x_80_sg_up;
  wire [1:0] _add_map_x_80_sg_down;
  wire [1:0] _add_map_x_80_sg_left;
  wire [1:0] _add_map_x_80_sg_right;
  wire _add_map_x_80_wall_t_in;
  wire [9:0] _add_map_x_80_moto;
  wire [9:0] _add_map_x_80_up;
  wire [9:0] _add_map_x_80_right;
  wire [9:0] _add_map_x_80_down;
  wire [9:0] _add_map_x_80_left;
  wire [9:0] _add_map_x_80_start;
  wire [9:0] _add_map_x_80_goal;
  wire [9:0] _add_map_x_80_now;
  wire [9:0] _add_map_x_80_data_out;
  wire [9:0] _add_map_x_80_data_out_index;
  wire [9:0] _add_map_x_80_data_near;
  wire _add_map_x_80_wall_t_out;
  wire [9:0] _add_map_x_80_data_org;
  wire [9:0] _add_map_x_80_data_org_near;
  wire [1:0] _add_map_x_80_s_g;
  wire [1:0] _add_map_x_80_s_g_near;
  wire _add_map_x_80_add_exe;
  wire _add_map_x_80_p_reset;
  wire _add_map_x_80_m_clock;
  wire [9:0] _add_map_x_79_moto_org_near;
  wire [9:0] _add_map_x_79_moto_org_near1;
  wire [9:0] _add_map_x_79_moto_org_near2;
  wire [9:0] _add_map_x_79_moto_org_near3;
  wire [9:0] _add_map_x_79_moto_org;
  wire [1:0] _add_map_x_79_sg_up;
  wire [1:0] _add_map_x_79_sg_down;
  wire [1:0] _add_map_x_79_sg_left;
  wire [1:0] _add_map_x_79_sg_right;
  wire _add_map_x_79_wall_t_in;
  wire [9:0] _add_map_x_79_moto;
  wire [9:0] _add_map_x_79_up;
  wire [9:0] _add_map_x_79_right;
  wire [9:0] _add_map_x_79_down;
  wire [9:0] _add_map_x_79_left;
  wire [9:0] _add_map_x_79_start;
  wire [9:0] _add_map_x_79_goal;
  wire [9:0] _add_map_x_79_now;
  wire [9:0] _add_map_x_79_data_out;
  wire [9:0] _add_map_x_79_data_out_index;
  wire [9:0] _add_map_x_79_data_near;
  wire _add_map_x_79_wall_t_out;
  wire [9:0] _add_map_x_79_data_org;
  wire [9:0] _add_map_x_79_data_org_near;
  wire [1:0] _add_map_x_79_s_g;
  wire [1:0] _add_map_x_79_s_g_near;
  wire _add_map_x_79_add_exe;
  wire _add_map_x_79_p_reset;
  wire _add_map_x_79_m_clock;
  wire [9:0] _add_map_x_78_moto_org_near;
  wire [9:0] _add_map_x_78_moto_org_near1;
  wire [9:0] _add_map_x_78_moto_org_near2;
  wire [9:0] _add_map_x_78_moto_org_near3;
  wire [9:0] _add_map_x_78_moto_org;
  wire [1:0] _add_map_x_78_sg_up;
  wire [1:0] _add_map_x_78_sg_down;
  wire [1:0] _add_map_x_78_sg_left;
  wire [1:0] _add_map_x_78_sg_right;
  wire _add_map_x_78_wall_t_in;
  wire [9:0] _add_map_x_78_moto;
  wire [9:0] _add_map_x_78_up;
  wire [9:0] _add_map_x_78_right;
  wire [9:0] _add_map_x_78_down;
  wire [9:0] _add_map_x_78_left;
  wire [9:0] _add_map_x_78_start;
  wire [9:0] _add_map_x_78_goal;
  wire [9:0] _add_map_x_78_now;
  wire [9:0] _add_map_x_78_data_out;
  wire [9:0] _add_map_x_78_data_out_index;
  wire [9:0] _add_map_x_78_data_near;
  wire _add_map_x_78_wall_t_out;
  wire [9:0] _add_map_x_78_data_org;
  wire [9:0] _add_map_x_78_data_org_near;
  wire [1:0] _add_map_x_78_s_g;
  wire [1:0] _add_map_x_78_s_g_near;
  wire _add_map_x_78_add_exe;
  wire _add_map_x_78_p_reset;
  wire _add_map_x_78_m_clock;
  wire [9:0] _add_map_x_77_moto_org_near;
  wire [9:0] _add_map_x_77_moto_org_near1;
  wire [9:0] _add_map_x_77_moto_org_near2;
  wire [9:0] _add_map_x_77_moto_org_near3;
  wire [9:0] _add_map_x_77_moto_org;
  wire [1:0] _add_map_x_77_sg_up;
  wire [1:0] _add_map_x_77_sg_down;
  wire [1:0] _add_map_x_77_sg_left;
  wire [1:0] _add_map_x_77_sg_right;
  wire _add_map_x_77_wall_t_in;
  wire [9:0] _add_map_x_77_moto;
  wire [9:0] _add_map_x_77_up;
  wire [9:0] _add_map_x_77_right;
  wire [9:0] _add_map_x_77_down;
  wire [9:0] _add_map_x_77_left;
  wire [9:0] _add_map_x_77_start;
  wire [9:0] _add_map_x_77_goal;
  wire [9:0] _add_map_x_77_now;
  wire [9:0] _add_map_x_77_data_out;
  wire [9:0] _add_map_x_77_data_out_index;
  wire [9:0] _add_map_x_77_data_near;
  wire _add_map_x_77_wall_t_out;
  wire [9:0] _add_map_x_77_data_org;
  wire [9:0] _add_map_x_77_data_org_near;
  wire [1:0] _add_map_x_77_s_g;
  wire [1:0] _add_map_x_77_s_g_near;
  wire _add_map_x_77_add_exe;
  wire _add_map_x_77_p_reset;
  wire _add_map_x_77_m_clock;
  wire [9:0] _add_map_x_76_moto_org_near;
  wire [9:0] _add_map_x_76_moto_org_near1;
  wire [9:0] _add_map_x_76_moto_org_near2;
  wire [9:0] _add_map_x_76_moto_org_near3;
  wire [9:0] _add_map_x_76_moto_org;
  wire [1:0] _add_map_x_76_sg_up;
  wire [1:0] _add_map_x_76_sg_down;
  wire [1:0] _add_map_x_76_sg_left;
  wire [1:0] _add_map_x_76_sg_right;
  wire _add_map_x_76_wall_t_in;
  wire [9:0] _add_map_x_76_moto;
  wire [9:0] _add_map_x_76_up;
  wire [9:0] _add_map_x_76_right;
  wire [9:0] _add_map_x_76_down;
  wire [9:0] _add_map_x_76_left;
  wire [9:0] _add_map_x_76_start;
  wire [9:0] _add_map_x_76_goal;
  wire [9:0] _add_map_x_76_now;
  wire [9:0] _add_map_x_76_data_out;
  wire [9:0] _add_map_x_76_data_out_index;
  wire [9:0] _add_map_x_76_data_near;
  wire _add_map_x_76_wall_t_out;
  wire [9:0] _add_map_x_76_data_org;
  wire [9:0] _add_map_x_76_data_org_near;
  wire [1:0] _add_map_x_76_s_g;
  wire [1:0] _add_map_x_76_s_g_near;
  wire _add_map_x_76_add_exe;
  wire _add_map_x_76_p_reset;
  wire _add_map_x_76_m_clock;
  wire [9:0] _add_map_x_75_moto_org_near;
  wire [9:0] _add_map_x_75_moto_org_near1;
  wire [9:0] _add_map_x_75_moto_org_near2;
  wire [9:0] _add_map_x_75_moto_org_near3;
  wire [9:0] _add_map_x_75_moto_org;
  wire [1:0] _add_map_x_75_sg_up;
  wire [1:0] _add_map_x_75_sg_down;
  wire [1:0] _add_map_x_75_sg_left;
  wire [1:0] _add_map_x_75_sg_right;
  wire _add_map_x_75_wall_t_in;
  wire [9:0] _add_map_x_75_moto;
  wire [9:0] _add_map_x_75_up;
  wire [9:0] _add_map_x_75_right;
  wire [9:0] _add_map_x_75_down;
  wire [9:0] _add_map_x_75_left;
  wire [9:0] _add_map_x_75_start;
  wire [9:0] _add_map_x_75_goal;
  wire [9:0] _add_map_x_75_now;
  wire [9:0] _add_map_x_75_data_out;
  wire [9:0] _add_map_x_75_data_out_index;
  wire [9:0] _add_map_x_75_data_near;
  wire _add_map_x_75_wall_t_out;
  wire [9:0] _add_map_x_75_data_org;
  wire [9:0] _add_map_x_75_data_org_near;
  wire [1:0] _add_map_x_75_s_g;
  wire [1:0] _add_map_x_75_s_g_near;
  wire _add_map_x_75_add_exe;
  wire _add_map_x_75_p_reset;
  wire _add_map_x_75_m_clock;
  wire [9:0] _add_map_x_74_moto_org_near;
  wire [9:0] _add_map_x_74_moto_org_near1;
  wire [9:0] _add_map_x_74_moto_org_near2;
  wire [9:0] _add_map_x_74_moto_org_near3;
  wire [9:0] _add_map_x_74_moto_org;
  wire [1:0] _add_map_x_74_sg_up;
  wire [1:0] _add_map_x_74_sg_down;
  wire [1:0] _add_map_x_74_sg_left;
  wire [1:0] _add_map_x_74_sg_right;
  wire _add_map_x_74_wall_t_in;
  wire [9:0] _add_map_x_74_moto;
  wire [9:0] _add_map_x_74_up;
  wire [9:0] _add_map_x_74_right;
  wire [9:0] _add_map_x_74_down;
  wire [9:0] _add_map_x_74_left;
  wire [9:0] _add_map_x_74_start;
  wire [9:0] _add_map_x_74_goal;
  wire [9:0] _add_map_x_74_now;
  wire [9:0] _add_map_x_74_data_out;
  wire [9:0] _add_map_x_74_data_out_index;
  wire [9:0] _add_map_x_74_data_near;
  wire _add_map_x_74_wall_t_out;
  wire [9:0] _add_map_x_74_data_org;
  wire [9:0] _add_map_x_74_data_org_near;
  wire [1:0] _add_map_x_74_s_g;
  wire [1:0] _add_map_x_74_s_g_near;
  wire _add_map_x_74_add_exe;
  wire _add_map_x_74_p_reset;
  wire _add_map_x_74_m_clock;
  wire [9:0] _add_map_x_73_moto_org_near;
  wire [9:0] _add_map_x_73_moto_org_near1;
  wire [9:0] _add_map_x_73_moto_org_near2;
  wire [9:0] _add_map_x_73_moto_org_near3;
  wire [9:0] _add_map_x_73_moto_org;
  wire [1:0] _add_map_x_73_sg_up;
  wire [1:0] _add_map_x_73_sg_down;
  wire [1:0] _add_map_x_73_sg_left;
  wire [1:0] _add_map_x_73_sg_right;
  wire _add_map_x_73_wall_t_in;
  wire [9:0] _add_map_x_73_moto;
  wire [9:0] _add_map_x_73_up;
  wire [9:0] _add_map_x_73_right;
  wire [9:0] _add_map_x_73_down;
  wire [9:0] _add_map_x_73_left;
  wire [9:0] _add_map_x_73_start;
  wire [9:0] _add_map_x_73_goal;
  wire [9:0] _add_map_x_73_now;
  wire [9:0] _add_map_x_73_data_out;
  wire [9:0] _add_map_x_73_data_out_index;
  wire [9:0] _add_map_x_73_data_near;
  wire _add_map_x_73_wall_t_out;
  wire [9:0] _add_map_x_73_data_org;
  wire [9:0] _add_map_x_73_data_org_near;
  wire [1:0] _add_map_x_73_s_g;
  wire [1:0] _add_map_x_73_s_g_near;
  wire _add_map_x_73_add_exe;
  wire _add_map_x_73_p_reset;
  wire _add_map_x_73_m_clock;
  wire [9:0] _add_map_x_72_moto_org_near;
  wire [9:0] _add_map_x_72_moto_org_near1;
  wire [9:0] _add_map_x_72_moto_org_near2;
  wire [9:0] _add_map_x_72_moto_org_near3;
  wire [9:0] _add_map_x_72_moto_org;
  wire [1:0] _add_map_x_72_sg_up;
  wire [1:0] _add_map_x_72_sg_down;
  wire [1:0] _add_map_x_72_sg_left;
  wire [1:0] _add_map_x_72_sg_right;
  wire _add_map_x_72_wall_t_in;
  wire [9:0] _add_map_x_72_moto;
  wire [9:0] _add_map_x_72_up;
  wire [9:0] _add_map_x_72_right;
  wire [9:0] _add_map_x_72_down;
  wire [9:0] _add_map_x_72_left;
  wire [9:0] _add_map_x_72_start;
  wire [9:0] _add_map_x_72_goal;
  wire [9:0] _add_map_x_72_now;
  wire [9:0] _add_map_x_72_data_out;
  wire [9:0] _add_map_x_72_data_out_index;
  wire [9:0] _add_map_x_72_data_near;
  wire _add_map_x_72_wall_t_out;
  wire [9:0] _add_map_x_72_data_org;
  wire [9:0] _add_map_x_72_data_org_near;
  wire [1:0] _add_map_x_72_s_g;
  wire [1:0] _add_map_x_72_s_g_near;
  wire _add_map_x_72_add_exe;
  wire _add_map_x_72_p_reset;
  wire _add_map_x_72_m_clock;
  wire [9:0] _add_map_x_71_moto_org_near;
  wire [9:0] _add_map_x_71_moto_org_near1;
  wire [9:0] _add_map_x_71_moto_org_near2;
  wire [9:0] _add_map_x_71_moto_org_near3;
  wire [9:0] _add_map_x_71_moto_org;
  wire [1:0] _add_map_x_71_sg_up;
  wire [1:0] _add_map_x_71_sg_down;
  wire [1:0] _add_map_x_71_sg_left;
  wire [1:0] _add_map_x_71_sg_right;
  wire _add_map_x_71_wall_t_in;
  wire [9:0] _add_map_x_71_moto;
  wire [9:0] _add_map_x_71_up;
  wire [9:0] _add_map_x_71_right;
  wire [9:0] _add_map_x_71_down;
  wire [9:0] _add_map_x_71_left;
  wire [9:0] _add_map_x_71_start;
  wire [9:0] _add_map_x_71_goal;
  wire [9:0] _add_map_x_71_now;
  wire [9:0] _add_map_x_71_data_out;
  wire [9:0] _add_map_x_71_data_out_index;
  wire [9:0] _add_map_x_71_data_near;
  wire _add_map_x_71_wall_t_out;
  wire [9:0] _add_map_x_71_data_org;
  wire [9:0] _add_map_x_71_data_org_near;
  wire [1:0] _add_map_x_71_s_g;
  wire [1:0] _add_map_x_71_s_g_near;
  wire _add_map_x_71_add_exe;
  wire _add_map_x_71_p_reset;
  wire _add_map_x_71_m_clock;
  wire [9:0] _add_map_x_70_moto_org_near;
  wire [9:0] _add_map_x_70_moto_org_near1;
  wire [9:0] _add_map_x_70_moto_org_near2;
  wire [9:0] _add_map_x_70_moto_org_near3;
  wire [9:0] _add_map_x_70_moto_org;
  wire [1:0] _add_map_x_70_sg_up;
  wire [1:0] _add_map_x_70_sg_down;
  wire [1:0] _add_map_x_70_sg_left;
  wire [1:0] _add_map_x_70_sg_right;
  wire _add_map_x_70_wall_t_in;
  wire [9:0] _add_map_x_70_moto;
  wire [9:0] _add_map_x_70_up;
  wire [9:0] _add_map_x_70_right;
  wire [9:0] _add_map_x_70_down;
  wire [9:0] _add_map_x_70_left;
  wire [9:0] _add_map_x_70_start;
  wire [9:0] _add_map_x_70_goal;
  wire [9:0] _add_map_x_70_now;
  wire [9:0] _add_map_x_70_data_out;
  wire [9:0] _add_map_x_70_data_out_index;
  wire [9:0] _add_map_x_70_data_near;
  wire _add_map_x_70_wall_t_out;
  wire [9:0] _add_map_x_70_data_org;
  wire [9:0] _add_map_x_70_data_org_near;
  wire [1:0] _add_map_x_70_s_g;
  wire [1:0] _add_map_x_70_s_g_near;
  wire _add_map_x_70_add_exe;
  wire _add_map_x_70_p_reset;
  wire _add_map_x_70_m_clock;
  wire [9:0] _add_map_x_69_moto_org_near;
  wire [9:0] _add_map_x_69_moto_org_near1;
  wire [9:0] _add_map_x_69_moto_org_near2;
  wire [9:0] _add_map_x_69_moto_org_near3;
  wire [9:0] _add_map_x_69_moto_org;
  wire [1:0] _add_map_x_69_sg_up;
  wire [1:0] _add_map_x_69_sg_down;
  wire [1:0] _add_map_x_69_sg_left;
  wire [1:0] _add_map_x_69_sg_right;
  wire _add_map_x_69_wall_t_in;
  wire [9:0] _add_map_x_69_moto;
  wire [9:0] _add_map_x_69_up;
  wire [9:0] _add_map_x_69_right;
  wire [9:0] _add_map_x_69_down;
  wire [9:0] _add_map_x_69_left;
  wire [9:0] _add_map_x_69_start;
  wire [9:0] _add_map_x_69_goal;
  wire [9:0] _add_map_x_69_now;
  wire [9:0] _add_map_x_69_data_out;
  wire [9:0] _add_map_x_69_data_out_index;
  wire [9:0] _add_map_x_69_data_near;
  wire _add_map_x_69_wall_t_out;
  wire [9:0] _add_map_x_69_data_org;
  wire [9:0] _add_map_x_69_data_org_near;
  wire [1:0] _add_map_x_69_s_g;
  wire [1:0] _add_map_x_69_s_g_near;
  wire _add_map_x_69_add_exe;
  wire _add_map_x_69_p_reset;
  wire _add_map_x_69_m_clock;
  wire [9:0] _add_map_x_68_moto_org_near;
  wire [9:0] _add_map_x_68_moto_org_near1;
  wire [9:0] _add_map_x_68_moto_org_near2;
  wire [9:0] _add_map_x_68_moto_org_near3;
  wire [9:0] _add_map_x_68_moto_org;
  wire [1:0] _add_map_x_68_sg_up;
  wire [1:0] _add_map_x_68_sg_down;
  wire [1:0] _add_map_x_68_sg_left;
  wire [1:0] _add_map_x_68_sg_right;
  wire _add_map_x_68_wall_t_in;
  wire [9:0] _add_map_x_68_moto;
  wire [9:0] _add_map_x_68_up;
  wire [9:0] _add_map_x_68_right;
  wire [9:0] _add_map_x_68_down;
  wire [9:0] _add_map_x_68_left;
  wire [9:0] _add_map_x_68_start;
  wire [9:0] _add_map_x_68_goal;
  wire [9:0] _add_map_x_68_now;
  wire [9:0] _add_map_x_68_data_out;
  wire [9:0] _add_map_x_68_data_out_index;
  wire [9:0] _add_map_x_68_data_near;
  wire _add_map_x_68_wall_t_out;
  wire [9:0] _add_map_x_68_data_org;
  wire [9:0] _add_map_x_68_data_org_near;
  wire [1:0] _add_map_x_68_s_g;
  wire [1:0] _add_map_x_68_s_g_near;
  wire _add_map_x_68_add_exe;
  wire _add_map_x_68_p_reset;
  wire _add_map_x_68_m_clock;
  wire [9:0] _add_map_x_67_moto_org_near;
  wire [9:0] _add_map_x_67_moto_org_near1;
  wire [9:0] _add_map_x_67_moto_org_near2;
  wire [9:0] _add_map_x_67_moto_org_near3;
  wire [9:0] _add_map_x_67_moto_org;
  wire [1:0] _add_map_x_67_sg_up;
  wire [1:0] _add_map_x_67_sg_down;
  wire [1:0] _add_map_x_67_sg_left;
  wire [1:0] _add_map_x_67_sg_right;
  wire _add_map_x_67_wall_t_in;
  wire [9:0] _add_map_x_67_moto;
  wire [9:0] _add_map_x_67_up;
  wire [9:0] _add_map_x_67_right;
  wire [9:0] _add_map_x_67_down;
  wire [9:0] _add_map_x_67_left;
  wire [9:0] _add_map_x_67_start;
  wire [9:0] _add_map_x_67_goal;
  wire [9:0] _add_map_x_67_now;
  wire [9:0] _add_map_x_67_data_out;
  wire [9:0] _add_map_x_67_data_out_index;
  wire [9:0] _add_map_x_67_data_near;
  wire _add_map_x_67_wall_t_out;
  wire [9:0] _add_map_x_67_data_org;
  wire [9:0] _add_map_x_67_data_org_near;
  wire [1:0] _add_map_x_67_s_g;
  wire [1:0] _add_map_x_67_s_g_near;
  wire _add_map_x_67_add_exe;
  wire _add_map_x_67_p_reset;
  wire _add_map_x_67_m_clock;
  wire [9:0] _add_map_x_66_moto_org_near;
  wire [9:0] _add_map_x_66_moto_org_near1;
  wire [9:0] _add_map_x_66_moto_org_near2;
  wire [9:0] _add_map_x_66_moto_org_near3;
  wire [9:0] _add_map_x_66_moto_org;
  wire [1:0] _add_map_x_66_sg_up;
  wire [1:0] _add_map_x_66_sg_down;
  wire [1:0] _add_map_x_66_sg_left;
  wire [1:0] _add_map_x_66_sg_right;
  wire _add_map_x_66_wall_t_in;
  wire [9:0] _add_map_x_66_moto;
  wire [9:0] _add_map_x_66_up;
  wire [9:0] _add_map_x_66_right;
  wire [9:0] _add_map_x_66_down;
  wire [9:0] _add_map_x_66_left;
  wire [9:0] _add_map_x_66_start;
  wire [9:0] _add_map_x_66_goal;
  wire [9:0] _add_map_x_66_now;
  wire [9:0] _add_map_x_66_data_out;
  wire [9:0] _add_map_x_66_data_out_index;
  wire [9:0] _add_map_x_66_data_near;
  wire _add_map_x_66_wall_t_out;
  wire [9:0] _add_map_x_66_data_org;
  wire [9:0] _add_map_x_66_data_org_near;
  wire [1:0] _add_map_x_66_s_g;
  wire [1:0] _add_map_x_66_s_g_near;
  wire _add_map_x_66_add_exe;
  wire _add_map_x_66_p_reset;
  wire _add_map_x_66_m_clock;
  wire [9:0] _add_map_x_65_moto_org_near;
  wire [9:0] _add_map_x_65_moto_org_near1;
  wire [9:0] _add_map_x_65_moto_org_near2;
  wire [9:0] _add_map_x_65_moto_org_near3;
  wire [9:0] _add_map_x_65_moto_org;
  wire [1:0] _add_map_x_65_sg_up;
  wire [1:0] _add_map_x_65_sg_down;
  wire [1:0] _add_map_x_65_sg_left;
  wire [1:0] _add_map_x_65_sg_right;
  wire _add_map_x_65_wall_t_in;
  wire [9:0] _add_map_x_65_moto;
  wire [9:0] _add_map_x_65_up;
  wire [9:0] _add_map_x_65_right;
  wire [9:0] _add_map_x_65_down;
  wire [9:0] _add_map_x_65_left;
  wire [9:0] _add_map_x_65_start;
  wire [9:0] _add_map_x_65_goal;
  wire [9:0] _add_map_x_65_now;
  wire [9:0] _add_map_x_65_data_out;
  wire [9:0] _add_map_x_65_data_out_index;
  wire [9:0] _add_map_x_65_data_near;
  wire _add_map_x_65_wall_t_out;
  wire [9:0] _add_map_x_65_data_org;
  wire [9:0] _add_map_x_65_data_org_near;
  wire [1:0] _add_map_x_65_s_g;
  wire [1:0] _add_map_x_65_s_g_near;
  wire _add_map_x_65_add_exe;
  wire _add_map_x_65_p_reset;
  wire _add_map_x_65_m_clock;
  wire [9:0] _add_map_x_64_moto_org_near;
  wire [9:0] _add_map_x_64_moto_org_near1;
  wire [9:0] _add_map_x_64_moto_org_near2;
  wire [9:0] _add_map_x_64_moto_org_near3;
  wire [9:0] _add_map_x_64_moto_org;
  wire [1:0] _add_map_x_64_sg_up;
  wire [1:0] _add_map_x_64_sg_down;
  wire [1:0] _add_map_x_64_sg_left;
  wire [1:0] _add_map_x_64_sg_right;
  wire _add_map_x_64_wall_t_in;
  wire [9:0] _add_map_x_64_moto;
  wire [9:0] _add_map_x_64_up;
  wire [9:0] _add_map_x_64_right;
  wire [9:0] _add_map_x_64_down;
  wire [9:0] _add_map_x_64_left;
  wire [9:0] _add_map_x_64_start;
  wire [9:0] _add_map_x_64_goal;
  wire [9:0] _add_map_x_64_now;
  wire [9:0] _add_map_x_64_data_out;
  wire [9:0] _add_map_x_64_data_out_index;
  wire [9:0] _add_map_x_64_data_near;
  wire _add_map_x_64_wall_t_out;
  wire [9:0] _add_map_x_64_data_org;
  wire [9:0] _add_map_x_64_data_org_near;
  wire [1:0] _add_map_x_64_s_g;
  wire [1:0] _add_map_x_64_s_g_near;
  wire _add_map_x_64_add_exe;
  wire _add_map_x_64_p_reset;
  wire _add_map_x_64_m_clock;
  wire [9:0] _add_map_x_63_moto_org_near;
  wire [9:0] _add_map_x_63_moto_org_near1;
  wire [9:0] _add_map_x_63_moto_org_near2;
  wire [9:0] _add_map_x_63_moto_org_near3;
  wire [9:0] _add_map_x_63_moto_org;
  wire [1:0] _add_map_x_63_sg_up;
  wire [1:0] _add_map_x_63_sg_down;
  wire [1:0] _add_map_x_63_sg_left;
  wire [1:0] _add_map_x_63_sg_right;
  wire _add_map_x_63_wall_t_in;
  wire [9:0] _add_map_x_63_moto;
  wire [9:0] _add_map_x_63_up;
  wire [9:0] _add_map_x_63_right;
  wire [9:0] _add_map_x_63_down;
  wire [9:0] _add_map_x_63_left;
  wire [9:0] _add_map_x_63_start;
  wire [9:0] _add_map_x_63_goal;
  wire [9:0] _add_map_x_63_now;
  wire [9:0] _add_map_x_63_data_out;
  wire [9:0] _add_map_x_63_data_out_index;
  wire [9:0] _add_map_x_63_data_near;
  wire _add_map_x_63_wall_t_out;
  wire [9:0] _add_map_x_63_data_org;
  wire [9:0] _add_map_x_63_data_org_near;
  wire [1:0] _add_map_x_63_s_g;
  wire [1:0] _add_map_x_63_s_g_near;
  wire _add_map_x_63_add_exe;
  wire _add_map_x_63_p_reset;
  wire _add_map_x_63_m_clock;
  wire [9:0] _add_map_x_62_moto_org_near;
  wire [9:0] _add_map_x_62_moto_org_near1;
  wire [9:0] _add_map_x_62_moto_org_near2;
  wire [9:0] _add_map_x_62_moto_org_near3;
  wire [9:0] _add_map_x_62_moto_org;
  wire [1:0] _add_map_x_62_sg_up;
  wire [1:0] _add_map_x_62_sg_down;
  wire [1:0] _add_map_x_62_sg_left;
  wire [1:0] _add_map_x_62_sg_right;
  wire _add_map_x_62_wall_t_in;
  wire [9:0] _add_map_x_62_moto;
  wire [9:0] _add_map_x_62_up;
  wire [9:0] _add_map_x_62_right;
  wire [9:0] _add_map_x_62_down;
  wire [9:0] _add_map_x_62_left;
  wire [9:0] _add_map_x_62_start;
  wire [9:0] _add_map_x_62_goal;
  wire [9:0] _add_map_x_62_now;
  wire [9:0] _add_map_x_62_data_out;
  wire [9:0] _add_map_x_62_data_out_index;
  wire [9:0] _add_map_x_62_data_near;
  wire _add_map_x_62_wall_t_out;
  wire [9:0] _add_map_x_62_data_org;
  wire [9:0] _add_map_x_62_data_org_near;
  wire [1:0] _add_map_x_62_s_g;
  wire [1:0] _add_map_x_62_s_g_near;
  wire _add_map_x_62_add_exe;
  wire _add_map_x_62_p_reset;
  wire _add_map_x_62_m_clock;
  wire [9:0] _add_map_x_61_moto_org_near;
  wire [9:0] _add_map_x_61_moto_org_near1;
  wire [9:0] _add_map_x_61_moto_org_near2;
  wire [9:0] _add_map_x_61_moto_org_near3;
  wire [9:0] _add_map_x_61_moto_org;
  wire [1:0] _add_map_x_61_sg_up;
  wire [1:0] _add_map_x_61_sg_down;
  wire [1:0] _add_map_x_61_sg_left;
  wire [1:0] _add_map_x_61_sg_right;
  wire _add_map_x_61_wall_t_in;
  wire [9:0] _add_map_x_61_moto;
  wire [9:0] _add_map_x_61_up;
  wire [9:0] _add_map_x_61_right;
  wire [9:0] _add_map_x_61_down;
  wire [9:0] _add_map_x_61_left;
  wire [9:0] _add_map_x_61_start;
  wire [9:0] _add_map_x_61_goal;
  wire [9:0] _add_map_x_61_now;
  wire [9:0] _add_map_x_61_data_out;
  wire [9:0] _add_map_x_61_data_out_index;
  wire [9:0] _add_map_x_61_data_near;
  wire _add_map_x_61_wall_t_out;
  wire [9:0] _add_map_x_61_data_org;
  wire [9:0] _add_map_x_61_data_org_near;
  wire [1:0] _add_map_x_61_s_g;
  wire [1:0] _add_map_x_61_s_g_near;
  wire _add_map_x_61_add_exe;
  wire _add_map_x_61_p_reset;
  wire _add_map_x_61_m_clock;
  wire [9:0] _add_map_x_60_moto_org_near;
  wire [9:0] _add_map_x_60_moto_org_near1;
  wire [9:0] _add_map_x_60_moto_org_near2;
  wire [9:0] _add_map_x_60_moto_org_near3;
  wire [9:0] _add_map_x_60_moto_org;
  wire [1:0] _add_map_x_60_sg_up;
  wire [1:0] _add_map_x_60_sg_down;
  wire [1:0] _add_map_x_60_sg_left;
  wire [1:0] _add_map_x_60_sg_right;
  wire _add_map_x_60_wall_t_in;
  wire [9:0] _add_map_x_60_moto;
  wire [9:0] _add_map_x_60_up;
  wire [9:0] _add_map_x_60_right;
  wire [9:0] _add_map_x_60_down;
  wire [9:0] _add_map_x_60_left;
  wire [9:0] _add_map_x_60_start;
  wire [9:0] _add_map_x_60_goal;
  wire [9:0] _add_map_x_60_now;
  wire [9:0] _add_map_x_60_data_out;
  wire [9:0] _add_map_x_60_data_out_index;
  wire [9:0] _add_map_x_60_data_near;
  wire _add_map_x_60_wall_t_out;
  wire [9:0] _add_map_x_60_data_org;
  wire [9:0] _add_map_x_60_data_org_near;
  wire [1:0] _add_map_x_60_s_g;
  wire [1:0] _add_map_x_60_s_g_near;
  wire _add_map_x_60_add_exe;
  wire _add_map_x_60_p_reset;
  wire _add_map_x_60_m_clock;
  wire [9:0] _add_map_x_59_moto_org_near;
  wire [9:0] _add_map_x_59_moto_org_near1;
  wire [9:0] _add_map_x_59_moto_org_near2;
  wire [9:0] _add_map_x_59_moto_org_near3;
  wire [9:0] _add_map_x_59_moto_org;
  wire [1:0] _add_map_x_59_sg_up;
  wire [1:0] _add_map_x_59_sg_down;
  wire [1:0] _add_map_x_59_sg_left;
  wire [1:0] _add_map_x_59_sg_right;
  wire _add_map_x_59_wall_t_in;
  wire [9:0] _add_map_x_59_moto;
  wire [9:0] _add_map_x_59_up;
  wire [9:0] _add_map_x_59_right;
  wire [9:0] _add_map_x_59_down;
  wire [9:0] _add_map_x_59_left;
  wire [9:0] _add_map_x_59_start;
  wire [9:0] _add_map_x_59_goal;
  wire [9:0] _add_map_x_59_now;
  wire [9:0] _add_map_x_59_data_out;
  wire [9:0] _add_map_x_59_data_out_index;
  wire [9:0] _add_map_x_59_data_near;
  wire _add_map_x_59_wall_t_out;
  wire [9:0] _add_map_x_59_data_org;
  wire [9:0] _add_map_x_59_data_org_near;
  wire [1:0] _add_map_x_59_s_g;
  wire [1:0] _add_map_x_59_s_g_near;
  wire _add_map_x_59_add_exe;
  wire _add_map_x_59_p_reset;
  wire _add_map_x_59_m_clock;
  wire [9:0] _add_map_x_58_moto_org_near;
  wire [9:0] _add_map_x_58_moto_org_near1;
  wire [9:0] _add_map_x_58_moto_org_near2;
  wire [9:0] _add_map_x_58_moto_org_near3;
  wire [9:0] _add_map_x_58_moto_org;
  wire [1:0] _add_map_x_58_sg_up;
  wire [1:0] _add_map_x_58_sg_down;
  wire [1:0] _add_map_x_58_sg_left;
  wire [1:0] _add_map_x_58_sg_right;
  wire _add_map_x_58_wall_t_in;
  wire [9:0] _add_map_x_58_moto;
  wire [9:0] _add_map_x_58_up;
  wire [9:0] _add_map_x_58_right;
  wire [9:0] _add_map_x_58_down;
  wire [9:0] _add_map_x_58_left;
  wire [9:0] _add_map_x_58_start;
  wire [9:0] _add_map_x_58_goal;
  wire [9:0] _add_map_x_58_now;
  wire [9:0] _add_map_x_58_data_out;
  wire [9:0] _add_map_x_58_data_out_index;
  wire [9:0] _add_map_x_58_data_near;
  wire _add_map_x_58_wall_t_out;
  wire [9:0] _add_map_x_58_data_org;
  wire [9:0] _add_map_x_58_data_org_near;
  wire [1:0] _add_map_x_58_s_g;
  wire [1:0] _add_map_x_58_s_g_near;
  wire _add_map_x_58_add_exe;
  wire _add_map_x_58_p_reset;
  wire _add_map_x_58_m_clock;
  wire [9:0] _add_map_x_57_moto_org_near;
  wire [9:0] _add_map_x_57_moto_org_near1;
  wire [9:0] _add_map_x_57_moto_org_near2;
  wire [9:0] _add_map_x_57_moto_org_near3;
  wire [9:0] _add_map_x_57_moto_org;
  wire [1:0] _add_map_x_57_sg_up;
  wire [1:0] _add_map_x_57_sg_down;
  wire [1:0] _add_map_x_57_sg_left;
  wire [1:0] _add_map_x_57_sg_right;
  wire _add_map_x_57_wall_t_in;
  wire [9:0] _add_map_x_57_moto;
  wire [9:0] _add_map_x_57_up;
  wire [9:0] _add_map_x_57_right;
  wire [9:0] _add_map_x_57_down;
  wire [9:0] _add_map_x_57_left;
  wire [9:0] _add_map_x_57_start;
  wire [9:0] _add_map_x_57_goal;
  wire [9:0] _add_map_x_57_now;
  wire [9:0] _add_map_x_57_data_out;
  wire [9:0] _add_map_x_57_data_out_index;
  wire [9:0] _add_map_x_57_data_near;
  wire _add_map_x_57_wall_t_out;
  wire [9:0] _add_map_x_57_data_org;
  wire [9:0] _add_map_x_57_data_org_near;
  wire [1:0] _add_map_x_57_s_g;
  wire [1:0] _add_map_x_57_s_g_near;
  wire _add_map_x_57_add_exe;
  wire _add_map_x_57_p_reset;
  wire _add_map_x_57_m_clock;
  wire [9:0] _add_map_x_56_moto_org_near;
  wire [9:0] _add_map_x_56_moto_org_near1;
  wire [9:0] _add_map_x_56_moto_org_near2;
  wire [9:0] _add_map_x_56_moto_org_near3;
  wire [9:0] _add_map_x_56_moto_org;
  wire [1:0] _add_map_x_56_sg_up;
  wire [1:0] _add_map_x_56_sg_down;
  wire [1:0] _add_map_x_56_sg_left;
  wire [1:0] _add_map_x_56_sg_right;
  wire _add_map_x_56_wall_t_in;
  wire [9:0] _add_map_x_56_moto;
  wire [9:0] _add_map_x_56_up;
  wire [9:0] _add_map_x_56_right;
  wire [9:0] _add_map_x_56_down;
  wire [9:0] _add_map_x_56_left;
  wire [9:0] _add_map_x_56_start;
  wire [9:0] _add_map_x_56_goal;
  wire [9:0] _add_map_x_56_now;
  wire [9:0] _add_map_x_56_data_out;
  wire [9:0] _add_map_x_56_data_out_index;
  wire [9:0] _add_map_x_56_data_near;
  wire _add_map_x_56_wall_t_out;
  wire [9:0] _add_map_x_56_data_org;
  wire [9:0] _add_map_x_56_data_org_near;
  wire [1:0] _add_map_x_56_s_g;
  wire [1:0] _add_map_x_56_s_g_near;
  wire _add_map_x_56_add_exe;
  wire _add_map_x_56_p_reset;
  wire _add_map_x_56_m_clock;
  wire [9:0] _add_map_x_55_moto_org_near;
  wire [9:0] _add_map_x_55_moto_org_near1;
  wire [9:0] _add_map_x_55_moto_org_near2;
  wire [9:0] _add_map_x_55_moto_org_near3;
  wire [9:0] _add_map_x_55_moto_org;
  wire [1:0] _add_map_x_55_sg_up;
  wire [1:0] _add_map_x_55_sg_down;
  wire [1:0] _add_map_x_55_sg_left;
  wire [1:0] _add_map_x_55_sg_right;
  wire _add_map_x_55_wall_t_in;
  wire [9:0] _add_map_x_55_moto;
  wire [9:0] _add_map_x_55_up;
  wire [9:0] _add_map_x_55_right;
  wire [9:0] _add_map_x_55_down;
  wire [9:0] _add_map_x_55_left;
  wire [9:0] _add_map_x_55_start;
  wire [9:0] _add_map_x_55_goal;
  wire [9:0] _add_map_x_55_now;
  wire [9:0] _add_map_x_55_data_out;
  wire [9:0] _add_map_x_55_data_out_index;
  wire [9:0] _add_map_x_55_data_near;
  wire _add_map_x_55_wall_t_out;
  wire [9:0] _add_map_x_55_data_org;
  wire [9:0] _add_map_x_55_data_org_near;
  wire [1:0] _add_map_x_55_s_g;
  wire [1:0] _add_map_x_55_s_g_near;
  wire _add_map_x_55_add_exe;
  wire _add_map_x_55_p_reset;
  wire _add_map_x_55_m_clock;
  wire [9:0] _add_map_x_54_moto_org_near;
  wire [9:0] _add_map_x_54_moto_org_near1;
  wire [9:0] _add_map_x_54_moto_org_near2;
  wire [9:0] _add_map_x_54_moto_org_near3;
  wire [9:0] _add_map_x_54_moto_org;
  wire [1:0] _add_map_x_54_sg_up;
  wire [1:0] _add_map_x_54_sg_down;
  wire [1:0] _add_map_x_54_sg_left;
  wire [1:0] _add_map_x_54_sg_right;
  wire _add_map_x_54_wall_t_in;
  wire [9:0] _add_map_x_54_moto;
  wire [9:0] _add_map_x_54_up;
  wire [9:0] _add_map_x_54_right;
  wire [9:0] _add_map_x_54_down;
  wire [9:0] _add_map_x_54_left;
  wire [9:0] _add_map_x_54_start;
  wire [9:0] _add_map_x_54_goal;
  wire [9:0] _add_map_x_54_now;
  wire [9:0] _add_map_x_54_data_out;
  wire [9:0] _add_map_x_54_data_out_index;
  wire [9:0] _add_map_x_54_data_near;
  wire _add_map_x_54_wall_t_out;
  wire [9:0] _add_map_x_54_data_org;
  wire [9:0] _add_map_x_54_data_org_near;
  wire [1:0] _add_map_x_54_s_g;
  wire [1:0] _add_map_x_54_s_g_near;
  wire _add_map_x_54_add_exe;
  wire _add_map_x_54_p_reset;
  wire _add_map_x_54_m_clock;
  wire [9:0] _add_map_x_53_moto_org_near;
  wire [9:0] _add_map_x_53_moto_org_near1;
  wire [9:0] _add_map_x_53_moto_org_near2;
  wire [9:0] _add_map_x_53_moto_org_near3;
  wire [9:0] _add_map_x_53_moto_org;
  wire [1:0] _add_map_x_53_sg_up;
  wire [1:0] _add_map_x_53_sg_down;
  wire [1:0] _add_map_x_53_sg_left;
  wire [1:0] _add_map_x_53_sg_right;
  wire _add_map_x_53_wall_t_in;
  wire [9:0] _add_map_x_53_moto;
  wire [9:0] _add_map_x_53_up;
  wire [9:0] _add_map_x_53_right;
  wire [9:0] _add_map_x_53_down;
  wire [9:0] _add_map_x_53_left;
  wire [9:0] _add_map_x_53_start;
  wire [9:0] _add_map_x_53_goal;
  wire [9:0] _add_map_x_53_now;
  wire [9:0] _add_map_x_53_data_out;
  wire [9:0] _add_map_x_53_data_out_index;
  wire [9:0] _add_map_x_53_data_near;
  wire _add_map_x_53_wall_t_out;
  wire [9:0] _add_map_x_53_data_org;
  wire [9:0] _add_map_x_53_data_org_near;
  wire [1:0] _add_map_x_53_s_g;
  wire [1:0] _add_map_x_53_s_g_near;
  wire _add_map_x_53_add_exe;
  wire _add_map_x_53_p_reset;
  wire _add_map_x_53_m_clock;
  wire [9:0] _add_map_x_52_moto_org_near;
  wire [9:0] _add_map_x_52_moto_org_near1;
  wire [9:0] _add_map_x_52_moto_org_near2;
  wire [9:0] _add_map_x_52_moto_org_near3;
  wire [9:0] _add_map_x_52_moto_org;
  wire [1:0] _add_map_x_52_sg_up;
  wire [1:0] _add_map_x_52_sg_down;
  wire [1:0] _add_map_x_52_sg_left;
  wire [1:0] _add_map_x_52_sg_right;
  wire _add_map_x_52_wall_t_in;
  wire [9:0] _add_map_x_52_moto;
  wire [9:0] _add_map_x_52_up;
  wire [9:0] _add_map_x_52_right;
  wire [9:0] _add_map_x_52_down;
  wire [9:0] _add_map_x_52_left;
  wire [9:0] _add_map_x_52_start;
  wire [9:0] _add_map_x_52_goal;
  wire [9:0] _add_map_x_52_now;
  wire [9:0] _add_map_x_52_data_out;
  wire [9:0] _add_map_x_52_data_out_index;
  wire [9:0] _add_map_x_52_data_near;
  wire _add_map_x_52_wall_t_out;
  wire [9:0] _add_map_x_52_data_org;
  wire [9:0] _add_map_x_52_data_org_near;
  wire [1:0] _add_map_x_52_s_g;
  wire [1:0] _add_map_x_52_s_g_near;
  wire _add_map_x_52_add_exe;
  wire _add_map_x_52_p_reset;
  wire _add_map_x_52_m_clock;
  wire [9:0] _add_map_x_51_moto_org_near;
  wire [9:0] _add_map_x_51_moto_org_near1;
  wire [9:0] _add_map_x_51_moto_org_near2;
  wire [9:0] _add_map_x_51_moto_org_near3;
  wire [9:0] _add_map_x_51_moto_org;
  wire [1:0] _add_map_x_51_sg_up;
  wire [1:0] _add_map_x_51_sg_down;
  wire [1:0] _add_map_x_51_sg_left;
  wire [1:0] _add_map_x_51_sg_right;
  wire _add_map_x_51_wall_t_in;
  wire [9:0] _add_map_x_51_moto;
  wire [9:0] _add_map_x_51_up;
  wire [9:0] _add_map_x_51_right;
  wire [9:0] _add_map_x_51_down;
  wire [9:0] _add_map_x_51_left;
  wire [9:0] _add_map_x_51_start;
  wire [9:0] _add_map_x_51_goal;
  wire [9:0] _add_map_x_51_now;
  wire [9:0] _add_map_x_51_data_out;
  wire [9:0] _add_map_x_51_data_out_index;
  wire [9:0] _add_map_x_51_data_near;
  wire _add_map_x_51_wall_t_out;
  wire [9:0] _add_map_x_51_data_org;
  wire [9:0] _add_map_x_51_data_org_near;
  wire [1:0] _add_map_x_51_s_g;
  wire [1:0] _add_map_x_51_s_g_near;
  wire _add_map_x_51_add_exe;
  wire _add_map_x_51_p_reset;
  wire _add_map_x_51_m_clock;
  wire [9:0] _add_map_x_50_moto_org_near;
  wire [9:0] _add_map_x_50_moto_org_near1;
  wire [9:0] _add_map_x_50_moto_org_near2;
  wire [9:0] _add_map_x_50_moto_org_near3;
  wire [9:0] _add_map_x_50_moto_org;
  wire [1:0] _add_map_x_50_sg_up;
  wire [1:0] _add_map_x_50_sg_down;
  wire [1:0] _add_map_x_50_sg_left;
  wire [1:0] _add_map_x_50_sg_right;
  wire _add_map_x_50_wall_t_in;
  wire [9:0] _add_map_x_50_moto;
  wire [9:0] _add_map_x_50_up;
  wire [9:0] _add_map_x_50_right;
  wire [9:0] _add_map_x_50_down;
  wire [9:0] _add_map_x_50_left;
  wire [9:0] _add_map_x_50_start;
  wire [9:0] _add_map_x_50_goal;
  wire [9:0] _add_map_x_50_now;
  wire [9:0] _add_map_x_50_data_out;
  wire [9:0] _add_map_x_50_data_out_index;
  wire [9:0] _add_map_x_50_data_near;
  wire _add_map_x_50_wall_t_out;
  wire [9:0] _add_map_x_50_data_org;
  wire [9:0] _add_map_x_50_data_org_near;
  wire [1:0] _add_map_x_50_s_g;
  wire [1:0] _add_map_x_50_s_g_near;
  wire _add_map_x_50_add_exe;
  wire _add_map_x_50_p_reset;
  wire _add_map_x_50_m_clock;
  wire [9:0] _add_map_x_49_moto_org_near;
  wire [9:0] _add_map_x_49_moto_org_near1;
  wire [9:0] _add_map_x_49_moto_org_near2;
  wire [9:0] _add_map_x_49_moto_org_near3;
  wire [9:0] _add_map_x_49_moto_org;
  wire [1:0] _add_map_x_49_sg_up;
  wire [1:0] _add_map_x_49_sg_down;
  wire [1:0] _add_map_x_49_sg_left;
  wire [1:0] _add_map_x_49_sg_right;
  wire _add_map_x_49_wall_t_in;
  wire [9:0] _add_map_x_49_moto;
  wire [9:0] _add_map_x_49_up;
  wire [9:0] _add_map_x_49_right;
  wire [9:0] _add_map_x_49_down;
  wire [9:0] _add_map_x_49_left;
  wire [9:0] _add_map_x_49_start;
  wire [9:0] _add_map_x_49_goal;
  wire [9:0] _add_map_x_49_now;
  wire [9:0] _add_map_x_49_data_out;
  wire [9:0] _add_map_x_49_data_out_index;
  wire [9:0] _add_map_x_49_data_near;
  wire _add_map_x_49_wall_t_out;
  wire [9:0] _add_map_x_49_data_org;
  wire [9:0] _add_map_x_49_data_org_near;
  wire [1:0] _add_map_x_49_s_g;
  wire [1:0] _add_map_x_49_s_g_near;
  wire _add_map_x_49_add_exe;
  wire _add_map_x_49_p_reset;
  wire _add_map_x_49_m_clock;
  wire [9:0] _add_map_x_48_moto_org_near;
  wire [9:0] _add_map_x_48_moto_org_near1;
  wire [9:0] _add_map_x_48_moto_org_near2;
  wire [9:0] _add_map_x_48_moto_org_near3;
  wire [9:0] _add_map_x_48_moto_org;
  wire [1:0] _add_map_x_48_sg_up;
  wire [1:0] _add_map_x_48_sg_down;
  wire [1:0] _add_map_x_48_sg_left;
  wire [1:0] _add_map_x_48_sg_right;
  wire _add_map_x_48_wall_t_in;
  wire [9:0] _add_map_x_48_moto;
  wire [9:0] _add_map_x_48_up;
  wire [9:0] _add_map_x_48_right;
  wire [9:0] _add_map_x_48_down;
  wire [9:0] _add_map_x_48_left;
  wire [9:0] _add_map_x_48_start;
  wire [9:0] _add_map_x_48_goal;
  wire [9:0] _add_map_x_48_now;
  wire [9:0] _add_map_x_48_data_out;
  wire [9:0] _add_map_x_48_data_out_index;
  wire [9:0] _add_map_x_48_data_near;
  wire _add_map_x_48_wall_t_out;
  wire [9:0] _add_map_x_48_data_org;
  wire [9:0] _add_map_x_48_data_org_near;
  wire [1:0] _add_map_x_48_s_g;
  wire [1:0] _add_map_x_48_s_g_near;
  wire _add_map_x_48_add_exe;
  wire _add_map_x_48_p_reset;
  wire _add_map_x_48_m_clock;
  wire [9:0] _add_map_x_47_moto_org_near;
  wire [9:0] _add_map_x_47_moto_org_near1;
  wire [9:0] _add_map_x_47_moto_org_near2;
  wire [9:0] _add_map_x_47_moto_org_near3;
  wire [9:0] _add_map_x_47_moto_org;
  wire [1:0] _add_map_x_47_sg_up;
  wire [1:0] _add_map_x_47_sg_down;
  wire [1:0] _add_map_x_47_sg_left;
  wire [1:0] _add_map_x_47_sg_right;
  wire _add_map_x_47_wall_t_in;
  wire [9:0] _add_map_x_47_moto;
  wire [9:0] _add_map_x_47_up;
  wire [9:0] _add_map_x_47_right;
  wire [9:0] _add_map_x_47_down;
  wire [9:0] _add_map_x_47_left;
  wire [9:0] _add_map_x_47_start;
  wire [9:0] _add_map_x_47_goal;
  wire [9:0] _add_map_x_47_now;
  wire [9:0] _add_map_x_47_data_out;
  wire [9:0] _add_map_x_47_data_out_index;
  wire [9:0] _add_map_x_47_data_near;
  wire _add_map_x_47_wall_t_out;
  wire [9:0] _add_map_x_47_data_org;
  wire [9:0] _add_map_x_47_data_org_near;
  wire [1:0] _add_map_x_47_s_g;
  wire [1:0] _add_map_x_47_s_g_near;
  wire _add_map_x_47_add_exe;
  wire _add_map_x_47_p_reset;
  wire _add_map_x_47_m_clock;
  wire [9:0] _add_map_x_46_moto_org_near;
  wire [9:0] _add_map_x_46_moto_org_near1;
  wire [9:0] _add_map_x_46_moto_org_near2;
  wire [9:0] _add_map_x_46_moto_org_near3;
  wire [9:0] _add_map_x_46_moto_org;
  wire [1:0] _add_map_x_46_sg_up;
  wire [1:0] _add_map_x_46_sg_down;
  wire [1:0] _add_map_x_46_sg_left;
  wire [1:0] _add_map_x_46_sg_right;
  wire _add_map_x_46_wall_t_in;
  wire [9:0] _add_map_x_46_moto;
  wire [9:0] _add_map_x_46_up;
  wire [9:0] _add_map_x_46_right;
  wire [9:0] _add_map_x_46_down;
  wire [9:0] _add_map_x_46_left;
  wire [9:0] _add_map_x_46_start;
  wire [9:0] _add_map_x_46_goal;
  wire [9:0] _add_map_x_46_now;
  wire [9:0] _add_map_x_46_data_out;
  wire [9:0] _add_map_x_46_data_out_index;
  wire [9:0] _add_map_x_46_data_near;
  wire _add_map_x_46_wall_t_out;
  wire [9:0] _add_map_x_46_data_org;
  wire [9:0] _add_map_x_46_data_org_near;
  wire [1:0] _add_map_x_46_s_g;
  wire [1:0] _add_map_x_46_s_g_near;
  wire _add_map_x_46_add_exe;
  wire _add_map_x_46_p_reset;
  wire _add_map_x_46_m_clock;
  wire [9:0] _add_map_x_45_moto_org_near;
  wire [9:0] _add_map_x_45_moto_org_near1;
  wire [9:0] _add_map_x_45_moto_org_near2;
  wire [9:0] _add_map_x_45_moto_org_near3;
  wire [9:0] _add_map_x_45_moto_org;
  wire [1:0] _add_map_x_45_sg_up;
  wire [1:0] _add_map_x_45_sg_down;
  wire [1:0] _add_map_x_45_sg_left;
  wire [1:0] _add_map_x_45_sg_right;
  wire _add_map_x_45_wall_t_in;
  wire [9:0] _add_map_x_45_moto;
  wire [9:0] _add_map_x_45_up;
  wire [9:0] _add_map_x_45_right;
  wire [9:0] _add_map_x_45_down;
  wire [9:0] _add_map_x_45_left;
  wire [9:0] _add_map_x_45_start;
  wire [9:0] _add_map_x_45_goal;
  wire [9:0] _add_map_x_45_now;
  wire [9:0] _add_map_x_45_data_out;
  wire [9:0] _add_map_x_45_data_out_index;
  wire [9:0] _add_map_x_45_data_near;
  wire _add_map_x_45_wall_t_out;
  wire [9:0] _add_map_x_45_data_org;
  wire [9:0] _add_map_x_45_data_org_near;
  wire [1:0] _add_map_x_45_s_g;
  wire [1:0] _add_map_x_45_s_g_near;
  wire _add_map_x_45_add_exe;
  wire _add_map_x_45_p_reset;
  wire _add_map_x_45_m_clock;
  wire [9:0] _add_map_x_44_moto_org_near;
  wire [9:0] _add_map_x_44_moto_org_near1;
  wire [9:0] _add_map_x_44_moto_org_near2;
  wire [9:0] _add_map_x_44_moto_org_near3;
  wire [9:0] _add_map_x_44_moto_org;
  wire [1:0] _add_map_x_44_sg_up;
  wire [1:0] _add_map_x_44_sg_down;
  wire [1:0] _add_map_x_44_sg_left;
  wire [1:0] _add_map_x_44_sg_right;
  wire _add_map_x_44_wall_t_in;
  wire [9:0] _add_map_x_44_moto;
  wire [9:0] _add_map_x_44_up;
  wire [9:0] _add_map_x_44_right;
  wire [9:0] _add_map_x_44_down;
  wire [9:0] _add_map_x_44_left;
  wire [9:0] _add_map_x_44_start;
  wire [9:0] _add_map_x_44_goal;
  wire [9:0] _add_map_x_44_now;
  wire [9:0] _add_map_x_44_data_out;
  wire [9:0] _add_map_x_44_data_out_index;
  wire [9:0] _add_map_x_44_data_near;
  wire _add_map_x_44_wall_t_out;
  wire [9:0] _add_map_x_44_data_org;
  wire [9:0] _add_map_x_44_data_org_near;
  wire [1:0] _add_map_x_44_s_g;
  wire [1:0] _add_map_x_44_s_g_near;
  wire _add_map_x_44_add_exe;
  wire _add_map_x_44_p_reset;
  wire _add_map_x_44_m_clock;
  wire [9:0] _add_map_x_43_moto_org_near;
  wire [9:0] _add_map_x_43_moto_org_near1;
  wire [9:0] _add_map_x_43_moto_org_near2;
  wire [9:0] _add_map_x_43_moto_org_near3;
  wire [9:0] _add_map_x_43_moto_org;
  wire [1:0] _add_map_x_43_sg_up;
  wire [1:0] _add_map_x_43_sg_down;
  wire [1:0] _add_map_x_43_sg_left;
  wire [1:0] _add_map_x_43_sg_right;
  wire _add_map_x_43_wall_t_in;
  wire [9:0] _add_map_x_43_moto;
  wire [9:0] _add_map_x_43_up;
  wire [9:0] _add_map_x_43_right;
  wire [9:0] _add_map_x_43_down;
  wire [9:0] _add_map_x_43_left;
  wire [9:0] _add_map_x_43_start;
  wire [9:0] _add_map_x_43_goal;
  wire [9:0] _add_map_x_43_now;
  wire [9:0] _add_map_x_43_data_out;
  wire [9:0] _add_map_x_43_data_out_index;
  wire [9:0] _add_map_x_43_data_near;
  wire _add_map_x_43_wall_t_out;
  wire [9:0] _add_map_x_43_data_org;
  wire [9:0] _add_map_x_43_data_org_near;
  wire [1:0] _add_map_x_43_s_g;
  wire [1:0] _add_map_x_43_s_g_near;
  wire _add_map_x_43_add_exe;
  wire _add_map_x_43_p_reset;
  wire _add_map_x_43_m_clock;
  wire [9:0] _add_map_x_42_moto_org_near;
  wire [9:0] _add_map_x_42_moto_org_near1;
  wire [9:0] _add_map_x_42_moto_org_near2;
  wire [9:0] _add_map_x_42_moto_org_near3;
  wire [9:0] _add_map_x_42_moto_org;
  wire [1:0] _add_map_x_42_sg_up;
  wire [1:0] _add_map_x_42_sg_down;
  wire [1:0] _add_map_x_42_sg_left;
  wire [1:0] _add_map_x_42_sg_right;
  wire _add_map_x_42_wall_t_in;
  wire [9:0] _add_map_x_42_moto;
  wire [9:0] _add_map_x_42_up;
  wire [9:0] _add_map_x_42_right;
  wire [9:0] _add_map_x_42_down;
  wire [9:0] _add_map_x_42_left;
  wire [9:0] _add_map_x_42_start;
  wire [9:0] _add_map_x_42_goal;
  wire [9:0] _add_map_x_42_now;
  wire [9:0] _add_map_x_42_data_out;
  wire [9:0] _add_map_x_42_data_out_index;
  wire [9:0] _add_map_x_42_data_near;
  wire _add_map_x_42_wall_t_out;
  wire [9:0] _add_map_x_42_data_org;
  wire [9:0] _add_map_x_42_data_org_near;
  wire [1:0] _add_map_x_42_s_g;
  wire [1:0] _add_map_x_42_s_g_near;
  wire _add_map_x_42_add_exe;
  wire _add_map_x_42_p_reset;
  wire _add_map_x_42_m_clock;
  wire [9:0] _add_map_x_41_moto_org_near;
  wire [9:0] _add_map_x_41_moto_org_near1;
  wire [9:0] _add_map_x_41_moto_org_near2;
  wire [9:0] _add_map_x_41_moto_org_near3;
  wire [9:0] _add_map_x_41_moto_org;
  wire [1:0] _add_map_x_41_sg_up;
  wire [1:0] _add_map_x_41_sg_down;
  wire [1:0] _add_map_x_41_sg_left;
  wire [1:0] _add_map_x_41_sg_right;
  wire _add_map_x_41_wall_t_in;
  wire [9:0] _add_map_x_41_moto;
  wire [9:0] _add_map_x_41_up;
  wire [9:0] _add_map_x_41_right;
  wire [9:0] _add_map_x_41_down;
  wire [9:0] _add_map_x_41_left;
  wire [9:0] _add_map_x_41_start;
  wire [9:0] _add_map_x_41_goal;
  wire [9:0] _add_map_x_41_now;
  wire [9:0] _add_map_x_41_data_out;
  wire [9:0] _add_map_x_41_data_out_index;
  wire [9:0] _add_map_x_41_data_near;
  wire _add_map_x_41_wall_t_out;
  wire [9:0] _add_map_x_41_data_org;
  wire [9:0] _add_map_x_41_data_org_near;
  wire [1:0] _add_map_x_41_s_g;
  wire [1:0] _add_map_x_41_s_g_near;
  wire _add_map_x_41_add_exe;
  wire _add_map_x_41_p_reset;
  wire _add_map_x_41_m_clock;
  wire [9:0] _add_map_x_40_moto_org_near;
  wire [9:0] _add_map_x_40_moto_org_near1;
  wire [9:0] _add_map_x_40_moto_org_near2;
  wire [9:0] _add_map_x_40_moto_org_near3;
  wire [9:0] _add_map_x_40_moto_org;
  wire [1:0] _add_map_x_40_sg_up;
  wire [1:0] _add_map_x_40_sg_down;
  wire [1:0] _add_map_x_40_sg_left;
  wire [1:0] _add_map_x_40_sg_right;
  wire _add_map_x_40_wall_t_in;
  wire [9:0] _add_map_x_40_moto;
  wire [9:0] _add_map_x_40_up;
  wire [9:0] _add_map_x_40_right;
  wire [9:0] _add_map_x_40_down;
  wire [9:0] _add_map_x_40_left;
  wire [9:0] _add_map_x_40_start;
  wire [9:0] _add_map_x_40_goal;
  wire [9:0] _add_map_x_40_now;
  wire [9:0] _add_map_x_40_data_out;
  wire [9:0] _add_map_x_40_data_out_index;
  wire [9:0] _add_map_x_40_data_near;
  wire _add_map_x_40_wall_t_out;
  wire [9:0] _add_map_x_40_data_org;
  wire [9:0] _add_map_x_40_data_org_near;
  wire [1:0] _add_map_x_40_s_g;
  wire [1:0] _add_map_x_40_s_g_near;
  wire _add_map_x_40_add_exe;
  wire _add_map_x_40_p_reset;
  wire _add_map_x_40_m_clock;
  wire [9:0] _add_map_x_39_moto_org_near;
  wire [9:0] _add_map_x_39_moto_org_near1;
  wire [9:0] _add_map_x_39_moto_org_near2;
  wire [9:0] _add_map_x_39_moto_org_near3;
  wire [9:0] _add_map_x_39_moto_org;
  wire [1:0] _add_map_x_39_sg_up;
  wire [1:0] _add_map_x_39_sg_down;
  wire [1:0] _add_map_x_39_sg_left;
  wire [1:0] _add_map_x_39_sg_right;
  wire _add_map_x_39_wall_t_in;
  wire [9:0] _add_map_x_39_moto;
  wire [9:0] _add_map_x_39_up;
  wire [9:0] _add_map_x_39_right;
  wire [9:0] _add_map_x_39_down;
  wire [9:0] _add_map_x_39_left;
  wire [9:0] _add_map_x_39_start;
  wire [9:0] _add_map_x_39_goal;
  wire [9:0] _add_map_x_39_now;
  wire [9:0] _add_map_x_39_data_out;
  wire [9:0] _add_map_x_39_data_out_index;
  wire [9:0] _add_map_x_39_data_near;
  wire _add_map_x_39_wall_t_out;
  wire [9:0] _add_map_x_39_data_org;
  wire [9:0] _add_map_x_39_data_org_near;
  wire [1:0] _add_map_x_39_s_g;
  wire [1:0] _add_map_x_39_s_g_near;
  wire _add_map_x_39_add_exe;
  wire _add_map_x_39_p_reset;
  wire _add_map_x_39_m_clock;
  wire [9:0] _add_map_x_38_moto_org_near;
  wire [9:0] _add_map_x_38_moto_org_near1;
  wire [9:0] _add_map_x_38_moto_org_near2;
  wire [9:0] _add_map_x_38_moto_org_near3;
  wire [9:0] _add_map_x_38_moto_org;
  wire [1:0] _add_map_x_38_sg_up;
  wire [1:0] _add_map_x_38_sg_down;
  wire [1:0] _add_map_x_38_sg_left;
  wire [1:0] _add_map_x_38_sg_right;
  wire _add_map_x_38_wall_t_in;
  wire [9:0] _add_map_x_38_moto;
  wire [9:0] _add_map_x_38_up;
  wire [9:0] _add_map_x_38_right;
  wire [9:0] _add_map_x_38_down;
  wire [9:0] _add_map_x_38_left;
  wire [9:0] _add_map_x_38_start;
  wire [9:0] _add_map_x_38_goal;
  wire [9:0] _add_map_x_38_now;
  wire [9:0] _add_map_x_38_data_out;
  wire [9:0] _add_map_x_38_data_out_index;
  wire [9:0] _add_map_x_38_data_near;
  wire _add_map_x_38_wall_t_out;
  wire [9:0] _add_map_x_38_data_org;
  wire [9:0] _add_map_x_38_data_org_near;
  wire [1:0] _add_map_x_38_s_g;
  wire [1:0] _add_map_x_38_s_g_near;
  wire _add_map_x_38_add_exe;
  wire _add_map_x_38_p_reset;
  wire _add_map_x_38_m_clock;
  wire [9:0] _add_map_x_37_moto_org_near;
  wire [9:0] _add_map_x_37_moto_org_near1;
  wire [9:0] _add_map_x_37_moto_org_near2;
  wire [9:0] _add_map_x_37_moto_org_near3;
  wire [9:0] _add_map_x_37_moto_org;
  wire [1:0] _add_map_x_37_sg_up;
  wire [1:0] _add_map_x_37_sg_down;
  wire [1:0] _add_map_x_37_sg_left;
  wire [1:0] _add_map_x_37_sg_right;
  wire _add_map_x_37_wall_t_in;
  wire [9:0] _add_map_x_37_moto;
  wire [9:0] _add_map_x_37_up;
  wire [9:0] _add_map_x_37_right;
  wire [9:0] _add_map_x_37_down;
  wire [9:0] _add_map_x_37_left;
  wire [9:0] _add_map_x_37_start;
  wire [9:0] _add_map_x_37_goal;
  wire [9:0] _add_map_x_37_now;
  wire [9:0] _add_map_x_37_data_out;
  wire [9:0] _add_map_x_37_data_out_index;
  wire [9:0] _add_map_x_37_data_near;
  wire _add_map_x_37_wall_t_out;
  wire [9:0] _add_map_x_37_data_org;
  wire [9:0] _add_map_x_37_data_org_near;
  wire [1:0] _add_map_x_37_s_g;
  wire [1:0] _add_map_x_37_s_g_near;
  wire _add_map_x_37_add_exe;
  wire _add_map_x_37_p_reset;
  wire _add_map_x_37_m_clock;
  wire [9:0] _add_map_x_36_moto_org_near;
  wire [9:0] _add_map_x_36_moto_org_near1;
  wire [9:0] _add_map_x_36_moto_org_near2;
  wire [9:0] _add_map_x_36_moto_org_near3;
  wire [9:0] _add_map_x_36_moto_org;
  wire [1:0] _add_map_x_36_sg_up;
  wire [1:0] _add_map_x_36_sg_down;
  wire [1:0] _add_map_x_36_sg_left;
  wire [1:0] _add_map_x_36_sg_right;
  wire _add_map_x_36_wall_t_in;
  wire [9:0] _add_map_x_36_moto;
  wire [9:0] _add_map_x_36_up;
  wire [9:0] _add_map_x_36_right;
  wire [9:0] _add_map_x_36_down;
  wire [9:0] _add_map_x_36_left;
  wire [9:0] _add_map_x_36_start;
  wire [9:0] _add_map_x_36_goal;
  wire [9:0] _add_map_x_36_now;
  wire [9:0] _add_map_x_36_data_out;
  wire [9:0] _add_map_x_36_data_out_index;
  wire [9:0] _add_map_x_36_data_near;
  wire _add_map_x_36_wall_t_out;
  wire [9:0] _add_map_x_36_data_org;
  wire [9:0] _add_map_x_36_data_org_near;
  wire [1:0] _add_map_x_36_s_g;
  wire [1:0] _add_map_x_36_s_g_near;
  wire _add_map_x_36_add_exe;
  wire _add_map_x_36_p_reset;
  wire _add_map_x_36_m_clock;
  wire [9:0] _add_map_x_35_moto_org_near;
  wire [9:0] _add_map_x_35_moto_org_near1;
  wire [9:0] _add_map_x_35_moto_org_near2;
  wire [9:0] _add_map_x_35_moto_org_near3;
  wire [9:0] _add_map_x_35_moto_org;
  wire [1:0] _add_map_x_35_sg_up;
  wire [1:0] _add_map_x_35_sg_down;
  wire [1:0] _add_map_x_35_sg_left;
  wire [1:0] _add_map_x_35_sg_right;
  wire _add_map_x_35_wall_t_in;
  wire [9:0] _add_map_x_35_moto;
  wire [9:0] _add_map_x_35_up;
  wire [9:0] _add_map_x_35_right;
  wire [9:0] _add_map_x_35_down;
  wire [9:0] _add_map_x_35_left;
  wire [9:0] _add_map_x_35_start;
  wire [9:0] _add_map_x_35_goal;
  wire [9:0] _add_map_x_35_now;
  wire [9:0] _add_map_x_35_data_out;
  wire [9:0] _add_map_x_35_data_out_index;
  wire [9:0] _add_map_x_35_data_near;
  wire _add_map_x_35_wall_t_out;
  wire [9:0] _add_map_x_35_data_org;
  wire [9:0] _add_map_x_35_data_org_near;
  wire [1:0] _add_map_x_35_s_g;
  wire [1:0] _add_map_x_35_s_g_near;
  wire _add_map_x_35_add_exe;
  wire _add_map_x_35_p_reset;
  wire _add_map_x_35_m_clock;
  wire [9:0] _add_map_x_34_moto_org_near;
  wire [9:0] _add_map_x_34_moto_org_near1;
  wire [9:0] _add_map_x_34_moto_org_near2;
  wire [9:0] _add_map_x_34_moto_org_near3;
  wire [9:0] _add_map_x_34_moto_org;
  wire [1:0] _add_map_x_34_sg_up;
  wire [1:0] _add_map_x_34_sg_down;
  wire [1:0] _add_map_x_34_sg_left;
  wire [1:0] _add_map_x_34_sg_right;
  wire _add_map_x_34_wall_t_in;
  wire [9:0] _add_map_x_34_moto;
  wire [9:0] _add_map_x_34_up;
  wire [9:0] _add_map_x_34_right;
  wire [9:0] _add_map_x_34_down;
  wire [9:0] _add_map_x_34_left;
  wire [9:0] _add_map_x_34_start;
  wire [9:0] _add_map_x_34_goal;
  wire [9:0] _add_map_x_34_now;
  wire [9:0] _add_map_x_34_data_out;
  wire [9:0] _add_map_x_34_data_out_index;
  wire [9:0] _add_map_x_34_data_near;
  wire _add_map_x_34_wall_t_out;
  wire [9:0] _add_map_x_34_data_org;
  wire [9:0] _add_map_x_34_data_org_near;
  wire [1:0] _add_map_x_34_s_g;
  wire [1:0] _add_map_x_34_s_g_near;
  wire _add_map_x_34_add_exe;
  wire _add_map_x_34_p_reset;
  wire _add_map_x_34_m_clock;
  wire [9:0] _add_map_x_33_moto_org_near;
  wire [9:0] _add_map_x_33_moto_org_near1;
  wire [9:0] _add_map_x_33_moto_org_near2;
  wire [9:0] _add_map_x_33_moto_org_near3;
  wire [9:0] _add_map_x_33_moto_org;
  wire [1:0] _add_map_x_33_sg_up;
  wire [1:0] _add_map_x_33_sg_down;
  wire [1:0] _add_map_x_33_sg_left;
  wire [1:0] _add_map_x_33_sg_right;
  wire _add_map_x_33_wall_t_in;
  wire [9:0] _add_map_x_33_moto;
  wire [9:0] _add_map_x_33_up;
  wire [9:0] _add_map_x_33_right;
  wire [9:0] _add_map_x_33_down;
  wire [9:0] _add_map_x_33_left;
  wire [9:0] _add_map_x_33_start;
  wire [9:0] _add_map_x_33_goal;
  wire [9:0] _add_map_x_33_now;
  wire [9:0] _add_map_x_33_data_out;
  wire [9:0] _add_map_x_33_data_out_index;
  wire [9:0] _add_map_x_33_data_near;
  wire _add_map_x_33_wall_t_out;
  wire [9:0] _add_map_x_33_data_org;
  wire [9:0] _add_map_x_33_data_org_near;
  wire [1:0] _add_map_x_33_s_g;
  wire [1:0] _add_map_x_33_s_g_near;
  wire _add_map_x_33_add_exe;
  wire _add_map_x_33_p_reset;
  wire _add_map_x_33_m_clock;
  wire [9:0] _add_map_x_32_moto_org_near;
  wire [9:0] _add_map_x_32_moto_org_near1;
  wire [9:0] _add_map_x_32_moto_org_near2;
  wire [9:0] _add_map_x_32_moto_org_near3;
  wire [9:0] _add_map_x_32_moto_org;
  wire [1:0] _add_map_x_32_sg_up;
  wire [1:0] _add_map_x_32_sg_down;
  wire [1:0] _add_map_x_32_sg_left;
  wire [1:0] _add_map_x_32_sg_right;
  wire _add_map_x_32_wall_t_in;
  wire [9:0] _add_map_x_32_moto;
  wire [9:0] _add_map_x_32_up;
  wire [9:0] _add_map_x_32_right;
  wire [9:0] _add_map_x_32_down;
  wire [9:0] _add_map_x_32_left;
  wire [9:0] _add_map_x_32_start;
  wire [9:0] _add_map_x_32_goal;
  wire [9:0] _add_map_x_32_now;
  wire [9:0] _add_map_x_32_data_out;
  wire [9:0] _add_map_x_32_data_out_index;
  wire [9:0] _add_map_x_32_data_near;
  wire _add_map_x_32_wall_t_out;
  wire [9:0] _add_map_x_32_data_org;
  wire [9:0] _add_map_x_32_data_org_near;
  wire [1:0] _add_map_x_32_s_g;
  wire [1:0] _add_map_x_32_s_g_near;
  wire _add_map_x_32_add_exe;
  wire _add_map_x_32_p_reset;
  wire _add_map_x_32_m_clock;
  wire [9:0] _add_map_x_31_moto_org_near;
  wire [9:0] _add_map_x_31_moto_org_near1;
  wire [9:0] _add_map_x_31_moto_org_near2;
  wire [9:0] _add_map_x_31_moto_org_near3;
  wire [9:0] _add_map_x_31_moto_org;
  wire [1:0] _add_map_x_31_sg_up;
  wire [1:0] _add_map_x_31_sg_down;
  wire [1:0] _add_map_x_31_sg_left;
  wire [1:0] _add_map_x_31_sg_right;
  wire _add_map_x_31_wall_t_in;
  wire [9:0] _add_map_x_31_moto;
  wire [9:0] _add_map_x_31_up;
  wire [9:0] _add_map_x_31_right;
  wire [9:0] _add_map_x_31_down;
  wire [9:0] _add_map_x_31_left;
  wire [9:0] _add_map_x_31_start;
  wire [9:0] _add_map_x_31_goal;
  wire [9:0] _add_map_x_31_now;
  wire [9:0] _add_map_x_31_data_out;
  wire [9:0] _add_map_x_31_data_out_index;
  wire [9:0] _add_map_x_31_data_near;
  wire _add_map_x_31_wall_t_out;
  wire [9:0] _add_map_x_31_data_org;
  wire [9:0] _add_map_x_31_data_org_near;
  wire [1:0] _add_map_x_31_s_g;
  wire [1:0] _add_map_x_31_s_g_near;
  wire _add_map_x_31_add_exe;
  wire _add_map_x_31_p_reset;
  wire _add_map_x_31_m_clock;
  wire [9:0] _add_map_x_30_moto_org_near;
  wire [9:0] _add_map_x_30_moto_org_near1;
  wire [9:0] _add_map_x_30_moto_org_near2;
  wire [9:0] _add_map_x_30_moto_org_near3;
  wire [9:0] _add_map_x_30_moto_org;
  wire [1:0] _add_map_x_30_sg_up;
  wire [1:0] _add_map_x_30_sg_down;
  wire [1:0] _add_map_x_30_sg_left;
  wire [1:0] _add_map_x_30_sg_right;
  wire _add_map_x_30_wall_t_in;
  wire [9:0] _add_map_x_30_moto;
  wire [9:0] _add_map_x_30_up;
  wire [9:0] _add_map_x_30_right;
  wire [9:0] _add_map_x_30_down;
  wire [9:0] _add_map_x_30_left;
  wire [9:0] _add_map_x_30_start;
  wire [9:0] _add_map_x_30_goal;
  wire [9:0] _add_map_x_30_now;
  wire [9:0] _add_map_x_30_data_out;
  wire [9:0] _add_map_x_30_data_out_index;
  wire [9:0] _add_map_x_30_data_near;
  wire _add_map_x_30_wall_t_out;
  wire [9:0] _add_map_x_30_data_org;
  wire [9:0] _add_map_x_30_data_org_near;
  wire [1:0] _add_map_x_30_s_g;
  wire [1:0] _add_map_x_30_s_g_near;
  wire _add_map_x_30_add_exe;
  wire _add_map_x_30_p_reset;
  wire _add_map_x_30_m_clock;
  wire [9:0] _add_map_x_29_moto_org_near;
  wire [9:0] _add_map_x_29_moto_org_near1;
  wire [9:0] _add_map_x_29_moto_org_near2;
  wire [9:0] _add_map_x_29_moto_org_near3;
  wire [9:0] _add_map_x_29_moto_org;
  wire [1:0] _add_map_x_29_sg_up;
  wire [1:0] _add_map_x_29_sg_down;
  wire [1:0] _add_map_x_29_sg_left;
  wire [1:0] _add_map_x_29_sg_right;
  wire _add_map_x_29_wall_t_in;
  wire [9:0] _add_map_x_29_moto;
  wire [9:0] _add_map_x_29_up;
  wire [9:0] _add_map_x_29_right;
  wire [9:0] _add_map_x_29_down;
  wire [9:0] _add_map_x_29_left;
  wire [9:0] _add_map_x_29_start;
  wire [9:0] _add_map_x_29_goal;
  wire [9:0] _add_map_x_29_now;
  wire [9:0] _add_map_x_29_data_out;
  wire [9:0] _add_map_x_29_data_out_index;
  wire [9:0] _add_map_x_29_data_near;
  wire _add_map_x_29_wall_t_out;
  wire [9:0] _add_map_x_29_data_org;
  wire [9:0] _add_map_x_29_data_org_near;
  wire [1:0] _add_map_x_29_s_g;
  wire [1:0] _add_map_x_29_s_g_near;
  wire _add_map_x_29_add_exe;
  wire _add_map_x_29_p_reset;
  wire _add_map_x_29_m_clock;
  wire [9:0] _add_map_x_28_moto_org_near;
  wire [9:0] _add_map_x_28_moto_org_near1;
  wire [9:0] _add_map_x_28_moto_org_near2;
  wire [9:0] _add_map_x_28_moto_org_near3;
  wire [9:0] _add_map_x_28_moto_org;
  wire [1:0] _add_map_x_28_sg_up;
  wire [1:0] _add_map_x_28_sg_down;
  wire [1:0] _add_map_x_28_sg_left;
  wire [1:0] _add_map_x_28_sg_right;
  wire _add_map_x_28_wall_t_in;
  wire [9:0] _add_map_x_28_moto;
  wire [9:0] _add_map_x_28_up;
  wire [9:0] _add_map_x_28_right;
  wire [9:0] _add_map_x_28_down;
  wire [9:0] _add_map_x_28_left;
  wire [9:0] _add_map_x_28_start;
  wire [9:0] _add_map_x_28_goal;
  wire [9:0] _add_map_x_28_now;
  wire [9:0] _add_map_x_28_data_out;
  wire [9:0] _add_map_x_28_data_out_index;
  wire [9:0] _add_map_x_28_data_near;
  wire _add_map_x_28_wall_t_out;
  wire [9:0] _add_map_x_28_data_org;
  wire [9:0] _add_map_x_28_data_org_near;
  wire [1:0] _add_map_x_28_s_g;
  wire [1:0] _add_map_x_28_s_g_near;
  wire _add_map_x_28_add_exe;
  wire _add_map_x_28_p_reset;
  wire _add_map_x_28_m_clock;
  wire [9:0] _add_map_x_27_moto_org_near;
  wire [9:0] _add_map_x_27_moto_org_near1;
  wire [9:0] _add_map_x_27_moto_org_near2;
  wire [9:0] _add_map_x_27_moto_org_near3;
  wire [9:0] _add_map_x_27_moto_org;
  wire [1:0] _add_map_x_27_sg_up;
  wire [1:0] _add_map_x_27_sg_down;
  wire [1:0] _add_map_x_27_sg_left;
  wire [1:0] _add_map_x_27_sg_right;
  wire _add_map_x_27_wall_t_in;
  wire [9:0] _add_map_x_27_moto;
  wire [9:0] _add_map_x_27_up;
  wire [9:0] _add_map_x_27_right;
  wire [9:0] _add_map_x_27_down;
  wire [9:0] _add_map_x_27_left;
  wire [9:0] _add_map_x_27_start;
  wire [9:0] _add_map_x_27_goal;
  wire [9:0] _add_map_x_27_now;
  wire [9:0] _add_map_x_27_data_out;
  wire [9:0] _add_map_x_27_data_out_index;
  wire [9:0] _add_map_x_27_data_near;
  wire _add_map_x_27_wall_t_out;
  wire [9:0] _add_map_x_27_data_org;
  wire [9:0] _add_map_x_27_data_org_near;
  wire [1:0] _add_map_x_27_s_g;
  wire [1:0] _add_map_x_27_s_g_near;
  wire _add_map_x_27_add_exe;
  wire _add_map_x_27_p_reset;
  wire _add_map_x_27_m_clock;
  wire [9:0] _add_map_x_26_moto_org_near;
  wire [9:0] _add_map_x_26_moto_org_near1;
  wire [9:0] _add_map_x_26_moto_org_near2;
  wire [9:0] _add_map_x_26_moto_org_near3;
  wire [9:0] _add_map_x_26_moto_org;
  wire [1:0] _add_map_x_26_sg_up;
  wire [1:0] _add_map_x_26_sg_down;
  wire [1:0] _add_map_x_26_sg_left;
  wire [1:0] _add_map_x_26_sg_right;
  wire _add_map_x_26_wall_t_in;
  wire [9:0] _add_map_x_26_moto;
  wire [9:0] _add_map_x_26_up;
  wire [9:0] _add_map_x_26_right;
  wire [9:0] _add_map_x_26_down;
  wire [9:0] _add_map_x_26_left;
  wire [9:0] _add_map_x_26_start;
  wire [9:0] _add_map_x_26_goal;
  wire [9:0] _add_map_x_26_now;
  wire [9:0] _add_map_x_26_data_out;
  wire [9:0] _add_map_x_26_data_out_index;
  wire [9:0] _add_map_x_26_data_near;
  wire _add_map_x_26_wall_t_out;
  wire [9:0] _add_map_x_26_data_org;
  wire [9:0] _add_map_x_26_data_org_near;
  wire [1:0] _add_map_x_26_s_g;
  wire [1:0] _add_map_x_26_s_g_near;
  wire _add_map_x_26_add_exe;
  wire _add_map_x_26_p_reset;
  wire _add_map_x_26_m_clock;
  wire [9:0] _add_map_x_25_moto_org_near;
  wire [9:0] _add_map_x_25_moto_org_near1;
  wire [9:0] _add_map_x_25_moto_org_near2;
  wire [9:0] _add_map_x_25_moto_org_near3;
  wire [9:0] _add_map_x_25_moto_org;
  wire [1:0] _add_map_x_25_sg_up;
  wire [1:0] _add_map_x_25_sg_down;
  wire [1:0] _add_map_x_25_sg_left;
  wire [1:0] _add_map_x_25_sg_right;
  wire _add_map_x_25_wall_t_in;
  wire [9:0] _add_map_x_25_moto;
  wire [9:0] _add_map_x_25_up;
  wire [9:0] _add_map_x_25_right;
  wire [9:0] _add_map_x_25_down;
  wire [9:0] _add_map_x_25_left;
  wire [9:0] _add_map_x_25_start;
  wire [9:0] _add_map_x_25_goal;
  wire [9:0] _add_map_x_25_now;
  wire [9:0] _add_map_x_25_data_out;
  wire [9:0] _add_map_x_25_data_out_index;
  wire [9:0] _add_map_x_25_data_near;
  wire _add_map_x_25_wall_t_out;
  wire [9:0] _add_map_x_25_data_org;
  wire [9:0] _add_map_x_25_data_org_near;
  wire [1:0] _add_map_x_25_s_g;
  wire [1:0] _add_map_x_25_s_g_near;
  wire _add_map_x_25_add_exe;
  wire _add_map_x_25_p_reset;
  wire _add_map_x_25_m_clock;
  wire [9:0] _add_map_x_24_moto_org_near;
  wire [9:0] _add_map_x_24_moto_org_near1;
  wire [9:0] _add_map_x_24_moto_org_near2;
  wire [9:0] _add_map_x_24_moto_org_near3;
  wire [9:0] _add_map_x_24_moto_org;
  wire [1:0] _add_map_x_24_sg_up;
  wire [1:0] _add_map_x_24_sg_down;
  wire [1:0] _add_map_x_24_sg_left;
  wire [1:0] _add_map_x_24_sg_right;
  wire _add_map_x_24_wall_t_in;
  wire [9:0] _add_map_x_24_moto;
  wire [9:0] _add_map_x_24_up;
  wire [9:0] _add_map_x_24_right;
  wire [9:0] _add_map_x_24_down;
  wire [9:0] _add_map_x_24_left;
  wire [9:0] _add_map_x_24_start;
  wire [9:0] _add_map_x_24_goal;
  wire [9:0] _add_map_x_24_now;
  wire [9:0] _add_map_x_24_data_out;
  wire [9:0] _add_map_x_24_data_out_index;
  wire [9:0] _add_map_x_24_data_near;
  wire _add_map_x_24_wall_t_out;
  wire [9:0] _add_map_x_24_data_org;
  wire [9:0] _add_map_x_24_data_org_near;
  wire [1:0] _add_map_x_24_s_g;
  wire [1:0] _add_map_x_24_s_g_near;
  wire _add_map_x_24_add_exe;
  wire _add_map_x_24_p_reset;
  wire _add_map_x_24_m_clock;
  wire [9:0] _add_map_x_23_moto_org_near;
  wire [9:0] _add_map_x_23_moto_org_near1;
  wire [9:0] _add_map_x_23_moto_org_near2;
  wire [9:0] _add_map_x_23_moto_org_near3;
  wire [9:0] _add_map_x_23_moto_org;
  wire [1:0] _add_map_x_23_sg_up;
  wire [1:0] _add_map_x_23_sg_down;
  wire [1:0] _add_map_x_23_sg_left;
  wire [1:0] _add_map_x_23_sg_right;
  wire _add_map_x_23_wall_t_in;
  wire [9:0] _add_map_x_23_moto;
  wire [9:0] _add_map_x_23_up;
  wire [9:0] _add_map_x_23_right;
  wire [9:0] _add_map_x_23_down;
  wire [9:0] _add_map_x_23_left;
  wire [9:0] _add_map_x_23_start;
  wire [9:0] _add_map_x_23_goal;
  wire [9:0] _add_map_x_23_now;
  wire [9:0] _add_map_x_23_data_out;
  wire [9:0] _add_map_x_23_data_out_index;
  wire [9:0] _add_map_x_23_data_near;
  wire _add_map_x_23_wall_t_out;
  wire [9:0] _add_map_x_23_data_org;
  wire [9:0] _add_map_x_23_data_org_near;
  wire [1:0] _add_map_x_23_s_g;
  wire [1:0] _add_map_x_23_s_g_near;
  wire _add_map_x_23_add_exe;
  wire _add_map_x_23_p_reset;
  wire _add_map_x_23_m_clock;
  wire [9:0] _add_map_x_22_moto_org_near;
  wire [9:0] _add_map_x_22_moto_org_near1;
  wire [9:0] _add_map_x_22_moto_org_near2;
  wire [9:0] _add_map_x_22_moto_org_near3;
  wire [9:0] _add_map_x_22_moto_org;
  wire [1:0] _add_map_x_22_sg_up;
  wire [1:0] _add_map_x_22_sg_down;
  wire [1:0] _add_map_x_22_sg_left;
  wire [1:0] _add_map_x_22_sg_right;
  wire _add_map_x_22_wall_t_in;
  wire [9:0] _add_map_x_22_moto;
  wire [9:0] _add_map_x_22_up;
  wire [9:0] _add_map_x_22_right;
  wire [9:0] _add_map_x_22_down;
  wire [9:0] _add_map_x_22_left;
  wire [9:0] _add_map_x_22_start;
  wire [9:0] _add_map_x_22_goal;
  wire [9:0] _add_map_x_22_now;
  wire [9:0] _add_map_x_22_data_out;
  wire [9:0] _add_map_x_22_data_out_index;
  wire [9:0] _add_map_x_22_data_near;
  wire _add_map_x_22_wall_t_out;
  wire [9:0] _add_map_x_22_data_org;
  wire [9:0] _add_map_x_22_data_org_near;
  wire [1:0] _add_map_x_22_s_g;
  wire [1:0] _add_map_x_22_s_g_near;
  wire _add_map_x_22_add_exe;
  wire _add_map_x_22_p_reset;
  wire _add_map_x_22_m_clock;
  wire [9:0] _add_map_x_21_moto_org_near;
  wire [9:0] _add_map_x_21_moto_org_near1;
  wire [9:0] _add_map_x_21_moto_org_near2;
  wire [9:0] _add_map_x_21_moto_org_near3;
  wire [9:0] _add_map_x_21_moto_org;
  wire [1:0] _add_map_x_21_sg_up;
  wire [1:0] _add_map_x_21_sg_down;
  wire [1:0] _add_map_x_21_sg_left;
  wire [1:0] _add_map_x_21_sg_right;
  wire _add_map_x_21_wall_t_in;
  wire [9:0] _add_map_x_21_moto;
  wire [9:0] _add_map_x_21_up;
  wire [9:0] _add_map_x_21_right;
  wire [9:0] _add_map_x_21_down;
  wire [9:0] _add_map_x_21_left;
  wire [9:0] _add_map_x_21_start;
  wire [9:0] _add_map_x_21_goal;
  wire [9:0] _add_map_x_21_now;
  wire [9:0] _add_map_x_21_data_out;
  wire [9:0] _add_map_x_21_data_out_index;
  wire [9:0] _add_map_x_21_data_near;
  wire _add_map_x_21_wall_t_out;
  wire [9:0] _add_map_x_21_data_org;
  wire [9:0] _add_map_x_21_data_org_near;
  wire [1:0] _add_map_x_21_s_g;
  wire [1:0] _add_map_x_21_s_g_near;
  wire _add_map_x_21_add_exe;
  wire _add_map_x_21_p_reset;
  wire _add_map_x_21_m_clock;
  wire [9:0] _add_map_x_20_moto_org_near;
  wire [9:0] _add_map_x_20_moto_org_near1;
  wire [9:0] _add_map_x_20_moto_org_near2;
  wire [9:0] _add_map_x_20_moto_org_near3;
  wire [9:0] _add_map_x_20_moto_org;
  wire [1:0] _add_map_x_20_sg_up;
  wire [1:0] _add_map_x_20_sg_down;
  wire [1:0] _add_map_x_20_sg_left;
  wire [1:0] _add_map_x_20_sg_right;
  wire _add_map_x_20_wall_t_in;
  wire [9:0] _add_map_x_20_moto;
  wire [9:0] _add_map_x_20_up;
  wire [9:0] _add_map_x_20_right;
  wire [9:0] _add_map_x_20_down;
  wire [9:0] _add_map_x_20_left;
  wire [9:0] _add_map_x_20_start;
  wire [9:0] _add_map_x_20_goal;
  wire [9:0] _add_map_x_20_now;
  wire [9:0] _add_map_x_20_data_out;
  wire [9:0] _add_map_x_20_data_out_index;
  wire [9:0] _add_map_x_20_data_near;
  wire _add_map_x_20_wall_t_out;
  wire [9:0] _add_map_x_20_data_org;
  wire [9:0] _add_map_x_20_data_org_near;
  wire [1:0] _add_map_x_20_s_g;
  wire [1:0] _add_map_x_20_s_g_near;
  wire _add_map_x_20_add_exe;
  wire _add_map_x_20_p_reset;
  wire _add_map_x_20_m_clock;
  wire [9:0] _add_map_x_19_moto_org_near;
  wire [9:0] _add_map_x_19_moto_org_near1;
  wire [9:0] _add_map_x_19_moto_org_near2;
  wire [9:0] _add_map_x_19_moto_org_near3;
  wire [9:0] _add_map_x_19_moto_org;
  wire [1:0] _add_map_x_19_sg_up;
  wire [1:0] _add_map_x_19_sg_down;
  wire [1:0] _add_map_x_19_sg_left;
  wire [1:0] _add_map_x_19_sg_right;
  wire _add_map_x_19_wall_t_in;
  wire [9:0] _add_map_x_19_moto;
  wire [9:0] _add_map_x_19_up;
  wire [9:0] _add_map_x_19_right;
  wire [9:0] _add_map_x_19_down;
  wire [9:0] _add_map_x_19_left;
  wire [9:0] _add_map_x_19_start;
  wire [9:0] _add_map_x_19_goal;
  wire [9:0] _add_map_x_19_now;
  wire [9:0] _add_map_x_19_data_out;
  wire [9:0] _add_map_x_19_data_out_index;
  wire [9:0] _add_map_x_19_data_near;
  wire _add_map_x_19_wall_t_out;
  wire [9:0] _add_map_x_19_data_org;
  wire [9:0] _add_map_x_19_data_org_near;
  wire [1:0] _add_map_x_19_s_g;
  wire [1:0] _add_map_x_19_s_g_near;
  wire _add_map_x_19_add_exe;
  wire _add_map_x_19_p_reset;
  wire _add_map_x_19_m_clock;
  wire [9:0] _add_map_x_18_moto_org_near;
  wire [9:0] _add_map_x_18_moto_org_near1;
  wire [9:0] _add_map_x_18_moto_org_near2;
  wire [9:0] _add_map_x_18_moto_org_near3;
  wire [9:0] _add_map_x_18_moto_org;
  wire [1:0] _add_map_x_18_sg_up;
  wire [1:0] _add_map_x_18_sg_down;
  wire [1:0] _add_map_x_18_sg_left;
  wire [1:0] _add_map_x_18_sg_right;
  wire _add_map_x_18_wall_t_in;
  wire [9:0] _add_map_x_18_moto;
  wire [9:0] _add_map_x_18_up;
  wire [9:0] _add_map_x_18_right;
  wire [9:0] _add_map_x_18_down;
  wire [9:0] _add_map_x_18_left;
  wire [9:0] _add_map_x_18_start;
  wire [9:0] _add_map_x_18_goal;
  wire [9:0] _add_map_x_18_now;
  wire [9:0] _add_map_x_18_data_out;
  wire [9:0] _add_map_x_18_data_out_index;
  wire [9:0] _add_map_x_18_data_near;
  wire _add_map_x_18_wall_t_out;
  wire [9:0] _add_map_x_18_data_org;
  wire [9:0] _add_map_x_18_data_org_near;
  wire [1:0] _add_map_x_18_s_g;
  wire [1:0] _add_map_x_18_s_g_near;
  wire _add_map_x_18_add_exe;
  wire _add_map_x_18_p_reset;
  wire _add_map_x_18_m_clock;
  wire [9:0] _add_map_x_17_moto_org_near;
  wire [9:0] _add_map_x_17_moto_org_near1;
  wire [9:0] _add_map_x_17_moto_org_near2;
  wire [9:0] _add_map_x_17_moto_org_near3;
  wire [9:0] _add_map_x_17_moto_org;
  wire [1:0] _add_map_x_17_sg_up;
  wire [1:0] _add_map_x_17_sg_down;
  wire [1:0] _add_map_x_17_sg_left;
  wire [1:0] _add_map_x_17_sg_right;
  wire _add_map_x_17_wall_t_in;
  wire [9:0] _add_map_x_17_moto;
  wire [9:0] _add_map_x_17_up;
  wire [9:0] _add_map_x_17_right;
  wire [9:0] _add_map_x_17_down;
  wire [9:0] _add_map_x_17_left;
  wire [9:0] _add_map_x_17_start;
  wire [9:0] _add_map_x_17_goal;
  wire [9:0] _add_map_x_17_now;
  wire [9:0] _add_map_x_17_data_out;
  wire [9:0] _add_map_x_17_data_out_index;
  wire [9:0] _add_map_x_17_data_near;
  wire _add_map_x_17_wall_t_out;
  wire [9:0] _add_map_x_17_data_org;
  wire [9:0] _add_map_x_17_data_org_near;
  wire [1:0] _add_map_x_17_s_g;
  wire [1:0] _add_map_x_17_s_g_near;
  wire _add_map_x_17_add_exe;
  wire _add_map_x_17_p_reset;
  wire _add_map_x_17_m_clock;
  wire [9:0] _add_map_x_16_moto_org_near;
  wire [9:0] _add_map_x_16_moto_org_near1;
  wire [9:0] _add_map_x_16_moto_org_near2;
  wire [9:0] _add_map_x_16_moto_org_near3;
  wire [9:0] _add_map_x_16_moto_org;
  wire [1:0] _add_map_x_16_sg_up;
  wire [1:0] _add_map_x_16_sg_down;
  wire [1:0] _add_map_x_16_sg_left;
  wire [1:0] _add_map_x_16_sg_right;
  wire _add_map_x_16_wall_t_in;
  wire [9:0] _add_map_x_16_moto;
  wire [9:0] _add_map_x_16_up;
  wire [9:0] _add_map_x_16_right;
  wire [9:0] _add_map_x_16_down;
  wire [9:0] _add_map_x_16_left;
  wire [9:0] _add_map_x_16_start;
  wire [9:0] _add_map_x_16_goal;
  wire [9:0] _add_map_x_16_now;
  wire [9:0] _add_map_x_16_data_out;
  wire [9:0] _add_map_x_16_data_out_index;
  wire [9:0] _add_map_x_16_data_near;
  wire _add_map_x_16_wall_t_out;
  wire [9:0] _add_map_x_16_data_org;
  wire [9:0] _add_map_x_16_data_org_near;
  wire [1:0] _add_map_x_16_s_g;
  wire [1:0] _add_map_x_16_s_g_near;
  wire _add_map_x_16_add_exe;
  wire _add_map_x_16_p_reset;
  wire _add_map_x_16_m_clock;
  wire [9:0] _add_map_x_15_moto_org_near;
  wire [9:0] _add_map_x_15_moto_org_near1;
  wire [9:0] _add_map_x_15_moto_org_near2;
  wire [9:0] _add_map_x_15_moto_org_near3;
  wire [9:0] _add_map_x_15_moto_org;
  wire [1:0] _add_map_x_15_sg_up;
  wire [1:0] _add_map_x_15_sg_down;
  wire [1:0] _add_map_x_15_sg_left;
  wire [1:0] _add_map_x_15_sg_right;
  wire _add_map_x_15_wall_t_in;
  wire [9:0] _add_map_x_15_moto;
  wire [9:0] _add_map_x_15_up;
  wire [9:0] _add_map_x_15_right;
  wire [9:0] _add_map_x_15_down;
  wire [9:0] _add_map_x_15_left;
  wire [9:0] _add_map_x_15_start;
  wire [9:0] _add_map_x_15_goal;
  wire [9:0] _add_map_x_15_now;
  wire [9:0] _add_map_x_15_data_out;
  wire [9:0] _add_map_x_15_data_out_index;
  wire [9:0] _add_map_x_15_data_near;
  wire _add_map_x_15_wall_t_out;
  wire [9:0] _add_map_x_15_data_org;
  wire [9:0] _add_map_x_15_data_org_near;
  wire [1:0] _add_map_x_15_s_g;
  wire [1:0] _add_map_x_15_s_g_near;
  wire _add_map_x_15_add_exe;
  wire _add_map_x_15_p_reset;
  wire _add_map_x_15_m_clock;
  wire [9:0] _add_map_x_14_moto_org_near;
  wire [9:0] _add_map_x_14_moto_org_near1;
  wire [9:0] _add_map_x_14_moto_org_near2;
  wire [9:0] _add_map_x_14_moto_org_near3;
  wire [9:0] _add_map_x_14_moto_org;
  wire [1:0] _add_map_x_14_sg_up;
  wire [1:0] _add_map_x_14_sg_down;
  wire [1:0] _add_map_x_14_sg_left;
  wire [1:0] _add_map_x_14_sg_right;
  wire _add_map_x_14_wall_t_in;
  wire [9:0] _add_map_x_14_moto;
  wire [9:0] _add_map_x_14_up;
  wire [9:0] _add_map_x_14_right;
  wire [9:0] _add_map_x_14_down;
  wire [9:0] _add_map_x_14_left;
  wire [9:0] _add_map_x_14_start;
  wire [9:0] _add_map_x_14_goal;
  wire [9:0] _add_map_x_14_now;
  wire [9:0] _add_map_x_14_data_out;
  wire [9:0] _add_map_x_14_data_out_index;
  wire [9:0] _add_map_x_14_data_near;
  wire _add_map_x_14_wall_t_out;
  wire [9:0] _add_map_x_14_data_org;
  wire [9:0] _add_map_x_14_data_org_near;
  wire [1:0] _add_map_x_14_s_g;
  wire [1:0] _add_map_x_14_s_g_near;
  wire _add_map_x_14_add_exe;
  wire _add_map_x_14_p_reset;
  wire _add_map_x_14_m_clock;
  wire [9:0] _add_map_x_13_moto_org_near;
  wire [9:0] _add_map_x_13_moto_org_near1;
  wire [9:0] _add_map_x_13_moto_org_near2;
  wire [9:0] _add_map_x_13_moto_org_near3;
  wire [9:0] _add_map_x_13_moto_org;
  wire [1:0] _add_map_x_13_sg_up;
  wire [1:0] _add_map_x_13_sg_down;
  wire [1:0] _add_map_x_13_sg_left;
  wire [1:0] _add_map_x_13_sg_right;
  wire _add_map_x_13_wall_t_in;
  wire [9:0] _add_map_x_13_moto;
  wire [9:0] _add_map_x_13_up;
  wire [9:0] _add_map_x_13_right;
  wire [9:0] _add_map_x_13_down;
  wire [9:0] _add_map_x_13_left;
  wire [9:0] _add_map_x_13_start;
  wire [9:0] _add_map_x_13_goal;
  wire [9:0] _add_map_x_13_now;
  wire [9:0] _add_map_x_13_data_out;
  wire [9:0] _add_map_x_13_data_out_index;
  wire [9:0] _add_map_x_13_data_near;
  wire _add_map_x_13_wall_t_out;
  wire [9:0] _add_map_x_13_data_org;
  wire [9:0] _add_map_x_13_data_org_near;
  wire [1:0] _add_map_x_13_s_g;
  wire [1:0] _add_map_x_13_s_g_near;
  wire _add_map_x_13_add_exe;
  wire _add_map_x_13_p_reset;
  wire _add_map_x_13_m_clock;
  wire [9:0] _add_map_x_12_moto_org_near;
  wire [9:0] _add_map_x_12_moto_org_near1;
  wire [9:0] _add_map_x_12_moto_org_near2;
  wire [9:0] _add_map_x_12_moto_org_near3;
  wire [9:0] _add_map_x_12_moto_org;
  wire [1:0] _add_map_x_12_sg_up;
  wire [1:0] _add_map_x_12_sg_down;
  wire [1:0] _add_map_x_12_sg_left;
  wire [1:0] _add_map_x_12_sg_right;
  wire _add_map_x_12_wall_t_in;
  wire [9:0] _add_map_x_12_moto;
  wire [9:0] _add_map_x_12_up;
  wire [9:0] _add_map_x_12_right;
  wire [9:0] _add_map_x_12_down;
  wire [9:0] _add_map_x_12_left;
  wire [9:0] _add_map_x_12_start;
  wire [9:0] _add_map_x_12_goal;
  wire [9:0] _add_map_x_12_now;
  wire [9:0] _add_map_x_12_data_out;
  wire [9:0] _add_map_x_12_data_out_index;
  wire [9:0] _add_map_x_12_data_near;
  wire _add_map_x_12_wall_t_out;
  wire [9:0] _add_map_x_12_data_org;
  wire [9:0] _add_map_x_12_data_org_near;
  wire [1:0] _add_map_x_12_s_g;
  wire [1:0] _add_map_x_12_s_g_near;
  wire _add_map_x_12_add_exe;
  wire _add_map_x_12_p_reset;
  wire _add_map_x_12_m_clock;
  wire [9:0] _add_map_x_11_moto_org_near;
  wire [9:0] _add_map_x_11_moto_org_near1;
  wire [9:0] _add_map_x_11_moto_org_near2;
  wire [9:0] _add_map_x_11_moto_org_near3;
  wire [9:0] _add_map_x_11_moto_org;
  wire [1:0] _add_map_x_11_sg_up;
  wire [1:0] _add_map_x_11_sg_down;
  wire [1:0] _add_map_x_11_sg_left;
  wire [1:0] _add_map_x_11_sg_right;
  wire _add_map_x_11_wall_t_in;
  wire [9:0] _add_map_x_11_moto;
  wire [9:0] _add_map_x_11_up;
  wire [9:0] _add_map_x_11_right;
  wire [9:0] _add_map_x_11_down;
  wire [9:0] _add_map_x_11_left;
  wire [9:0] _add_map_x_11_start;
  wire [9:0] _add_map_x_11_goal;
  wire [9:0] _add_map_x_11_now;
  wire [9:0] _add_map_x_11_data_out;
  wire [9:0] _add_map_x_11_data_out_index;
  wire [9:0] _add_map_x_11_data_near;
  wire _add_map_x_11_wall_t_out;
  wire [9:0] _add_map_x_11_data_org;
  wire [9:0] _add_map_x_11_data_org_near;
  wire [1:0] _add_map_x_11_s_g;
  wire [1:0] _add_map_x_11_s_g_near;
  wire _add_map_x_11_add_exe;
  wire _add_map_x_11_p_reset;
  wire _add_map_x_11_m_clock;
  wire [9:0] _add_map_x_10_moto_org_near;
  wire [9:0] _add_map_x_10_moto_org_near1;
  wire [9:0] _add_map_x_10_moto_org_near2;
  wire [9:0] _add_map_x_10_moto_org_near3;
  wire [9:0] _add_map_x_10_moto_org;
  wire [1:0] _add_map_x_10_sg_up;
  wire [1:0] _add_map_x_10_sg_down;
  wire [1:0] _add_map_x_10_sg_left;
  wire [1:0] _add_map_x_10_sg_right;
  wire _add_map_x_10_wall_t_in;
  wire [9:0] _add_map_x_10_moto;
  wire [9:0] _add_map_x_10_up;
  wire [9:0] _add_map_x_10_right;
  wire [9:0] _add_map_x_10_down;
  wire [9:0] _add_map_x_10_left;
  wire [9:0] _add_map_x_10_start;
  wire [9:0] _add_map_x_10_goal;
  wire [9:0] _add_map_x_10_now;
  wire [9:0] _add_map_x_10_data_out;
  wire [9:0] _add_map_x_10_data_out_index;
  wire [9:0] _add_map_x_10_data_near;
  wire _add_map_x_10_wall_t_out;
  wire [9:0] _add_map_x_10_data_org;
  wire [9:0] _add_map_x_10_data_org_near;
  wire [1:0] _add_map_x_10_s_g;
  wire [1:0] _add_map_x_10_s_g_near;
  wire _add_map_x_10_add_exe;
  wire _add_map_x_10_p_reset;
  wire _add_map_x_10_m_clock;
  wire [9:0] _add_map_x_9_moto_org_near;
  wire [9:0] _add_map_x_9_moto_org_near1;
  wire [9:0] _add_map_x_9_moto_org_near2;
  wire [9:0] _add_map_x_9_moto_org_near3;
  wire [9:0] _add_map_x_9_moto_org;
  wire [1:0] _add_map_x_9_sg_up;
  wire [1:0] _add_map_x_9_sg_down;
  wire [1:0] _add_map_x_9_sg_left;
  wire [1:0] _add_map_x_9_sg_right;
  wire _add_map_x_9_wall_t_in;
  wire [9:0] _add_map_x_9_moto;
  wire [9:0] _add_map_x_9_up;
  wire [9:0] _add_map_x_9_right;
  wire [9:0] _add_map_x_9_down;
  wire [9:0] _add_map_x_9_left;
  wire [9:0] _add_map_x_9_start;
  wire [9:0] _add_map_x_9_goal;
  wire [9:0] _add_map_x_9_now;
  wire [9:0] _add_map_x_9_data_out;
  wire [9:0] _add_map_x_9_data_out_index;
  wire [9:0] _add_map_x_9_data_near;
  wire _add_map_x_9_wall_t_out;
  wire [9:0] _add_map_x_9_data_org;
  wire [9:0] _add_map_x_9_data_org_near;
  wire [1:0] _add_map_x_9_s_g;
  wire [1:0] _add_map_x_9_s_g_near;
  wire _add_map_x_9_add_exe;
  wire _add_map_x_9_p_reset;
  wire _add_map_x_9_m_clock;
  wire [9:0] _add_map_x_8_moto_org_near;
  wire [9:0] _add_map_x_8_moto_org_near1;
  wire [9:0] _add_map_x_8_moto_org_near2;
  wire [9:0] _add_map_x_8_moto_org_near3;
  wire [9:0] _add_map_x_8_moto_org;
  wire [1:0] _add_map_x_8_sg_up;
  wire [1:0] _add_map_x_8_sg_down;
  wire [1:0] _add_map_x_8_sg_left;
  wire [1:0] _add_map_x_8_sg_right;
  wire _add_map_x_8_wall_t_in;
  wire [9:0] _add_map_x_8_moto;
  wire [9:0] _add_map_x_8_up;
  wire [9:0] _add_map_x_8_right;
  wire [9:0] _add_map_x_8_down;
  wire [9:0] _add_map_x_8_left;
  wire [9:0] _add_map_x_8_start;
  wire [9:0] _add_map_x_8_goal;
  wire [9:0] _add_map_x_8_now;
  wire [9:0] _add_map_x_8_data_out;
  wire [9:0] _add_map_x_8_data_out_index;
  wire [9:0] _add_map_x_8_data_near;
  wire _add_map_x_8_wall_t_out;
  wire [9:0] _add_map_x_8_data_org;
  wire [9:0] _add_map_x_8_data_org_near;
  wire [1:0] _add_map_x_8_s_g;
  wire [1:0] _add_map_x_8_s_g_near;
  wire _add_map_x_8_add_exe;
  wire _add_map_x_8_p_reset;
  wire _add_map_x_8_m_clock;
  wire [9:0] _add_map_x_7_moto_org_near;
  wire [9:0] _add_map_x_7_moto_org_near1;
  wire [9:0] _add_map_x_7_moto_org_near2;
  wire [9:0] _add_map_x_7_moto_org_near3;
  wire [9:0] _add_map_x_7_moto_org;
  wire [1:0] _add_map_x_7_sg_up;
  wire [1:0] _add_map_x_7_sg_down;
  wire [1:0] _add_map_x_7_sg_left;
  wire [1:0] _add_map_x_7_sg_right;
  wire _add_map_x_7_wall_t_in;
  wire [9:0] _add_map_x_7_moto;
  wire [9:0] _add_map_x_7_up;
  wire [9:0] _add_map_x_7_right;
  wire [9:0] _add_map_x_7_down;
  wire [9:0] _add_map_x_7_left;
  wire [9:0] _add_map_x_7_start;
  wire [9:0] _add_map_x_7_goal;
  wire [9:0] _add_map_x_7_now;
  wire [9:0] _add_map_x_7_data_out;
  wire [9:0] _add_map_x_7_data_out_index;
  wire [9:0] _add_map_x_7_data_near;
  wire _add_map_x_7_wall_t_out;
  wire [9:0] _add_map_x_7_data_org;
  wire [9:0] _add_map_x_7_data_org_near;
  wire [1:0] _add_map_x_7_s_g;
  wire [1:0] _add_map_x_7_s_g_near;
  wire _add_map_x_7_add_exe;
  wire _add_map_x_7_p_reset;
  wire _add_map_x_7_m_clock;
  wire [9:0] _add_map_x_6_moto_org_near;
  wire [9:0] _add_map_x_6_moto_org_near1;
  wire [9:0] _add_map_x_6_moto_org_near2;
  wire [9:0] _add_map_x_6_moto_org_near3;
  wire [9:0] _add_map_x_6_moto_org;
  wire [1:0] _add_map_x_6_sg_up;
  wire [1:0] _add_map_x_6_sg_down;
  wire [1:0] _add_map_x_6_sg_left;
  wire [1:0] _add_map_x_6_sg_right;
  wire _add_map_x_6_wall_t_in;
  wire [9:0] _add_map_x_6_moto;
  wire [9:0] _add_map_x_6_up;
  wire [9:0] _add_map_x_6_right;
  wire [9:0] _add_map_x_6_down;
  wire [9:0] _add_map_x_6_left;
  wire [9:0] _add_map_x_6_start;
  wire [9:0] _add_map_x_6_goal;
  wire [9:0] _add_map_x_6_now;
  wire [9:0] _add_map_x_6_data_out;
  wire [9:0] _add_map_x_6_data_out_index;
  wire [9:0] _add_map_x_6_data_near;
  wire _add_map_x_6_wall_t_out;
  wire [9:0] _add_map_x_6_data_org;
  wire [9:0] _add_map_x_6_data_org_near;
  wire [1:0] _add_map_x_6_s_g;
  wire [1:0] _add_map_x_6_s_g_near;
  wire _add_map_x_6_add_exe;
  wire _add_map_x_6_p_reset;
  wire _add_map_x_6_m_clock;
  wire [9:0] _add_map_x_5_moto_org_near;
  wire [9:0] _add_map_x_5_moto_org_near1;
  wire [9:0] _add_map_x_5_moto_org_near2;
  wire [9:0] _add_map_x_5_moto_org_near3;
  wire [9:0] _add_map_x_5_moto_org;
  wire [1:0] _add_map_x_5_sg_up;
  wire [1:0] _add_map_x_5_sg_down;
  wire [1:0] _add_map_x_5_sg_left;
  wire [1:0] _add_map_x_5_sg_right;
  wire _add_map_x_5_wall_t_in;
  wire [9:0] _add_map_x_5_moto;
  wire [9:0] _add_map_x_5_up;
  wire [9:0] _add_map_x_5_right;
  wire [9:0] _add_map_x_5_down;
  wire [9:0] _add_map_x_5_left;
  wire [9:0] _add_map_x_5_start;
  wire [9:0] _add_map_x_5_goal;
  wire [9:0] _add_map_x_5_now;
  wire [9:0] _add_map_x_5_data_out;
  wire [9:0] _add_map_x_5_data_out_index;
  wire [9:0] _add_map_x_5_data_near;
  wire _add_map_x_5_wall_t_out;
  wire [9:0] _add_map_x_5_data_org;
  wire [9:0] _add_map_x_5_data_org_near;
  wire [1:0] _add_map_x_5_s_g;
  wire [1:0] _add_map_x_5_s_g_near;
  wire _add_map_x_5_add_exe;
  wire _add_map_x_5_p_reset;
  wire _add_map_x_5_m_clock;
  wire [9:0] _add_map_x_4_moto_org_near;
  wire [9:0] _add_map_x_4_moto_org_near1;
  wire [9:0] _add_map_x_4_moto_org_near2;
  wire [9:0] _add_map_x_4_moto_org_near3;
  wire [9:0] _add_map_x_4_moto_org;
  wire [1:0] _add_map_x_4_sg_up;
  wire [1:0] _add_map_x_4_sg_down;
  wire [1:0] _add_map_x_4_sg_left;
  wire [1:0] _add_map_x_4_sg_right;
  wire _add_map_x_4_wall_t_in;
  wire [9:0] _add_map_x_4_moto;
  wire [9:0] _add_map_x_4_up;
  wire [9:0] _add_map_x_4_right;
  wire [9:0] _add_map_x_4_down;
  wire [9:0] _add_map_x_4_left;
  wire [9:0] _add_map_x_4_start;
  wire [9:0] _add_map_x_4_goal;
  wire [9:0] _add_map_x_4_now;
  wire [9:0] _add_map_x_4_data_out;
  wire [9:0] _add_map_x_4_data_out_index;
  wire [9:0] _add_map_x_4_data_near;
  wire _add_map_x_4_wall_t_out;
  wire [9:0] _add_map_x_4_data_org;
  wire [9:0] _add_map_x_4_data_org_near;
  wire [1:0] _add_map_x_4_s_g;
  wire [1:0] _add_map_x_4_s_g_near;
  wire _add_map_x_4_add_exe;
  wire _add_map_x_4_p_reset;
  wire _add_map_x_4_m_clock;
  wire [9:0] _add_map_x_3_moto_org_near;
  wire [9:0] _add_map_x_3_moto_org_near1;
  wire [9:0] _add_map_x_3_moto_org_near2;
  wire [9:0] _add_map_x_3_moto_org_near3;
  wire [9:0] _add_map_x_3_moto_org;
  wire [1:0] _add_map_x_3_sg_up;
  wire [1:0] _add_map_x_3_sg_down;
  wire [1:0] _add_map_x_3_sg_left;
  wire [1:0] _add_map_x_3_sg_right;
  wire _add_map_x_3_wall_t_in;
  wire [9:0] _add_map_x_3_moto;
  wire [9:0] _add_map_x_3_up;
  wire [9:0] _add_map_x_3_right;
  wire [9:0] _add_map_x_3_down;
  wire [9:0] _add_map_x_3_left;
  wire [9:0] _add_map_x_3_start;
  wire [9:0] _add_map_x_3_goal;
  wire [9:0] _add_map_x_3_now;
  wire [9:0] _add_map_x_3_data_out;
  wire [9:0] _add_map_x_3_data_out_index;
  wire [9:0] _add_map_x_3_data_near;
  wire _add_map_x_3_wall_t_out;
  wire [9:0] _add_map_x_3_data_org;
  wire [9:0] _add_map_x_3_data_org_near;
  wire [1:0] _add_map_x_3_s_g;
  wire [1:0] _add_map_x_3_s_g_near;
  wire _add_map_x_3_add_exe;
  wire _add_map_x_3_p_reset;
  wire _add_map_x_3_m_clock;
  wire [9:0] _add_map_x_2_moto_org_near;
  wire [9:0] _add_map_x_2_moto_org_near1;
  wire [9:0] _add_map_x_2_moto_org_near2;
  wire [9:0] _add_map_x_2_moto_org_near3;
  wire [9:0] _add_map_x_2_moto_org;
  wire [1:0] _add_map_x_2_sg_up;
  wire [1:0] _add_map_x_2_sg_down;
  wire [1:0] _add_map_x_2_sg_left;
  wire [1:0] _add_map_x_2_sg_right;
  wire _add_map_x_2_wall_t_in;
  wire [9:0] _add_map_x_2_moto;
  wire [9:0] _add_map_x_2_up;
  wire [9:0] _add_map_x_2_right;
  wire [9:0] _add_map_x_2_down;
  wire [9:0] _add_map_x_2_left;
  wire [9:0] _add_map_x_2_start;
  wire [9:0] _add_map_x_2_goal;
  wire [9:0] _add_map_x_2_now;
  wire [9:0] _add_map_x_2_data_out;
  wire [9:0] _add_map_x_2_data_out_index;
  wire [9:0] _add_map_x_2_data_near;
  wire _add_map_x_2_wall_t_out;
  wire [9:0] _add_map_x_2_data_org;
  wire [9:0] _add_map_x_2_data_org_near;
  wire [1:0] _add_map_x_2_s_g;
  wire [1:0] _add_map_x_2_s_g_near;
  wire _add_map_x_2_add_exe;
  wire _add_map_x_2_p_reset;
  wire _add_map_x_2_m_clock;
  wire [9:0] _add_map_x_1_moto_org_near;
  wire [9:0] _add_map_x_1_moto_org_near1;
  wire [9:0] _add_map_x_1_moto_org_near2;
  wire [9:0] _add_map_x_1_moto_org_near3;
  wire [9:0] _add_map_x_1_moto_org;
  wire [1:0] _add_map_x_1_sg_up;
  wire [1:0] _add_map_x_1_sg_down;
  wire [1:0] _add_map_x_1_sg_left;
  wire [1:0] _add_map_x_1_sg_right;
  wire _add_map_x_1_wall_t_in;
  wire [9:0] _add_map_x_1_moto;
  wire [9:0] _add_map_x_1_up;
  wire [9:0] _add_map_x_1_right;
  wire [9:0] _add_map_x_1_down;
  wire [9:0] _add_map_x_1_left;
  wire [9:0] _add_map_x_1_start;
  wire [9:0] _add_map_x_1_goal;
  wire [9:0] _add_map_x_1_now;
  wire [9:0] _add_map_x_1_data_out;
  wire [9:0] _add_map_x_1_data_out_index;
  wire [9:0] _add_map_x_1_data_near;
  wire _add_map_x_1_wall_t_out;
  wire [9:0] _add_map_x_1_data_org;
  wire [9:0] _add_map_x_1_data_org_near;
  wire [1:0] _add_map_x_1_s_g;
  wire [1:0] _add_map_x_1_s_g_near;
  wire _add_map_x_1_add_exe;
  wire _add_map_x_1_p_reset;
  wire _add_map_x_1_m_clock;
  wire _net_0;
  wire _net_1;
  wire _net_2;
  wire _net_3;
  wire _net_4;
  wire _net_5;
  wire _net_6;
  wire _net_7;
  wire _net_8;
  wire _net_9;
  wire _net_10;
  wire _net_11;
  wire _net_12;
  wire _net_13;
  wire _net_14;
  wire _net_15;
  wire _net_16;
  wire _net_17;
  wire _net_18;
  wire _net_19;
  wire _net_20;
  wire _net_21;
  wire _net_22;
  wire _net_23;
  wire _net_24;
  wire _net_25;
  wire _net_26;
  wire _net_27;
  wire _net_28;
  wire _net_29;
  wire _net_30;
  wire _net_31;
  wire _net_32;
  wire _net_33;
  wire _net_34;
  wire _net_35;
  wire _net_36;
  wire _net_37;
  wire _net_38;
  wire _net_39;
  wire _net_40;
  wire _net_41;
  wire _net_42;
  wire _net_43;
  wire _net_44;
  wire _net_45;
  wire _net_46;
  wire _net_47;
  wire _net_48;
  wire _net_49;
  wire _net_50;
  wire _net_51;
  wire _net_52;
  wire _net_53;
  wire _net_54;
  wire _net_55;
  wire _net_56;
  wire _net_57;
  wire _net_58;
  wire _net_59;
  wire _net_60;
  wire _net_61;
  wire _net_62;
  wire _net_63;
  wire _net_64;
  wire _net_65;
  wire _net_66;
  wire _net_67;
  wire _net_68;
  wire _net_69;
  wire _net_70;
  wire _net_71;
  wire _net_72;
  wire _net_73;
  wire _net_74;
  wire _net_75;
  wire _net_76;
  wire _net_77;
  wire _net_78;
  wire _net_79;
  wire _net_80;
  wire _net_81;
  wire _net_82;
  wire _net_83;
  wire _net_84;
  wire _net_85;
  wire _net_86;
  wire _net_87;
  wire _net_88;
  wire _net_89;
  wire _net_90;
  wire _net_91;
  wire _net_92;
  wire _net_93;
  wire _net_94;
  wire _net_95;
  wire _net_96;
  wire _net_97;
  wire _net_98;
  wire _net_99;
  wire _net_100;
  wire _net_101;
  wire _net_102;
  wire _net_103;
  wire _net_104;
  wire _net_105;
  wire _net_106;
  wire _net_107;
  wire _net_108;
  wire _net_109;
  wire _net_110;
  wire _net_111;
  wire _net_112;
  wire _net_113;
  wire _net_114;
  wire _net_115;
  wire _net_116;
  wire _net_117;
  wire _net_118;
  wire _net_119;
  wire _net_120;
  wire _net_121;
  wire _net_122;
  wire _net_123;
  wire _net_124;
  wire _net_125;
  wire _net_126;
  wire _net_127;
  wire _net_128;
  wire _net_129;
  wire _net_130;
  wire _net_131;
  wire _net_132;
  wire _net_133;
  wire _net_134;
  wire _net_135;
  wire _net_136;
  wire _net_137;
  wire _net_138;
  wire _net_139;
  wire _net_140;
  wire _net_141;
  wire _net_142;
  wire _net_143;
  wire _net_144;
  wire _net_145;
  wire _net_146;
  wire _net_147;
  wire _net_148;
  wire _net_149;
  wire _net_150;
  wire _net_151;
  wire _net_152;
  wire _net_153;
  wire _net_154;
  wire _net_155;
  wire _net_156;
  wire _net_157;
  wire _net_158;
  wire _net_159;
  wire _net_160;
  wire _net_161;
  wire _net_162;
  wire _net_163;
  wire _net_164;
  wire _net_165;
  wire _net_166;
  wire _net_167;
  wire _net_168;
  wire _net_169;
  wire _net_170;
  wire _net_171;
  wire _net_172;
  wire _net_173;
  wire _net_174;
  wire _net_175;
  wire _net_176;
  wire _net_177;
  wire _net_178;
  wire _net_179;
  wire _net_180;
  wire _net_181;
  wire _net_182;
  wire _net_183;
  wire _net_184;
  wire _net_185;
  wire _net_186;
  wire _net_187;
  wire _net_188;
  wire _net_189;
  wire _net_190;
  wire _net_191;
  wire _net_192;
  wire _net_193;
  wire _net_194;
  wire _net_195;
  wire _net_196;
  wire _net_197;
  wire _net_198;
  wire _net_199;
  wire _net_200;
  wire _net_201;
  wire _net_202;
  wire _net_203;
  wire _net_204;
  wire _net_205;
  wire _net_206;
  wire _net_207;
  wire _net_208;
  wire _net_209;
  wire _net_210;
  wire _net_211;
  wire _net_212;
  wire _net_213;
  wire _net_214;
  wire _net_215;
  wire _net_216;
  wire _net_217;
  wire _net_218;
  wire _net_219;
  wire _net_220;
  wire _net_221;
  wire _net_222;
  wire _net_223;
  wire _net_224;
  wire _net_225;
  wire _net_226;
  wire _net_227;
  wire _net_228;
  wire _net_229;
  wire _net_230;
  wire _net_231;
  wire _net_232;
  wire _net_233;
  wire _net_234;
  wire _net_235;
  wire _net_236;
  wire _net_237;
  wire _net_238;
  wire _net_239;
  wire _net_240;
  wire _net_241;
  wire _net_242;
  wire _net_243;
  wire _net_244;
  wire _net_245;
  wire _net_246;
  wire _net_247;
  wire _net_248;
  wire _net_249;
  wire _net_250;
  wire _net_251;
  wire _net_252;
  wire _net_253;
  wire _net_254;
  wire _net_255;
  wire _net_256;
  wire _net_257;
  wire _net_258;
  wire _net_259;
  wire _net_260;
  wire _net_261;
  wire _net_262;
  wire _net_263;
  wire _net_264;
  wire _net_265;
  wire _net_266;
  wire _net_267;
  wire _net_268;
  wire _net_269;
  wire _net_270;
  wire _net_271;
  wire _net_272;
  wire _net_273;
  wire _net_274;
  wire _net_275;
  wire _net_276;
  wire _net_277;
  wire _net_278;
  wire _net_279;
  wire _net_280;
  wire _net_281;
  wire _net_282;
  wire _net_283;
  wire _net_284;
  wire _net_285;
  wire _net_286;
  wire _net_287;
  wire _net_288;
  wire _net_289;
  wire _net_290;
  wire _net_291;
  wire _net_292;
  wire _net_293;
  wire _net_294;
  wire _net_295;
  wire _net_296;
  wire _net_297;
  wire _net_298;
  wire _net_299;
  wire _net_300;
  wire _net_301;
  wire _net_302;
  wire _net_303;
  wire _net_304;
  wire _net_305;
  wire _net_306;
  wire _net_307;
  wire _net_308;
  wire _net_309;
  wire _net_310;
  wire _net_311;
  wire _net_312;
  wire _net_313;
  wire _net_314;
  wire _net_315;
  wire _net_316;
  wire _net_317;
  wire _net_318;
  wire _net_319;
  wire _net_320;
  wire _net_321;
  wire _net_322;
  wire _net_323;
  wire _net_324;
  wire _net_325;
  wire _net_326;
  wire _net_327;
  wire _net_328;
  wire _net_329;
  wire _net_330;
  wire _net_331;
  wire _net_332;
  wire _net_333;
  wire _net_334;
  wire _net_335;
  wire _net_336;
  wire _net_337;
  wire _net_338;
  wire _net_339;
  wire _net_340;
  wire _net_341;
  wire _net_342;
  wire _net_343;
  wire _net_344;
  wire _net_345;
  wire _net_346;
  wire _net_347;
  wire _net_348;
  wire _net_349;
  wire _net_350;
  wire _net_351;
  wire _net_352;
  wire _net_353;
  wire _net_354;
  wire _net_355;
  wire _net_356;
  wire _net_357;
  wire _net_358;
  wire _net_359;
  wire _net_360;
  wire _net_361;
  wire _net_362;
  wire _net_363;
  wire _net_364;
  wire _net_365;
  wire _net_366;
  wire _net_367;
  wire _net_368;
  wire _net_369;
  wire _net_370;
  wire _net_371;
  wire _net_372;
  wire _net_373;
  wire _net_374;
  wire _net_375;
  wire _net_376;
  wire _net_377;
  wire _net_378;
  wire _net_379;
  wire _net_380;
  wire _net_381;
  wire _net_382;
  wire _net_383;
  wire _net_384;
  wire _net_385;
  wire _net_386;
  wire _net_387;
  wire _net_388;
  wire _net_389;
  wire _net_390;
  wire _net_391;
  wire _net_392;
  wire _net_393;
  wire _net_394;
  wire _net_395;
  wire _net_396;
  wire _net_397;
  wire _net_398;
  wire _net_399;
  wire _net_400;
  wire _net_401;
  wire _net_402;
  wire _net_403;
  wire _net_404;
  wire _net_405;
  wire _net_406;
  wire _net_407;
  wire _net_408;
  wire _net_409;
  wire _net_410;
  wire _net_411;
  wire _net_412;
  wire _net_413;
  wire _net_414;
  wire _net_415;
  wire _net_416;
  wire _net_417;
  wire _net_418;
  wire _net_419;
  wire _net_420;
  wire _net_421;
  wire _net_422;
  wire _net_423;
  wire _net_424;
  wire _net_425;
  wire _net_426;
  wire _net_427;
  wire _net_428;
  wire _net_429;
  wire _net_430;
  wire _net_431;
  wire _net_432;
  wire _net_433;
  wire _net_434;
  wire _net_435;
  wire _net_436;
  wire _net_437;
  wire _net_438;
  wire _net_439;
  wire _net_440;
  wire _net_441;
  wire _net_442;
  wire _net_443;
  wire _net_444;
  wire _net_445;
  wire _net_446;
  wire _net_447;
  wire _net_448;
  wire _net_449;
  wire _net_450;
  wire _net_451;
  wire _net_452;
  wire _net_453;
  wire _net_454;
  wire _net_455;
  wire _net_456;
  wire _net_457;
  wire _net_458;
  wire _net_459;
  wire _net_460;
  wire _net_461;
  wire _net_462;
  wire _net_463;
  wire _net_464;
  wire _net_465;
  wire _net_466;
  wire _net_467;
  wire _net_468;
  wire _net_469;
  wire _net_470;
  wire _net_471;
  wire _net_472;
  wire _net_473;
  wire _net_474;
  wire _net_475;
  wire _net_476;
  wire _net_477;
  wire _net_478;
  wire _net_479;
  wire _net_480;
  wire _net_481;
  wire _net_482;
  wire _net_483;
  wire _net_484;
  wire _net_485;
  wire _net_486;
  wire _net_487;
  wire _net_488;
  wire _net_489;
  wire _net_490;
  wire _net_491;
  wire _net_492;
  wire _net_493;
  wire _net_494;
  wire _net_495;
  wire _net_496;
  wire _net_497;
  wire _net_498;
  wire _net_499;
  wire _net_500;
  wire _net_501;
  wire _net_502;
  wire _net_503;
  wire _net_504;
  wire _net_505;
  wire _net_506;
  wire _net_507;
  wire _net_508;
  wire _net_509;
  wire _net_510;
  wire _net_511;
  wire _net_512;
  wire _net_513;
  wire _net_514;
  wire _net_515;
  wire _net_516;
  wire _net_517;
  wire _net_518;
  wire _net_519;
  wire _net_520;
  wire _net_521;
  wire _net_522;
  wire _net_523;
  wire _net_524;
  wire _net_525;
  wire _net_526;
  wire _net_527;
  wire _net_528;
  wire _net_529;
  wire _net_530;
  wire _net_531;
  wire _net_532;
  wire _net_533;
  wire _net_534;
  wire _net_535;
  wire _net_536;
  wire _net_537;
  wire _net_538;
  wire _net_539;
  wire _net_540;
  wire _net_541;
  wire _net_542;
  wire _net_543;
  wire _net_544;
  wire _net_545;
  wire _net_546;
  wire _net_547;
  wire _net_548;
  wire _net_549;
  wire _net_550;
  wire _net_551;
  wire _net_552;
  wire _net_553;
  wire _net_554;
  wire _net_555;
  wire _net_556;
  wire _net_557;
  wire _net_558;
  wire _net_559;
  wire _net_560;
  wire _net_561;
  wire _net_562;
  wire _net_563;
  wire _net_564;
  wire _net_565;
  wire _net_566;
  wire _net_567;
  wire _net_568;
  wire _net_569;
  wire _net_570;
  wire _net_571;
  wire _net_572;
  wire _net_573;
  wire _net_574;
  wire _net_575;
  wire _net_576;
  wire _net_577;
  wire _net_578;
  wire _net_579;
  wire _net_580;
  wire _net_581;
  wire _net_582;
  wire _net_583;
  wire _net_584;
  wire _net_585;
  wire _net_586;
  wire _net_587;
  wire _net_588;
  wire _net_589;
  wire _net_590;
  wire _net_591;
  wire _net_592;
  wire _net_593;
  wire _net_594;
  wire _net_595;
  wire _net_596;
  wire _net_597;
  wire _net_598;
  wire _net_599;
  wire _net_600;
  wire _net_601;
  wire _net_602;
  wire _net_603;
  wire _net_604;
  wire _net_605;
  wire _net_606;
  wire _net_607;
  wire _net_608;
  wire _net_609;
  wire _net_610;
  wire _net_611;
  wire _net_612;
  wire _net_613;
  wire _net_614;
  wire _net_615;
  wire _net_616;
  wire _net_617;
  wire _net_618;
  wire _net_619;
  wire _net_620;
  wire _net_621;
  wire _net_622;
  wire _net_623;
  wire _net_624;
  wire _net_625;
  wire _net_626;
  wire _net_627;
  wire _net_628;
  wire _net_629;
  wire _net_630;
  wire _net_631;
  wire _net_632;
  wire _net_633;
  wire _net_634;
  wire _net_635;
  wire _net_636;
  wire _net_637;
  wire _net_638;
  wire _net_639;
  wire _net_640;
  wire _net_641;
  wire _net_642;
  wire _net_643;
  wire _net_644;
  wire _net_645;
  wire _net_646;
  wire _net_647;
  wire _net_648;
  wire _net_649;
  wire _net_650;
  wire _net_651;
  wire _net_652;
  wire _net_653;
  wire _net_654;
  wire _net_655;
  wire _net_656;
  wire _net_657;
  wire _net_658;
  wire _net_659;
  wire _net_660;
  wire _net_661;
  wire _net_662;
  wire _net_663;
  wire _net_664;
  wire _net_665;
  wire _net_666;
  wire _net_667;
  wire _net_668;
  wire _net_669;
  wire _net_670;
  wire _net_671;
  wire _net_672;
  wire _net_673;
  wire _net_674;
  wire _net_675;
  wire _net_676;
  wire _net_677;
  wire _net_678;
  wire _net_679;
  wire _net_680;
  wire _net_681;
  wire _net_682;
  wire _net_683;
  wire _net_684;
  wire _net_685;
  wire _net_686;
  wire _net_687;
  wire _net_688;
  wire _net_689;
  wire _net_690;
  wire _net_691;
  wire _net_692;
  wire _net_693;
  wire _net_694;
  wire _net_695;
  wire _net_696;
  wire _net_697;
  wire _net_698;
  wire _net_699;
  wire _net_700;
  wire _net_701;
  wire _net_702;
  wire _net_703;
  wire _net_704;
  wire _net_705;
  wire _net_706;
  wire _net_707;
  wire _net_708;
  wire _net_709;
  wire _net_710;
  wire _net_711;
  wire _net_712;
  wire _net_713;
  wire _net_714;
  wire _net_715;
  wire _net_716;
  wire _net_717;
  wire _net_718;
  wire _net_719;
  wire _net_720;
  wire _net_721;
  wire _net_722;
  wire _net_723;
  wire _net_724;
  wire _net_725;
  wire _net_726;
  wire _net_727;
  wire _net_728;
  wire _net_729;
  wire _net_730;
  wire _net_731;
  wire _net_732;
  wire _net_733;
  wire _net_734;
  wire _net_735;
  wire _net_736;
  wire _net_737;
  wire _net_738;
  wire _net_739;
  wire _net_740;
  wire _net_741;
  wire _net_742;
  wire _net_743;
  wire _net_744;
  wire _net_745;
  wire _net_746;
  wire _net_747;
  wire _net_748;
  wire _net_749;
  wire _net_750;
  wire _net_751;
  wire _net_752;
  wire _net_753;
  wire _net_754;
  wire _net_755;
  wire _net_756;
  wire _net_757;
  wire _net_758;
  wire _net_759;
  wire _net_760;
  wire _net_761;
  wire _net_762;
  wire _net_763;
  wire _net_764;
  wire _net_765;
  wire _net_766;
  wire _net_767;
  wire _net_768;
  wire _net_769;
  wire _net_770;
  wire _net_771;
  wire _net_772;
  wire _net_773;
  wire _net_774;
  wire _net_775;
  wire _net_776;
  wire _net_777;
  wire _net_778;
  wire _net_779;
  wire _net_780;
  wire _net_781;
  wire _net_782;
  wire _net_783;
  wire _net_784;
  wire _net_785;
  wire _net_786;
  wire _net_787;
  wire _net_788;
  wire _net_789;
  wire _net_790;
  wire _net_791;
  wire _net_792;
  wire _net_793;
  wire _net_794;
  wire _net_795;
  wire _net_796;
  wire _net_797;
  wire _net_798;
  wire _net_799;
  wire _net_800;
  wire _net_801;
  wire _net_802;
  wire _net_803;
  wire _net_804;
  wire _net_805;
  wire _net_806;
  wire _net_807;
  wire _net_808;
  wire _net_809;
  wire _net_810;
  wire _net_811;
  wire _net_812;
  wire _net_813;
  wire _net_814;
  wire _net_815;
  wire _net_816;
  wire _net_817;
  wire _net_818;
  wire _net_819;
  wire _net_820;
  wire _net_821;
  wire _net_822;
  wire _net_823;
  wire _net_824;
  wire _net_825;
  wire _net_826;
  wire _net_827;
  wire _net_828;
  wire _net_829;
  wire _net_830;
  wire _net_831;
  wire _net_832;
  wire _net_833;
  wire _net_834;
  wire _net_835;
  wire _net_836;
  wire _net_837;
  wire _net_838;
  wire _net_839;
  wire _net_840;
  wire _net_841;
  wire _net_842;
  wire _net_843;
  wire _net_844;
  wire _net_845;
  wire _net_846;
  wire _net_847;
  wire _net_848;
  wire _net_849;
  wire _net_850;
  wire _net_851;
  wire _net_852;
  wire _net_853;
  wire _net_854;
  wire _net_855;
  wire _net_856;
  wire _net_857;
  wire _net_858;
  wire _net_859;
  wire _net_860;
  wire _net_861;
  wire _net_862;
  wire _net_863;
  wire _net_864;
  wire _net_865;
  wire _net_866;
  wire _net_867;
  wire _net_868;
  wire _net_869;
  wire _net_870;
  wire _net_871;
  wire _net_872;
  wire _net_873;
  wire _net_874;
  wire _net_875;
  wire _net_876;
  wire _net_877;
  wire _net_878;
  wire _net_879;
  wire _net_880;
  wire _net_881;
  wire _net_882;
  wire _net_883;
  wire _net_884;
  wire _net_885;
  wire _net_886;
  wire _net_887;
  wire _net_888;
  wire _net_889;
  wire _net_890;
  wire _net_891;
  wire _net_892;
  wire _net_893;
  wire _net_894;
  wire _net_895;
  wire _net_896;
  wire _net_897;
  wire _net_898;
  wire _net_899;
  wire _net_900;
  wire _net_901;
  wire _net_902;
  wire _net_903;
  wire _net_904;
  wire _net_905;
  wire _net_906;
  wire _net_907;
  wire _net_908;
  wire _net_909;
  wire _net_910;
  wire _net_911;
  wire _net_912;
  wire _net_913;
  wire _net_914;
  wire _net_915;
  wire _net_916;
  wire _net_917;
  wire _net_918;
  wire _net_919;
  wire _net_920;
  wire _net_921;
  wire _net_922;
  wire _net_923;
  wire _net_924;
  wire _net_925;
  wire _net_926;
  wire _net_927;
  wire _net_928;
  wire _net_929;
  wire _net_930;
  wire _net_931;
  wire _net_932;
  wire _net_933;
  wire _net_934;
  wire _net_935;
  wire _net_936;
  wire _net_937;
  wire _net_938;
  wire _net_939;
  wire _net_940;
  wire _net_941;
  wire _net_942;
  wire _net_943;
  wire _net_944;
  wire _net_945;
  wire _net_946;
  wire _net_947;
  wire _net_948;
  wire _net_949;
  wire _net_950;
  wire _net_951;
  wire _net_952;
  wire _net_953;
  wire _net_954;
  wire _net_955;
  wire _net_956;
  wire _net_957;
  wire _net_958;
  wire _net_959;
  wire _net_960;
  wire _net_961;
  wire _net_962;
  wire _net_963;
  wire _net_964;
  wire _net_965;
  wire _net_966;
  wire _net_967;
  wire _net_968;
  wire _net_969;
  wire _net_970;
  wire _net_971;
  wire _net_972;
  wire _net_973;
  wire _net_974;
  wire _net_975;
  wire _net_976;
  wire _net_977;
  wire _net_978;
  wire _net_979;
  wire _net_980;
  wire _net_981;
  wire _net_982;
  wire _net_983;
  wire _net_984;
  wire _net_985;
  wire _net_986;
  wire _net_987;
  wire _net_988;
  wire _net_989;
  wire _net_990;
  wire _net_991;
  wire _net_992;
  wire _net_993;
  wire _net_994;
  wire _net_995;
  wire _net_996;
  wire _net_997;
  wire _net_998;
  wire _net_999;
  wire _net_1000;
  wire _net_1001;
  wire _net_1002;
  wire _net_1003;
  wire _net_1004;
  wire _net_1005;
  wire _net_1006;
  wire _net_1007;
  wire _net_1008;
  wire _net_1009;
  wire _net_1010;
  wire _net_1011;
  wire _net_1012;
  wire _net_1013;
  wire _net_1014;
  wire _net_1015;
  wire _net_1016;
  wire _net_1017;
  wire _net_1018;
  wire _net_1019;
  wire _net_1020;
  wire _net_1021;
  wire _net_1022;
  wire _net_1023;
  wire _net_1024;
  wire _net_1025;
  wire _net_1026;
  wire _net_1027;
  wire _net_1028;
  wire _net_1029;
  wire _net_1030;
  wire _net_1031;
  wire _net_1032;
  wire _net_1033;
  wire _net_1034;
  wire _net_1035;
  wire _net_1036;
  wire _net_1037;
  wire _net_1038;
  wire _net_1039;
  wire _net_1040;
  wire _net_1041;
  wire _net_1042;
  wire _net_1043;
  wire _net_1044;
  wire _net_1045;
  wire _net_1046;
  wire _net_1047;
  wire _net_1048;
  wire _net_1049;
  wire _net_1050;
  wire _net_1051;
  wire _net_1052;
  wire _net_1053;
  wire _net_1054;
  wire _net_1055;
  wire _net_1056;
  wire _net_1057;
  wire _net_1058;
  wire _net_1059;
  wire _net_1060;
  wire _net_1061;
  wire _net_1062;
  wire _net_1063;
  wire _net_1064;
  wire _net_1065;
  wire _net_1066;
  wire _net_1067;
  wire _net_1068;
  wire _net_1069;
  wire _net_1070;
  wire _net_1071;
  wire _net_1072;
  wire _net_1073;
  wire _net_1074;
  wire _net_1075;
  wire _net_1076;
  wire _net_1077;
  wire _net_1078;
  wire _net_1079;
  wire _net_1080;
  wire _net_1081;
  wire _net_1082;
  wire _net_1083;
  wire _net_1084;
  wire _net_1085;
  wire _net_1086;
  wire _net_1087;
  wire _net_1088;
  wire _net_1089;
  wire _net_1090;
  wire _net_1091;
  wire _net_1092;
  wire _net_1093;
  wire _net_1094;
  wire _net_1095;
  wire _net_1096;
  wire _net_1097;
  wire _net_1098;
  wire _net_1099;
  wire _net_1100;
  wire _net_1101;
  wire _net_1102;
  wire _net_1103;
  wire _net_1104;
  wire _net_1105;
  wire _net_1106;
  wire _net_1107;
  wire _net_1108;
  wire _net_1109;
  wire _net_1110;
  wire _net_1111;
  wire _net_1112;
  wire _net_1113;
  wire _net_1114;
  wire _net_1115;
  wire _net_1116;
  wire _net_1117;
  wire _net_1118;
  wire _net_1119;
  wire _net_1120;
  wire _net_1121;
  wire _net_1122;
  wire _net_1123;
  wire _net_1124;
  wire _net_1125;
  wire _net_1126;
  wire _net_1127;
  wire _net_1128;
  wire _net_1129;
  wire _net_1130;
  wire _net_1131;
  wire _net_1132;
  wire _net_1133;
  wire _net_1134;
  wire _net_1135;
  wire _net_1136;
  wire _net_1137;
  wire _net_1138;
  wire _net_1139;
  wire _net_1140;
  wire _net_1141;
  wire _net_1142;
  wire _net_1143;
  wire _net_1144;
  wire _net_1145;
  wire _net_1146;
  wire _net_1147;
  wire _net_1148;
  wire _net_1149;
  wire _net_1150;
  wire _net_1151;
  wire _net_1152;
  wire _net_1153;
  wire _net_1154;
  wire _net_1155;
  wire _net_1156;
  wire _net_1157;
  wire _net_1158;
  wire _net_1159;
  wire _net_1160;
  wire _net_1161;
  wire _net_1162;
  wire _net_1163;
  wire _net_1164;
  wire _net_1165;
  wire _net_1166;
  wire _net_1167;
  wire _net_1168;
  wire _net_1169;
  wire _net_1170;
  wire _net_1171;
  wire _net_1172;
  wire _net_1173;
  wire _net_1174;
  wire _net_1175;
  wire _net_1176;
  wire _net_1177;
  wire _net_1178;
  wire _net_1179;
  wire _net_1180;
  wire _net_1181;
  wire _net_1182;
  wire _net_1183;
  wire _net_1184;
  wire _net_1185;
  wire _net_1186;
  wire _net_1187;
  wire _net_1188;
  wire _net_1189;
  wire _net_1190;
  wire _net_1191;
  wire _net_1192;
  wire _net_1193;
  wire _net_1194;
  wire _net_1195;
  wire _net_1196;
  wire _net_1197;
  wire _net_1198;
  wire _net_1199;
  wire _net_1200;
  wire _net_1201;
  wire _net_1202;
  wire _net_1203;
  wire _net_1204;
  wire _net_1205;
  wire _net_1206;
  wire _net_1207;
  wire _net_1208;
  wire _net_1209;
  wire _net_1210;
  wire _net_1211;
  wire _net_1212;
  wire _net_1213;
  wire _net_1214;
  wire _net_1215;
  wire _net_1216;
  wire _net_1217;
  wire _net_1218;
  wire _net_1219;
  wire _net_1220;
  wire _net_1221;
  wire _net_1222;
  wire _net_1223;
  wire _net_1224;
  wire _net_1225;
  wire _net_1226;
  wire _net_1227;
  wire _net_1228;
  wire _net_1229;
  wire _net_1230;
  wire _net_1231;
  wire _net_1232;
  wire _net_1233;
  wire _net_1234;
  wire _net_1235;
  wire _net_1236;
  wire _net_1237;
  wire _net_1238;
  wire _net_1239;
  wire _net_1240;
  wire _net_1241;
  wire _net_1242;
  wire _net_1243;
  wire _net_1244;
  wire _net_1245;
  wire _net_1246;
  wire _net_1247;
  wire _net_1248;
  wire _net_1249;
  wire _net_1250;
  wire _net_1251;
  wire _net_1252;
  wire _net_1253;
  wire _net_1254;
  wire _net_1255;
  wire _net_1256;
  wire _net_1257;
  wire _net_1258;
  wire _net_1259;
  wire _net_1260;
  wire _net_1261;
  wire _net_1262;
  wire _net_1263;
  wire _net_1264;
  wire _net_1265;
  wire _net_1266;
  wire _net_1267;
  wire _net_1268;
  wire _net_1269;
  wire _net_1270;
  wire _net_1271;
  wire _net_1272;
  wire _net_1273;
  wire _net_1274;
  wire _net_1275;
  wire _net_1276;
  wire _net_1277;
  wire _net_1278;
  wire _net_1279;
  wire _net_1280;
  wire _net_1281;
  wire _net_1282;
  wire _net_1283;
  wire _net_1284;
  wire _net_1285;
  wire _net_1286;
  wire _net_1287;
  wire _net_1288;
  wire _net_1289;
  wire _net_1290;
  wire _net_1291;
  wire _net_1292;
  wire _net_1293;
  wire _net_1294;
  wire _net_1295;
  wire _net_1296;
  wire _net_1297;
  wire _net_1298;
  wire _net_1299;
  wire _net_1300;
  wire _net_1301;
  wire _net_1302;
  wire _net_1303;
  wire _net_1304;
  wire _net_1305;
  wire _net_1306;
  wire _net_1307;
  wire _net_1308;
  wire _net_1309;
  wire _net_1310;
  wire _net_1311;
  wire _net_1312;
  wire _net_1313;
  wire _net_1314;
  wire _net_1315;
  wire _net_1316;
  wire _net_1317;
  wire _net_1318;
  wire _net_1319;
  wire _net_1320;
  wire _net_1321;
  wire _net_1322;
  wire _net_1323;
  wire _net_1324;
  wire _net_1325;
  wire _net_1326;
  wire _net_1327;
  wire _net_1328;
  wire _net_1329;
  wire _net_1330;
  wire _net_1331;
  wire _net_1332;
  wire _net_1333;
  wire _net_1334;
  wire _net_1335;
  wire _net_1336;
  wire _net_1337;
  wire _net_1338;
  wire _net_1339;
  wire _net_1340;
  wire _net_1341;
  wire _net_1342;
  wire _net_1343;
  wire _net_1344;
  wire _net_1345;
  wire _net_1346;
  wire _net_1347;
  wire _net_1348;
  wire _net_1349;
  wire _net_1350;
  wire _net_1351;
  wire _net_1352;
  wire _net_1353;
  wire _net_1354;
  wire _net_1355;
  wire _net_1356;
  wire _net_1357;
  wire _net_1358;
  wire _net_1359;
  wire _net_1360;
  wire _net_1361;
  wire _net_1362;
  wire _net_1363;
  wire _net_1364;
  wire _net_1365;
  wire _net_1366;
  wire _net_1367;
  wire _net_1368;
  wire _net_1369;
  wire _net_1370;
  wire _net_1371;
  wire _net_1372;
  wire _net_1373;
  wire _net_1374;
  wire _net_1375;
  wire _net_1376;
  wire _net_1377;
  wire _net_1378;
  wire _net_1379;
  wire _net_1380;
  wire _net_1381;
  wire _net_1382;
  wire _net_1383;
  wire _net_1384;
  wire _net_1385;
  wire _net_1386;
  wire _net_1387;
  wire _net_1388;
  wire _net_1389;
  wire _net_1390;
  wire _net_1391;
  wire _net_1392;
  wire _net_1393;
  wire _net_1394;
  wire _net_1395;
  wire _net_1396;
  wire _net_1397;
  wire _net_1398;
  wire _net_1399;
  wire _net_1400;
  wire _net_1401;
  wire _net_1402;
  wire _net_1403;
  wire _net_1404;
  wire _net_1405;
  wire _net_1406;
  wire _net_1407;
  wire _net_1408;
  wire _net_1409;
  wire _net_1410;
  wire _net_1411;
  wire _net_1412;
  wire _net_1413;
  wire _net_1414;
  wire _net_1415;
  wire _net_1416;
  wire _net_1417;
  wire _net_1418;
  wire _net_1419;
  wire _net_1420;
  wire _net_1421;
  wire _net_1422;
  wire _net_1423;
  wire _net_1424;
  wire _net_1425;
  wire _net_1426;
  wire _net_1427;
  wire _net_1428;
  wire _net_1429;
  wire _net_1430;
  wire _net_1431;
  wire _net_1432;
  wire _net_1433;
  wire _net_1434;
  wire _net_1435;
  wire _net_1436;
  wire _net_1437;
  wire _net_1438;
  wire _net_1439;
  wire _net_1440;
  wire _net_1441;
  wire _net_1442;
  wire _net_1443;
  wire _net_1444;
  wire _net_1445;
  wire _net_1446;
  wire _net_1447;
  wire _net_1448;
  wire _net_1449;
  wire _net_1450;
  wire _net_1451;
  wire _net_1452;
  wire _net_1453;
  wire _net_1454;
  wire _net_1455;
  wire _net_1456;
  wire _net_1457;
  wire _net_1458;
  wire _net_1459;
  wire _net_1460;
  wire _net_1461;
  wire _net_1462;
  wire _net_1463;
  wire _net_1464;
  wire _net_1465;
  wire _net_1466;
  wire _net_1467;
  wire _net_1468;
  wire _net_1469;
  wire _net_1470;
  wire _net_1471;
  wire _net_1472;
  wire _net_1473;
  wire _net_1474;
  wire _net_1475;
  wire _net_1476;
  wire _net_1477;
  wire _net_1478;
  wire _net_1479;
  wire _net_1480;
  wire _net_1481;
  wire _net_1482;
  wire _net_1483;
  wire _net_1484;
  wire _net_1485;
  wire _net_1486;
  wire _net_1487;
  wire _net_1488;
  wire _net_1489;
  wire _net_1490;
  wire _net_1491;
  wire _net_1492;
  wire _net_1493;
  wire _net_1494;
  wire _net_1495;
  wire _net_1496;
  wire _net_1497;
  wire _net_1498;
  wire _net_1499;
  wire _net_1500;
  wire _net_1501;
  wire _net_1502;
  wire _net_1503;
  wire _net_1504;
  wire _net_1505;
  wire _net_1506;
  wire _net_1507;
  wire _net_1508;
  wire _net_1509;
  wire _net_1510;
  wire _net_1511;
  wire _net_1512;
  wire _net_1513;
  wire _net_1514;
  wire _net_1515;
  wire _net_1516;
  wire _net_1517;
  wire _net_1518;
  wire _net_1519;
  wire _net_1520;
  wire _net_1521;
  wire _net_1522;
  wire _net_1523;
  wire _net_1524;
  wire _net_1525;
  wire _net_1526;
  wire _net_1527;
  wire _net_1528;
  wire _net_1529;
  wire _net_1530;
  wire _net_1531;
  wire _net_1532;
  wire _net_1533;
  wire _net_1534;
  wire _net_1535;
  wire _net_1536;
  wire _net_1537;
  wire _net_1538;
  wire _net_1539;
  wire _net_1540;
  wire _net_1541;
  wire _net_1542;
  wire _net_1543;
  wire _net_1544;
  wire _net_1545;
  wire _net_1546;
  wire _net_1547;
  wire _net_1548;
  wire _net_1549;
  wire _net_1550;
  wire _net_1551;
  wire _net_1552;
  wire _net_1553;
  wire _net_1554;
  wire _net_1555;
  wire _net_1556;
  wire _net_1557;
  wire _net_1558;
  wire _net_1559;
  wire _net_1560;
  wire _net_1561;
  wire _net_1562;
  wire _net_1563;
  wire _net_1564;
  wire _net_1565;
  wire _net_1566;
  wire _net_1567;
  wire _net_1568;
  wire _net_1569;
  wire _net_1570;
  wire _net_1571;
  wire _net_1572;
  wire _net_1573;
  wire _net_1574;
  wire _net_1575;
  wire _net_1576;
  wire _net_1577;
  wire _net_1578;
  wire _net_1579;
  wire _net_1580;
  wire _net_1581;
  wire _net_1582;
  wire _net_1583;
  wire _net_1584;
  wire _net_1585;
  wire _net_1586;
  wire _net_1587;
  wire _net_1588;
  wire _net_1589;
  wire _net_1590;
  wire _net_1591;
  wire _net_1592;
  wire _net_1593;
  wire _net_1594;
  wire _net_1595;
  wire _net_1596;
  wire _net_1597;
  wire _net_1598;
  wire _net_1599;
  wire _net_1600;
  wire _net_1601;
  wire _net_1602;
  wire _net_1603;
  wire _net_1604;
  wire _net_1605;
  wire _net_1606;
  wire _net_1607;
  wire _net_1608;
  wire _net_1609;
  wire _net_1610;
  wire _net_1611;
  wire _net_1612;
  wire _net_1613;
  wire _net_1614;
  wire _net_1615;
  wire _net_1616;
  wire _net_1617;
  wire _net_1618;
  wire _net_1619;
  wire _net_1620;
  wire _net_1621;
  wire _net_1622;
  wire _net_1623;
  wire _net_1624;
  wire _net_1625;
  wire _net_1626;
  wire _net_1627;
  wire _net_1628;
  wire _net_1629;
  wire _net_1630;
  wire _net_1631;
  wire _net_1632;
  wire _net_1633;
  wire _net_1634;
  wire _net_1635;
  wire _net_1636;
  wire _net_1637;
  wire _net_1638;
  wire _net_1639;
  wire _net_1640;
  wire _net_1641;
  wire _net_1642;
  wire _net_1643;
  wire _net_1644;
  wire _net_1645;
  wire _net_1646;
  wire _net_1647;
  wire _net_1648;
  wire _net_1649;
  wire _net_1650;
  wire _net_1651;
  wire _net_1652;
  wire _net_1653;
  wire _net_1654;
  wire _net_1655;
  wire _net_1656;
  wire _net_1657;
  wire _net_1658;
  wire _net_1659;
  wire _net_1660;
  wire _net_1661;
  wire _net_1662;
  wire _net_1663;
  wire _net_1664;
  wire _net_1665;
  wire _net_1666;
  wire _net_1667;
  wire _net_1668;
  wire _net_1669;
  wire _net_1670;
  wire _net_1671;
  wire _net_1672;
  wire _net_1673;
  wire _net_1674;
  wire _net_1675;
  wire _net_1676;
  wire _net_1677;
  wire _net_1678;
  wire _net_1679;
  wire _net_1680;
  wire _net_1681;
  wire _net_1682;
  wire _net_1683;
  wire _net_1684;
  wire _net_1685;
  wire _net_1686;
  wire _net_1687;
  wire _net_1688;
  wire _net_1689;
  wire _net_1690;
  wire _net_1691;
  wire _net_1692;
  wire _net_1693;
  wire _net_1694;
  wire _net_1695;
  wire _net_1696;
  wire _net_1697;
  wire _net_1698;
  wire _net_1699;
  wire _net_1700;
  wire _net_1701;
  wire _net_1702;
  wire _net_1703;
  wire _net_1704;
  wire _net_1705;
  wire _net_1706;
  wire _net_1707;
  wire _net_1708;
  wire _net_1709;
  wire _net_1710;
  wire _net_1711;
  wire _net_1712;
  wire _net_1713;
  wire _net_1714;
  wire _net_1715;
  wire _net_1716;
  wire _net_1717;
  wire _net_1718;
  wire _net_1719;
  wire _net_1720;
  wire _net_1721;
  wire _net_1722;
  wire _net_1723;
  wire _net_1724;
  wire _net_1725;
  wire _net_1726;
  wire _net_1727;
  wire _net_1728;
  wire _net_1729;
  wire _net_1730;
  wire _net_1731;
  wire _net_1732;
  wire _net_1733;
  wire _net_1734;
  wire _net_1735;
  wire _net_1736;
  wire _net_1737;
  wire _net_1738;
  wire _net_1739;
  wire _net_1740;
  wire _net_1741;
  wire _net_1742;
  wire _net_1743;
  wire _net_1744;
  wire _net_1745;
  wire _net_1746;
  wire _net_1747;
  wire _net_1748;
  wire _net_1749;
  wire _net_1750;
  wire _net_1751;
  wire _net_1752;
  wire _net_1753;
  wire _net_1754;
  wire _net_1755;
  wire _net_1756;
  wire _net_1757;
  wire _net_1758;
  wire _net_1759;
  wire _net_1760;
  wire _net_1761;
  wire _net_1762;
  wire _net_1763;
  wire _net_1764;
  wire _net_1765;
  wire _net_1766;
  wire _net_1767;
  wire _net_1768;
  wire _net_1769;
  wire _net_1770;
  wire _net_1771;
  wire _net_1772;
  wire _net_1773;
  wire _net_1774;
  wire _net_1775;
  wire _net_1776;
  wire _net_1777;
  wire _net_1778;
  wire _net_1779;
  wire _net_1780;
  wire _net_1781;
  wire _net_1782;
  wire _net_1783;
  wire _net_1784;
  wire _net_1785;
  wire _net_1786;
  wire _net_1787;
  wire _net_1788;
  wire _net_1789;
  wire _net_1790;
  wire _net_1791;
  wire _net_1792;
  wire _net_1793;
  wire _net_1794;
  wire _net_1795;
  wire _net_1796;
  wire _net_1797;
  wire _net_1798;
  wire _net_1799;
  wire _net_1800;
  wire _net_1801;
  wire _net_1802;
  wire _net_1803;
  wire _net_1804;
  wire _net_1805;
  wire _net_1806;
  wire _net_1807;
  wire _net_1808;
  wire _net_1809;
  wire _net_1810;
  wire _net_1811;
  wire _net_1812;
  wire _net_1813;
  wire _net_1814;
  wire _net_1815;
  wire _net_1816;
  wire _net_1817;
  wire _net_1818;
  wire _net_1819;
  wire _net_1820;
  wire _net_1821;
  wire _net_1822;
  wire _net_1823;
  wire _net_1824;
  wire _net_1825;
  wire _net_1826;
  wire _net_1827;
  wire _net_1828;
  wire _net_1829;
  wire _net_1830;
  wire _net_1831;
  wire _net_1832;
  wire _net_1833;
  wire _net_1834;
  wire _net_1835;
  wire _net_1836;
  wire _net_1837;
  wire _net_1838;
  wire _net_1839;
  wire _net_1840;
  wire _net_1841;
  wire _net_1842;
  wire _net_1843;
  wire _net_1844;
  wire _net_1845;
  wire _net_1846;
  wire _net_1847;
  wire _net_1848;
  wire _net_1849;
  wire _net_1850;
  wire _net_1851;
  wire _net_1852;
  wire _net_1853;
  wire _net_1854;
  wire _net_1855;
  wire _net_1856;
  wire _net_1857;
  wire _net_1858;
  wire _net_1859;
  wire _net_1860;
  wire _net_1861;
  wire _net_1862;
  wire _net_1863;
  wire _net_1864;
  wire _net_1865;
  wire _net_1866;
  wire _net_1867;
  wire _net_1868;
  wire _net_1869;
  wire _net_1870;
  wire _net_1871;
  wire _net_1872;
  wire _net_1873;
  wire _net_1874;
  wire _net_1875;
  wire _net_1876;
  wire _net_1877;
  wire _net_1878;
  wire _net_1879;
  wire _net_1880;
  wire _net_1881;
  wire _net_1882;
  wire _net_1883;
  wire _net_1884;
  wire _net_1885;
  wire _net_1886;
  wire _net_1887;
  wire _net_1888;
  wire _net_1889;
  wire _net_1890;
  wire _net_1891;
  wire _net_1892;
  wire _net_1893;
  wire _net_1894;
  wire _net_1895;
  wire _net_1896;
  wire _net_1897;
  wire _net_1898;
  wire _net_1899;
  wire _net_1900;
  wire _net_1901;
  wire _net_1902;
  wire _net_1903;
  wire _net_1904;
  wire _net_1905;
  wire _net_1906;
  wire _net_1907;
  wire _net_1908;
  wire _net_1909;
  wire _net_1910;
  wire _net_1911;
  wire _net_1912;
  wire _net_1913;
  wire _net_1914;
  wire _net_1915;
  wire _net_1916;
  wire _net_1917;
  wire _net_1918;
  wire _net_1919;
  wire _net_1920;
  wire _net_1921;
  wire _net_1922;
  wire _net_1923;
  wire _net_1924;
  wire _net_1925;
  wire _net_1926;
  wire _net_1927;
  wire _net_1928;
  wire _net_1929;
  wire _net_1930;
  wire _net_1931;
  wire _net_1932;
  wire _net_1933;
  wire _net_1934;
  wire _net_1935;
  wire _net_1936;
  wire _net_1937;
  wire _net_1938;
  wire _net_1939;
  wire _net_1940;
  wire _net_1941;
  wire _net_1942;
  wire _net_1943;
  wire _net_1944;
  wire _net_1945;
  wire _net_1946;
  wire _net_1947;
  wire _net_1948;
  wire _net_1949;
  wire _net_1950;
  wire _net_1951;
  wire _net_1952;
  wire _net_1953;
  wire _net_1954;
  wire _net_1955;
  wire _net_1956;
  wire _net_1957;
  wire _net_1958;
  wire _net_1959;
  wire _net_1960;
  wire _net_1961;
  wire _net_1962;
  wire _net_1963;
  wire _net_1964;
  wire _net_1965;
  wire _net_1966;
  wire _net_1967;
  wire _net_1968;
  wire _net_1969;
  wire _net_1970;
  wire _net_1971;
  wire _net_1972;
  wire _net_1973;
  wire _net_1974;
  wire _net_1975;
  wire _net_1976;
  wire _net_1977;
  wire _net_1978;
  wire _net_1979;
  wire _net_1980;
  wire _net_1981;
  wire _net_1982;
  wire _net_1983;
  wire _net_1984;
  wire _net_1985;
  wire _net_1986;
  wire _net_1987;
  wire _net_1988;
  wire _net_1989;
  wire _net_1990;
  wire _net_1991;
  wire _net_1992;
  wire _net_1993;
  wire _net_1994;
  wire _net_1995;
  wire _net_1996;
  wire _net_1997;
  wire _net_1998;
  wire _net_1999;
  wire _net_2000;
  wire _net_2001;
  wire _net_2002;
  wire _net_2003;
  wire _net_2004;
  wire _net_2005;
  wire _net_2006;
  wire _net_2007;
  wire _net_2008;
  wire _net_2009;
  wire _net_2010;
  wire _net_2011;
  wire _net_2012;
  wire _net_2013;
  wire _net_2014;
  wire _net_2015;
  wire _net_2016;
  wire _net_2017;
  wire _net_2018;
  wire _net_2019;
  wire _net_2020;
  wire _net_2021;
  wire _net_2022;
  wire _net_2023;
  wire _net_2024;
  wire _net_2025;
  wire _net_2026;
  wire _net_2027;
  wire _net_2028;
  wire _net_2029;
  wire _net_2030;
  wire _net_2031;
  wire _net_2032;
  wire _net_2033;
  wire _net_2034;
  wire _net_2035;
  wire _net_2036;
  wire _net_2037;
  wire _net_2038;
  wire _net_2039;
  wire _net_2040;
  wire _net_2041;
  wire _net_2042;
  wire _net_2043;
  wire _net_2044;
  wire _net_2045;
  wire _net_2046;
  wire _net_2047;
  wire _net_2048;
  wire _net_2049;
  wire _net_2050;
  wire _net_2051;
  wire _net_2052;
  wire _net_2053;
  wire _net_2054;
  wire _net_2055;
  wire _net_2056;
  wire _net_2057;
  wire _net_2058;
  wire _net_2059;
  wire _net_2060;
  wire _net_2061;
  wire _net_2062;
  wire _net_2063;
  wire _net_2064;
  wire _net_2065;
  wire _net_2066;
  wire _net_2067;
  wire _net_2068;
  wire _net_2069;
  wire _net_2070;
  wire _net_2071;
  wire _net_2072;
  wire _net_2073;
  wire _net_2074;
  wire _net_2075;
  wire _net_2076;
  wire _net_2077;
  wire _net_2078;
  wire _net_2079;
  wire _net_2080;
  wire _net_2081;
  wire _net_2082;
  wire _net_2083;
  wire _net_2084;
  wire _net_2085;
  wire _net_2086;
  wire _net_2087;
  wire _net_2088;
  wire _net_2089;
  wire _net_2090;
  wire _net_2091;
  wire _net_2092;
  wire _net_2093;
  wire _net_2094;
  wire _net_2095;
  wire _net_2096;
  wire _net_2097;
  wire _net_2098;
  wire _net_2099;
  wire _net_2100;
  wire _net_2101;
  wire _net_2102;
  wire _net_2103;
  wire _net_2104;
  wire _net_2105;
  wire _net_2106;
  wire _net_2107;
  wire _net_2108;
  wire _net_2109;
  wire _net_2110;
  wire _net_2111;
  wire _net_2112;
  wire _net_2113;
  wire _net_2114;
  wire _net_2115;
  wire _net_2116;
  wire _net_2117;
  wire _net_2118;
  wire _net_2119;
  wire _net_2120;
  wire _net_2121;
  wire _net_2122;
  wire _net_2123;
  wire _net_2124;
  wire _net_2125;
  wire _net_2126;
  wire _net_2127;
  wire _net_2128;
  wire _net_2129;
  wire _net_2130;
  wire _net_2131;
  wire _net_2132;
  wire _net_2133;
  wire _net_2134;
  wire _net_2135;
  wire _net_2136;
  wire _net_2137;
  wire _net_2138;
  wire _net_2139;
  wire _net_2140;
  wire _net_2141;
  wire _net_2142;
  wire _net_2143;
  wire _net_2144;
  wire _net_2145;
  wire _net_2146;
  wire _net_2147;
  wire _net_2148;
  wire _net_2149;
  wire _net_2150;
  wire _net_2151;
  wire _net_2152;
  wire _net_2153;
  wire _net_2154;
  wire _net_2155;
  wire _net_2156;
  wire _net_2157;
  wire _net_2158;
  wire _net_2159;
  wire _net_2160;
  wire _net_2161;
  wire _net_2162;
  wire _net_2163;
  wire _net_2164;
  wire _net_2165;
  wire _net_2166;
  wire _net_2167;
  wire _net_2168;
  wire _net_2169;
  wire _net_2170;
  wire _net_2171;
  wire _net_2172;
  wire _net_2173;
  wire _net_2174;
  wire _net_2175;
  wire _net_2176;
  wire _net_2177;
  wire _net_2178;
  wire _net_2179;
  wire _net_2180;
  wire _net_2181;
  wire _net_2182;
  wire _net_2183;
  wire _net_2184;
  wire _net_2185;
  wire _net_2186;
  wire _net_2187;
  wire _net_2188;
  wire _net_2189;
  wire _net_2190;
  wire _net_2191;
  wire _net_2192;
  wire _net_2193;
  wire _net_2194;
  wire _net_2195;
  wire _net_2196;
  wire _net_2197;
  wire _net_2198;
  wire _net_2199;
  wire _net_2200;
  wire _net_2201;
  wire _net_2202;
  wire _net_2203;
  wire _net_2204;
  wire _net_2205;
  wire _net_2206;
  wire _net_2207;
  wire _net_2208;
  wire _net_2209;
  wire _net_2210;
  wire _net_2211;
  wire _net_2212;
  wire _net_2213;
  wire _net_2214;
  wire _net_2215;
  wire _net_2216;
  wire _net_2217;
  wire _net_2218;
  wire _net_2219;
  wire _net_2220;
  wire _net_2221;
  wire _net_2222;
  wire _net_2223;
  wire _net_2224;
  wire _net_2225;
  wire _net_2226;
  wire _net_2227;
  wire _net_2228;
  wire _net_2229;
  wire _net_2230;
  wire _net_2231;
  wire _net_2232;
  wire _net_2233;
  wire _net_2234;
  wire _net_2235;
  wire _net_2236;
  wire _net_2237;
  wire _net_2238;
  wire _net_2239;
  wire _net_2240;
  wire _net_2241;
  wire _net_2242;
  wire _net_2243;
  wire _net_2244;
  wire _net_2245;
  wire _net_2246;
  wire _net_2247;
  wire _net_2248;
  wire _net_2249;
  wire _net_2250;
  wire _net_2251;
  wire _net_2252;
  wire _net_2253;
  wire _net_2254;
  wire _net_2255;
  wire _net_2256;
  wire _net_2257;
  wire _net_2258;
  wire _net_2259;
  wire _net_2260;
  wire _net_2261;
  wire _net_2262;
  wire _net_2263;
  wire _net_2264;
  wire _net_2265;
  wire _net_2266;
  wire _net_2267;
  wire _net_2268;
  wire _net_2269;
  wire _net_2270;
  wire _net_2271;
  wire _net_2272;
  wire _net_2273;
  wire _net_2274;
  wire _net_2275;
  wire _net_2276;
  wire _net_2277;
  wire _net_2278;
  wire _net_2279;
  wire _net_2280;
  wire _net_2281;
  wire _net_2282;
  wire _net_2283;
  wire _net_2284;
  wire _net_2285;
  wire _net_2286;
  wire _net_2287;
  wire _net_2288;
  wire _net_2289;
  wire _net_2290;
  wire _net_2291;
  wire _net_2292;
  wire _net_2293;
  wire _net_2294;
  wire _net_2295;
  wire _net_2296;
  wire _net_2297;
  wire _net_2298;
  wire _net_2299;
  wire _net_2300;
  wire _net_2301;
  wire _net_2302;
  wire _net_2303;
  wire _net_2304;
  wire _net_2305;
  wire _net_2306;
  wire _net_2307;
  wire _net_2308;
  wire _net_2309;
  wire _net_2310;
  wire _net_2311;
  wire _net_2312;
  wire _net_2313;
  wire _net_2314;
  wire _net_2315;
  wire _net_2316;
  wire _net_2317;
  wire _net_2318;
  wire _net_2319;
  wire _net_2320;
  wire _net_2321;
  wire _net_2322;
  wire _net_2323;
  wire _net_2324;
  wire _net_2325;
  wire _net_2326;
  wire _net_2327;
  wire _net_2328;
  wire _net_2329;
  wire _net_2330;
  wire _net_2331;
  wire _net_2332;
  wire _net_2333;
  wire _net_2334;
  wire _net_2335;
  wire _net_2336;
  wire _net_2337;
  wire _net_2338;
  wire _net_2339;
  wire _net_2340;
  wire _net_2341;
  wire _net_2342;
  wire _net_2343;
  wire _net_2344;
  wire _net_2345;
  wire _net_2346;
  wire _net_2347;
  wire _net_2348;
  wire _net_2349;
  wire _net_2350;
  wire _net_2351;
  wire _net_2352;
  wire _net_2353;
  wire _net_2354;
  wire _net_2355;
  wire _net_2356;
  wire _net_2357;
  wire _net_2358;
  wire _net_2359;
  wire _net_2360;
  wire _net_2361;
  wire _net_2362;
  wire _net_2363;
  wire _net_2364;
  wire _net_2365;
  wire _net_2366;
  wire _net_2367;
  wire _net_2368;
  wire _net_2369;
  wire _net_2370;
  wire _net_2371;
  wire _net_2372;
  wire _net_2373;
  wire _net_2374;
  wire _net_2375;
  wire _net_2376;
  wire _net_2377;
  wire _net_2378;
  wire _net_2379;
  wire _net_2380;
  wire _net_2381;
  wire _net_2382;
  wire _net_2383;
  wire _net_2384;
  wire _net_2385;
  wire _net_2386;
  wire _net_2387;
  wire _net_2388;
  wire _net_2389;
  wire _net_2390;
  wire _net_2391;
  wire _net_2392;
  wire _net_2393;
  wire _net_2394;
  wire _net_2395;
  wire _net_2396;
  wire _net_2397;
  wire _net_2398;
  wire _net_2399;
  wire _net_2400;
  wire _net_2401;
  wire _net_2402;
  wire _net_2403;
  wire _net_2404;
  wire _net_2405;
  wire _net_2406;
  wire _net_2407;
  wire _net_2408;
  wire _net_2409;
  wire _net_2410;
  wire _net_2411;
  wire _net_2412;
  wire _net_2413;
  wire _net_2414;
  wire _net_2415;
  wire _net_2416;
  wire _net_2417;
  wire _net_2418;
  wire _net_2419;
  wire _net_2420;
  wire _net_2421;
  wire _net_2422;
  wire _net_2423;
  wire _net_2424;
  wire _net_2425;
  wire _net_2426;
  wire _net_2427;
  wire _net_2428;
  wire _net_2429;
  wire _net_2430;
  wire _net_2431;
  wire _net_2432;
  wire _net_2433;
  wire _net_2434;
  wire _net_2435;
  wire _net_2436;
  wire _net_2437;
  wire _net_2438;
  wire _net_2439;
  wire _net_2440;
  wire _net_2441;
  wire _net_2442;
  wire _net_2443;
  wire _net_2444;
  wire _net_2445;
  wire _net_2446;
  wire _net_2447;
  wire _net_2448;
  wire _net_2449;
  wire _net_2450;
  wire _net_2451;
  wire _net_2452;
  wire _net_2453;
  wire _net_2454;
  wire _net_2455;
  wire _net_2456;
  wire _net_2457;
  wire _net_2458;
  wire _net_2459;
  wire _net_2460;
  wire _net_2461;
  wire _net_2462;
  wire _net_2463;
  wire _net_2464;
  wire _net_2465;
  wire _net_2466;
  wire _net_2467;
  wire _net_2468;
  wire _net_2469;
  wire _net_2470;
  wire _net_2471;
  wire _net_2472;
  wire _net_2473;
  wire _net_2474;
  wire _net_2475;
  wire _net_2476;
  wire _net_2477;
  wire _net_2478;
  wire _net_2479;
  wire _net_2480;
  wire _net_2481;
  wire _net_2482;
  wire _net_2483;
  wire _net_2484;
  wire _net_2485;
  wire _net_2486;
  wire _net_2487;
  wire _net_2488;
  wire _net_2489;
  wire _net_2490;
  wire _net_2491;
  wire _net_2492;
  wire _net_2493;
  wire _net_2494;
  wire _net_2495;
  wire _net_2496;
  wire _net_2497;
  wire _net_2498;
  wire _net_2499;
  wire _net_2500;
  wire _net_2501;
  wire _net_2502;
  wire _net_2503;
  wire _net_2504;
  wire _net_2505;
  wire _net_2506;
  wire _net_2507;
  wire _net_2508;
  wire _net_2509;
  wire _net_2510;
  wire _net_2511;
  wire _net_2512;
  wire _net_2513;
  wire _net_2514;
  wire _net_2515;
  wire _net_2516;
  wire _net_2517;
  wire _net_2518;
  wire _net_2519;
  wire _net_2520;
  wire _net_2521;
  wire _net_2522;
  wire _net_2523;
  wire _net_2524;
  wire _net_2525;
  wire _net_2526;
  wire _net_2527;
  wire _net_2528;
  wire _net_2529;
  wire _net_2530;
  wire _net_2531;
  wire _net_2532;
  wire _net_2533;
  wire _net_2534;
  wire _net_2535;
  wire _net_2536;
  wire _net_2537;
  wire _net_2538;
  wire _net_2539;
  wire _net_2540;
  wire _net_2541;
  wire _net_2542;
  wire _net_2543;
  wire _net_2544;
  wire _net_2545;
  wire _net_2546;
  wire _net_2547;
  wire _net_2548;
  wire _net_2549;
  wire _net_2550;
  wire _net_2551;
  wire _net_2552;
  wire _net_2553;
  wire _net_2554;
  wire _net_2555;
  wire _net_2556;
  wire _net_2557;
  wire _net_2558;
  wire _net_2559;
  wire _net_2560;
  wire _net_2561;
  wire _net_2562;
  wire _net_2563;
  wire _net_2564;
  wire _net_2565;
  wire _net_2566;
  wire _net_2567;
  wire _net_2568;
  wire _net_2569;
  wire _net_2570;
  wire _net_2571;
  wire _net_2572;
  wire _net_2573;
  wire _net_2574;
  wire _net_2575;
  wire _net_2576;
  wire _net_2577;
  wire _net_2578;
  wire _net_2579;
  wire _net_2580;
  wire _net_2581;
  wire _net_2582;
  wire _net_2583;
  wire _net_2584;
  wire _net_2585;
  wire _net_2586;
  wire _net_2587;
  wire _net_2588;
  wire _net_2589;
  wire _net_2590;
  wire _net_2591;
  wire _net_2592;
  wire _net_2593;
  wire _net_2594;
  wire _net_2595;
  wire _net_2596;
  wire _net_2597;
  wire _net_2598;
  wire _net_2599;
  wire _net_2600;
  wire _net_2601;
  wire _net_2602;
  wire _net_2603;
  wire _net_2604;
  wire _net_2605;
  wire _net_2606;
  wire _net_2607;
  wire _net_2608;
  wire _net_2609;
  wire _net_2610;
  wire _net_2611;
  wire _net_2612;
  wire _net_2613;
  wire _net_2614;
  wire _net_2615;
  wire _net_2616;
  wire _net_2617;
  wire _net_2618;
  wire _net_2619;
  wire _net_2620;
  wire _net_2621;
  wire _net_2622;
  wire _net_2623;
  wire _net_2624;
  wire _net_2625;
  wire _net_2626;
  wire _net_2627;
  wire _net_2628;
  wire _net_2629;
  wire _net_2630;
  wire _net_2631;
  wire _net_2632;
  wire _net_2633;
  wire _net_2634;
  wire _net_2635;
  wire _net_2636;
  wire _net_2637;
  wire _net_2638;
  wire _net_2639;
  wire _net_2640;
  wire _net_2641;
  wire _net_2642;
  wire _net_2643;
  wire _net_2644;
  wire _net_2645;
  wire _net_2646;
  wire _net_2647;
  wire _net_2648;
  wire _net_2649;
  wire _net_2650;
  wire _net_2651;
  wire _net_2652;
  wire _net_2653;
  wire _net_2654;
  wire _net_2655;
  wire _net_2656;
  wire _net_2657;
  wire _net_2658;
  wire _net_2659;
  wire _net_2660;
  wire _net_2661;
  wire _net_2662;
  wire _net_2663;
  wire _net_2664;
  wire _net_2665;
  wire _net_2666;
  wire _net_2667;
  wire _net_2668;
  wire _net_2669;
  wire _net_2670;
  wire _net_2671;
  wire _net_2672;
  wire _net_2673;
  wire _net_2674;
  wire _net_2675;
  wire _net_2676;
  wire _net_2677;
  wire _net_2678;
  wire _net_2679;
  wire _net_2680;
  wire _net_2681;
  wire _net_2682;
  wire _net_2683;
  wire _net_2684;
  wire _net_2685;
  wire _net_2686;
  wire _net_2687;
  wire _net_2688;
  wire _net_2689;
  wire _net_2690;
  wire _net_2691;
  wire _net_2692;
  wire _net_2693;
  wire _net_2694;
  wire _net_2695;
  wire _net_2696;
  wire _net_2697;
  wire _net_2698;
  wire _net_2699;
  wire _net_2700;
  wire _net_2701;
  wire _net_2702;
  wire _net_2703;
  wire _net_2704;
  wire _net_2705;
  wire _net_2706;
  wire _net_2707;
  wire _net_2708;
  wire _net_2709;
  wire _net_2710;
  wire _net_2711;
  wire _net_2712;
  wire _net_2713;
  wire _net_2714;
  wire _net_2715;
  wire _net_2716;
  wire _net_2717;
  wire _net_2718;
  wire _net_2719;
  wire _net_2720;
  wire _net_2721;
  wire _net_2722;
  wire _net_2723;
  wire _net_2724;
  wire _net_2725;
  wire _net_2726;
  wire _net_2727;
  wire _net_2728;
  wire _net_2729;
  wire _net_2730;
  wire _net_2731;
  wire _net_2732;
  wire _net_2733;
  wire _net_2734;
  wire _net_2735;
  wire _net_2736;
  wire _net_2737;
  wire _net_2738;
  wire _net_2739;
  wire _net_2740;
  wire _net_2741;
  wire _net_2742;
  wire _net_2743;
  wire _net_2744;
  wire _net_2745;
  wire _net_2746;
  wire _net_2747;
  wire _net_2748;
  wire _net_2749;
  wire _net_2750;
  wire _net_2751;
  wire _net_2752;
  wire _net_2753;
  wire _net_2754;
  wire _net_2755;
  wire _net_2756;
  wire _net_2757;
  wire _net_2758;
  wire _net_2759;
  wire _net_2760;
  wire _net_2761;
  wire _net_2762;
  wire _net_2763;
  wire _net_2764;
  wire _net_2765;
  wire _net_2766;
  wire _net_2767;
  wire _net_2768;
  wire _net_2769;
  wire _net_2770;
  wire _net_2771;
  wire _net_2772;
  wire _net_2773;
  wire _net_2774;
  wire _net_2775;
  wire _net_2776;
  wire _net_2777;
  wire _net_2778;
  wire _net_2779;
  wire _net_2780;
  wire _net_2781;
  wire _net_2782;
  wire _net_2783;
  wire _net_2784;
  wire _net_2785;
  wire _net_2786;
  wire _net_2787;
  wire _net_2788;
  wire _net_2789;
  wire _net_2790;
  wire _net_2791;
  wire _net_2792;
  wire _net_2793;
  wire _net_2794;
  wire _net_2795;
  wire _net_2796;
  wire _net_2797;
  wire _net_2798;
  wire _net_2799;
  wire _net_2800;
  wire _net_2801;
  wire _net_2802;
  wire _net_2803;
  wire _net_2804;
  wire _net_2805;
  wire _net_2806;
  wire _net_2807;
  wire _net_2808;
  wire _net_2809;
  wire _net_2810;
  wire _net_2811;
  wire _net_2812;
  wire _net_2813;
  wire _net_2814;
  wire _net_2815;
  wire _net_2816;
  wire _net_2817;
  wire _net_2818;
  wire _net_2819;
  wire _net_2820;
  wire _net_2821;
  wire _net_2822;
  wire _net_2823;
  wire _net_2824;
  wire _net_2825;
  wire _net_2826;
  wire _net_2827;
  wire _net_2828;
  wire _net_2829;
  wire _net_2830;
  wire _net_2831;
  wire _net_2832;
  wire _net_2833;
  wire _net_2834;
  wire _net_2835;
  wire _net_2836;
  wire _net_2837;
  wire _net_2838;
  wire _net_2839;
  wire _net_2840;
  wire _net_2841;
  wire _net_2842;
  wire _net_2843;
  wire _net_2844;
  wire _net_2845;
  wire _net_2846;
  wire _net_2847;
  wire _net_2848;
  wire _net_2849;
  wire _net_2850;
  wire _net_2851;
  wire _net_2852;
  wire _net_2853;
  wire _net_2854;
  wire _net_2855;
  wire _net_2856;
  wire _net_2857;
  wire _net_2858;
  wire _net_2859;
  wire _net_2860;
  wire _net_2861;
  wire _net_2862;
  wire _net_2863;
  wire _net_2864;
  wire _net_2865;
  wire _net_2866;
  wire _net_2867;
  wire _net_2868;
  wire _net_2869;
  wire _net_2870;
  wire _net_2871;
  wire _net_2872;
  wire _net_2873;
  wire _net_2874;
  wire _net_2875;
  wire _net_2876;
  wire _net_2877;
  wire _net_2878;
  wire _net_2879;
  wire _net_2880;
  wire _net_2881;
  wire _net_2882;
  wire _net_2883;
  wire _net_2884;
  wire _net_2885;
  wire _net_2886;
  wire _net_2887;
  wire _net_2888;
  wire _net_2889;
  wire _net_2890;
  wire _net_2891;
  wire _net_2892;
  wire _net_2893;
  wire _net_2894;
  wire _net_2895;
  wire _net_2896;
  wire _net_2897;
  wire _net_2898;
  wire _net_2899;
  wire _net_2900;
  wire _net_2901;
  wire _net_2902;
  wire _net_2903;
  wire _net_2904;
  wire _net_2905;
  wire _net_2906;
  wire _net_2907;
  wire _net_2908;
  wire _net_2909;
  wire _net_2910;
  wire _net_2911;
  wire _net_2912;
  wire _net_2913;
  wire _net_2914;
  wire _net_2915;
  wire _net_2916;
  wire _net_2917;
  wire _net_2918;
  wire _net_2919;
  wire _net_2920;
  wire _net_2921;
  wire _net_2922;
  wire _net_2923;
  wire _net_2924;
  wire _net_2925;
  wire _net_2926;
  wire _net_2927;
  wire _net_2928;
  wire _net_2929;
  wire _net_2930;
  wire _net_2931;
  wire _net_2932;
  wire _net_2933;
  wire _net_2934;
  wire _net_2935;
  wire _net_2936;
  wire _net_2937;
  wire _net_2938;
  wire _net_2939;
  wire _net_2940;
  wire _net_2941;
  wire _net_2942;
  wire _net_2943;
  wire _net_2944;
  wire _net_2945;
  wire _net_2946;
  wire _net_2947;
  wire _net_2948;
  wire _net_2949;
  wire _net_2950;
  wire _net_2951;
  wire _net_2952;
  wire _net_2953;
  wire _net_2954;
  wire _net_2955;
  wire _net_2956;
  wire _net_2957;
  wire _net_2958;
  wire _net_2959;
  wire _net_2960;
  wire _net_2961;
  wire _net_2962;
  wire _net_2963;
  wire _net_2964;
  wire _net_2965;
  wire _net_2966;
  wire _net_2967;
  wire _net_2968;
  wire _net_2969;
  wire _net_2970;
  wire _net_2971;
  wire _net_2972;
  wire _net_2973;
  wire _net_2974;
  wire _net_2975;
  wire _net_2976;
  wire _net_2977;
  wire _net_2978;
  wire _net_2979;
  wire _net_2980;
  wire _net_2981;
  wire _net_2982;
  wire _net_2983;
  wire _net_2984;
  wire _net_2985;
  wire _net_2986;
  wire _net_2987;
  wire _net_2988;
  wire _net_2989;
  wire _net_2990;
  wire _net_2991;
  wire _net_2992;
  wire _net_2993;
  wire _net_2994;
  wire _net_2995;
  wire _net_2996;
  wire _net_2997;
  wire _net_2998;
  wire _net_2999;
  wire _net_3000;
  wire _net_3001;
  wire _net_3002;
  wire _net_3003;
  wire _net_3004;
  wire _net_3005;
  wire _net_3006;
  wire _net_3007;
  wire _net_3008;
  wire _net_3009;
  wire _net_3010;
  wire _net_3011;
  wire _net_3012;
  wire _net_3013;
  wire _net_3014;
  wire _net_3015;
  wire _net_3016;
  wire _net_3017;
  wire _net_3018;
  wire _net_3019;
  wire _net_3020;
  wire _net_3021;
  wire _net_3022;
  wire _net_3023;
  wire _net_3024;
  wire _net_3025;
  wire _net_3026;
  wire _net_3027;
  wire _net_3028;
  wire _net_3029;
  wire _net_3030;
  wire _net_3031;
  wire _net_3032;
  wire _net_3033;
  wire _net_3034;
  wire _net_3035;
  wire _net_3036;
  wire _net_3037;
  wire _net_3038;
  wire _net_3039;
  wire _net_3040;
  wire _net_3041;
  wire _net_3042;
  wire _net_3043;
  wire _net_3044;
  wire _net_3045;
  wire _net_3046;
  wire _net_3047;
  wire _net_3048;
  wire _net_3049;
  wire _net_3050;
  wire _net_3051;
  wire _net_3052;
  wire _net_3053;
  wire _net_3054;
  wire _net_3055;
  wire _net_3056;
  wire _net_3057;
  wire _net_3058;
  wire _net_3059;
  wire _net_3060;
  wire _net_3061;
  wire _net_3062;
  wire _net_3063;
  wire _net_3064;
  wire _net_3065;
  wire _net_3066;
  wire _net_3067;
  wire _net_3068;
  wire _net_3069;
  wire _net_3070;
  wire _net_3071;
  wire _net_3072;
  wire _net_3073;
  wire _net_3074;
  wire _net_3075;
  wire _net_3076;
  wire _net_3077;
  wire _net_3078;
  wire _net_3079;
  wire _net_3080;
  wire _net_3081;
  wire _net_3082;
  wire _net_3083;
  wire _net_3084;
  wire _net_3085;
  wire _net_3086;
  wire _net_3087;
  wire _net_3088;
  wire _net_3089;
  wire _net_3090;
  wire _net_3091;
  wire _net_3092;
  wire _net_3093;
  wire _net_3094;
  wire _net_3095;
  wire _net_3096;
  wire _net_3097;
  wire _net_3098;
  wire _net_3099;
  wire _net_3100;
  wire _net_3101;
  wire _net_3102;
  wire _net_3103;
  wire _net_3104;
  wire _net_3105;
  wire _net_3106;
  wire _net_3107;
  wire _net_3108;
  wire _net_3109;
  wire _net_3110;
  wire _net_3111;
  wire _net_3112;
  wire _net_3113;
  wire _net_3114;
  wire _net_3115;
  wire _net_3116;
  wire _net_3117;
  wire _net_3118;
  wire _net_3119;
  wire _net_3120;
  wire _net_3121;
  wire _net_3122;
  wire _net_3123;
  wire _net_3124;
  wire _net_3125;
  wire _net_3126;
  wire _net_3127;
  wire _net_3128;
  wire _net_3129;
  wire _net_3130;
  wire _net_3131;
  wire _net_3132;
  wire _net_3133;
  wire _net_3134;
  wire _net_3135;
  wire _net_3136;
  wire _net_3137;
  wire _net_3138;
  wire _net_3139;
  wire _net_3140;
  wire _net_3141;
  wire _net_3142;
  wire _net_3143;
  wire _net_3144;
  wire _net_3145;
  wire _net_3146;
  wire _net_3147;
  wire _net_3148;
  wire _net_3149;
  wire _net_3150;
  wire _net_3151;
  wire _net_3152;
  wire _net_3153;
  wire _net_3154;
  wire _net_3155;
  wire _net_3156;
  wire _net_3157;
  wire _net_3158;
  wire _net_3159;
  wire _net_3160;
  wire _net_3161;
  wire _net_3162;
  wire _net_3163;
  wire _net_3164;
  wire _net_3165;
  wire _net_3166;
  wire _net_3167;
  wire _net_3168;
  wire _net_3169;
  wire _net_3170;
  wire _net_3171;
  wire _net_3172;
  wire _net_3173;
  wire _net_3174;
  wire _net_3175;
  wire _net_3176;
  wire _net_3177;
  wire _net_3178;
  wire _net_3179;
  wire _net_3180;
  wire _net_3181;
  wire _net_3182;
  wire _net_3183;
  wire _net_3184;
  wire _net_3185;
  wire _net_3186;
  wire _net_3187;
  wire _net_3188;
  wire _net_3189;
  wire _net_3190;
  wire _net_3191;
  wire _net_3192;
  wire _net_3193;
  wire _net_3194;
  wire _net_3195;
  wire _net_3196;
  wire _net_3197;
  wire _net_3198;
  wire _net_3199;
  wire _net_3200;
  wire _net_3201;
  wire _net_3202;
  wire _net_3203;
  wire _net_3204;
  wire _net_3205;
  wire _net_3206;
  wire _net_3207;
  wire _net_3208;
  wire _net_3209;
  wire _net_3210;
  wire _net_3211;
  wire _net_3212;
  wire _net_3213;
  wire _net_3214;
  wire _net_3215;
  wire _net_3216;
  wire _net_3217;
  wire _net_3218;
  wire _net_3219;
  wire _net_3220;
  wire _net_3221;
  wire _net_3222;
  wire _net_3223;
  wire _net_3224;
  wire _net_3225;
  wire _net_3226;
  wire _net_3227;
  wire _net_3228;
  wire _net_3229;
  wire _net_3230;
  wire _net_3231;
  wire _net_3232;
  wire _net_3233;
  wire _net_3234;
  wire _net_3235;
  wire _net_3236;
  wire _net_3237;
  wire _net_3238;
  wire _net_3239;
  wire _net_3240;
  wire _net_3241;
  wire _net_3242;
  wire _net_3243;
  wire _net_3244;
  wire _net_3245;
  wire _net_3246;
  wire _net_3247;
  wire _net_3248;
  wire _net_3249;
  wire _net_3250;
  wire _net_3251;
  wire _net_3252;
  wire _net_3253;
  wire _net_3254;
  wire _net_3255;
  wire _net_3256;
  wire _net_3257;
  wire _net_3258;
  wire _net_3259;
  wire _net_3260;
  wire _net_3261;
  wire _net_3262;
  wire _net_3263;
  wire _net_3264;
  wire _net_3265;
  wire _net_3266;
  wire _net_3267;
  wire _net_3268;
  wire _net_3269;
  wire _net_3270;
  wire _net_3271;
  wire _net_3272;
  wire _net_3273;
  wire _net_3274;
  wire _net_3275;
  wire _net_3276;
  wire _net_3277;
  wire _net_3278;
  wire _net_3279;
  wire _net_3280;
  wire _net_3281;
  wire _net_3282;
  wire _net_3283;
  wire _net_3284;
  wire _net_3285;
  wire _net_3286;
  wire _net_3287;
  wire _net_3288;
  wire _net_3289;
  wire _net_3290;
  wire _net_3291;
  wire _net_3292;
  wire _net_3293;
  wire _net_3294;
  wire _net_3295;
  wire _net_3296;
  wire _net_3297;
  wire _net_3298;
  wire _net_3299;
  wire _net_3300;
  wire _net_3301;
  wire _net_3302;
  wire _net_3303;
  wire _net_3304;
  wire _net_3305;
  wire _net_3306;
  wire _net_3307;
  wire _net_3308;
  wire _net_3309;
  wire _net_3310;
  wire _net_3311;
  wire _net_3312;
  wire _net_3313;
  wire _net_3314;
  wire _net_3315;
  wire _net_3316;
  wire _net_3317;
  wire _net_3318;
  wire _net_3319;
  wire _net_3320;
  wire _net_3321;
  wire _net_3322;
  wire _net_3323;
  wire _net_3324;
  wire _net_3325;
  wire _net_3326;
  wire _net_3327;
  wire _net_3328;
  wire _net_3329;
  wire _net_3330;
  wire _net_3331;
  wire _net_3332;
  wire _net_3333;
  wire _net_3334;
  wire _net_3335;
  wire _net_3336;
  wire _net_3337;
  wire _net_3338;
  wire _net_3339;
  wire _net_3340;
  wire _net_3341;
  wire _net_3342;
  wire _net_3343;
  wire _net_3344;
  wire _net_3345;
  wire _net_3346;
  wire _net_3347;
  wire _net_3348;
  wire _net_3349;
  wire _net_3350;
  wire _net_3351;
  wire _net_3352;
  wire _net_3353;
  wire _net_3354;
  wire _net_3355;
  wire _net_3356;
  wire _net_3357;
  wire _net_3358;
  wire _net_3359;
  wire _net_3360;
  wire _net_3361;
  wire _net_3362;
  wire _net_3363;
  wire _net_3364;
  wire _net_3365;
  wire _net_3366;
  wire _net_3367;
  wire _net_3368;
  wire _net_3369;
  wire _net_3370;
  wire _net_3371;
  wire _net_3372;
  wire _net_3373;
  wire _net_3374;
  wire _net_3375;
  wire _net_3376;
  wire _net_3377;
  wire _net_3378;
  wire _net_3379;
  wire _net_3380;
  wire _net_3381;
  wire _net_3382;
  wire _net_3383;
  wire _net_3384;
  wire _net_3385;
  wire _net_3386;
  wire _net_3387;
  wire _net_3388;
  wire _net_3389;
  wire _net_3390;
  wire _net_3391;
  wire _net_3392;
  wire _net_3393;
  wire _net_3394;
  wire _net_3395;
  wire _net_3396;
  wire _net_3397;
  wire _net_3398;
  wire _net_3399;
  wire _net_3400;
  wire _net_3401;
  wire _net_3402;
  wire _net_3403;
  wire _net_3404;
  wire _net_3405;
  wire _net_3406;
  wire _net_3407;
  wire _net_3408;
  wire _net_3409;
  wire _net_3410;
  wire _net_3411;
  wire _net_3412;
  wire _net_3413;
  wire _net_3414;
  wire _net_3415;
  wire _net_3416;
  wire _net_3417;
  wire _net_3418;
  wire _net_3419;
  wire _net_3420;
  wire _net_3421;
  wire _net_3422;
  wire _net_3423;
  wire _net_3424;
  wire _net_3425;
  wire _net_3426;
  wire _net_3427;
  wire _net_3428;
  wire _net_3429;
  wire _net_3430;
  wire _net_3431;
  wire _net_3432;
  wire _net_3433;
  wire _net_3434;
  wire _net_3435;
  wire _net_3436;
  wire _net_3437;
  wire _net_3438;
  wire _net_3439;
  wire _net_3440;
  wire _net_3441;
  wire _net_3442;
  wire _net_3443;
  wire _net_3444;
  wire _net_3445;
  wire _net_3446;
  wire _net_3447;
  wire _net_3448;
  wire _net_3449;
  wire _net_3450;
  wire _net_3451;
  wire _net_3452;
  wire _net_3453;
  wire _net_3454;
  wire _net_3455;
  wire _net_3456;
  wire _net_3457;
  wire _net_3458;
  wire _net_3459;
  wire _net_3460;
  wire _net_3461;
  wire _net_3462;
  wire _net_3463;
  wire _net_3464;
  wire _net_3465;
  wire _net_3466;
  wire _net_3467;
  wire _net_3468;
  wire _net_3469;
  wire _net_3470;
  wire _net_3471;
  wire _net_3472;
  wire _net_3473;
  wire _net_3474;
  wire _net_3475;
  wire _net_3476;
  wire _net_3477;
  wire _net_3478;
  wire _net_3479;
  wire _net_3480;
  wire _net_3481;
  wire _net_3482;
  wire _net_3483;
  wire _net_3484;
  wire _net_3485;
  wire _net_3486;
  wire _net_3487;
  wire _net_3488;
  wire _net_3489;
  wire _net_3490;
  wire _net_3491;
  wire _net_3492;
  wire _net_3493;
  wire _net_3494;
  wire _net_3495;
  wire _net_3496;
  wire _net_3497;
  wire _net_3498;
  wire _net_3499;
  wire _net_3500;
  wire _net_3501;
  wire _net_3502;
  wire _net_3503;
  wire _net_3504;
  wire _net_3505;
  wire _net_3506;
  wire _net_3507;
  wire _net_3508;
  wire _net_3509;
  wire _net_3510;
  wire _net_3511;
  wire _net_3512;
  wire _net_3513;
  wire _net_3514;
  wire _net_3515;
  wire _net_3516;
  wire _net_3517;
  wire _net_3518;
  wire _net_3519;
  wire _net_3520;
  wire _net_3521;
  wire _net_3522;
  wire _net_3523;
  wire _net_3524;
  wire _net_3525;
  wire _net_3526;
  wire _net_3527;
  wire _net_3528;
  wire _net_3529;
  wire _net_3530;
  wire _net_3531;
  wire _net_3532;
  wire _net_3533;
  wire _net_3534;
  wire _net_3535;
  wire _net_3536;
  wire _net_3537;
  wire _net_3538;
  wire _net_3539;
  wire _net_3540;
  wire _net_3541;
  wire _net_3542;
  wire _net_3543;
  wire _net_3544;
  wire _net_3545;
  wire _net_3546;
  wire _net_3547;
  wire _net_3548;
  wire _net_3549;
  wire _net_3550;
  wire _net_3551;
  wire _net_3552;
  wire _net_3553;
  wire _net_3554;
  wire _net_3555;
  wire _net_3556;
  wire _net_3557;
  wire _net_3558;
  wire _net_3559;
  wire _net_3560;
  wire _net_3561;
  wire _net_3562;
  wire _net_3563;
  wire _net_3564;
  wire _net_3565;
  wire _net_3566;
  wire _net_3567;
  wire _net_3568;
  wire _net_3569;
  wire _net_3570;
  wire _net_3571;
  wire _net_3572;
  wire _net_3573;
  wire _net_3574;
  wire _net_3575;
  wire _net_3576;
  wire _net_3577;
  wire _net_3578;
  wire _net_3579;
  wire _net_3580;
  wire _net_3581;
  wire _net_3582;
  wire _net_3583;
  wire _net_3584;
  wire _net_3585;
  wire _net_3586;
  wire _net_3587;
  wire _net_3588;
  wire _net_3589;
  wire _net_3590;
  wire _net_3591;
  wire _net_3592;
  wire _net_3593;
  wire _net_3594;
  wire _net_3595;
  wire _net_3596;
  wire _net_3597;
  wire _net_3598;
  wire _net_3599;
  wire _net_3600;
  wire _net_3601;
  wire _net_3602;
  wire _net_3603;
  wire _net_3604;
  wire _net_3605;
  wire _net_3606;
  wire _net_3607;
  wire _net_3608;
  wire _net_3609;
  wire _net_3610;
  wire _net_3611;
  wire _net_3612;
  wire _net_3613;
  wire _net_3614;
  wire _net_3615;
  wire _net_3616;
  wire _net_3617;
  wire _net_3618;
  wire _net_3619;
  wire _net_3620;
  wire _net_3621;
  wire _net_3622;
  wire _net_3623;
  wire _net_3624;
  wire _net_3625;
  wire _net_3626;
  wire _net_3627;
  wire _net_3628;
  wire _net_3629;
  wire _net_3630;
  wire _net_3631;
  wire _net_3632;
  wire _net_3633;
  wire _net_3634;
  wire _net_3635;
  wire _net_3636;
  wire _net_3637;
  wire _net_3638;
  wire _net_3639;
  wire _net_3640;
  wire _net_3641;
  wire _net_3642;
  wire _net_3643;
  wire _net_3644;
  wire _net_3645;
  wire _net_3646;
  wire _net_3647;
  wire _net_3648;
  wire _net_3649;
  wire _net_3650;
  wire _net_3651;
  wire _net_3652;
  wire _net_3653;
  wire _net_3654;
  wire _net_3655;
  wire _net_3656;
  wire _net_3657;
  wire _net_3658;
  wire _net_3659;
  wire _net_3660;
  wire _net_3661;
  wire _net_3662;
  wire _net_3663;
  wire _net_3664;
  wire _net_3665;
  wire _net_3666;
  wire _net_3667;
  wire _net_3668;
  wire _net_3669;
  wire _net_3670;
  wire _net_3671;
  wire _net_3672;
  wire _net_3673;
  wire _net_3674;
  wire _net_3675;
  wire _net_3676;
  wire _net_3677;
  wire _net_3678;
  wire _net_3679;
  wire _net_3680;
  wire _net_3681;
  wire _net_3682;
  wire _net_3683;
  wire _net_3684;
  wire _net_3685;
  wire _net_3686;
  wire _net_3687;
  wire _net_3688;
  wire _net_3689;
  wire _net_3690;
  wire _net_3691;
  wire _net_3692;
  wire _net_3693;
  wire _net_3694;
  wire _net_3695;
  wire _net_3696;
  wire _net_3697;
  wire _net_3698;
  wire _net_3699;
  wire _net_3700;
  wire _net_3701;
  wire _net_3702;
  wire _net_3703;
  wire _net_3704;
  wire _net_3705;
  wire _net_3706;
  wire _net_3707;
  wire _net_3708;
  wire _net_3709;
  wire _net_3710;
  wire _net_3711;
  wire _net_3712;
  wire _net_3713;
  wire _net_3714;
  wire _net_3715;
  wire _net_3716;
  wire _net_3717;
  wire _net_3718;
  wire _net_3719;
  wire _net_3720;
  wire _net_3721;
  wire _net_3722;
  wire _net_3723;
  wire _net_3724;
  wire _net_3725;
  wire _net_3726;
  wire _net_3727;
  wire _net_3728;
  wire _net_3729;
  wire _net_3730;
  wire _net_3731;
  wire _net_3732;
  wire _net_3733;
  wire _net_3734;
  wire _net_3735;
  wire _net_3736;
  wire _net_3737;
  wire _net_3738;
  wire _net_3739;
  wire _net_3740;
  wire _net_3741;
  wire _net_3742;
  wire _net_3743;
  wire _net_3744;
  wire _net_3745;
  wire _net_3746;
  wire _net_3747;
  wire _net_3748;
  wire _net_3749;
  wire _net_3750;
  wire _net_3751;
  wire _net_3752;
  wire _net_3753;
  wire _net_3754;
  wire _net_3755;
  wire _net_3756;
  wire _net_3757;
  wire _net_3758;
  wire _net_3759;
  wire _net_3760;
  wire _net_3761;
  wire _net_3762;
  wire _net_3763;
  wire _net_3764;
  wire _net_3765;
  wire _net_3766;
  wire _net_3767;
  wire _net_3768;
  wire _net_3769;
  wire _net_3770;
  wire _net_3771;
  wire _net_3772;
  wire _net_3773;
  wire _net_3774;
  wire _net_3775;
  wire _net_3776;
  wire _net_3777;
  wire _net_3778;
  wire _net_3779;
  wire _net_3780;
  wire _net_3781;
  wire _net_3782;
  wire _net_3783;
  wire _net_3784;
  wire _net_3785;
  wire _net_3786;
  wire _net_3787;
  wire _net_3788;
  wire _net_3789;
  wire _net_3790;
  wire _net_3791;
  wire _net_3792;
  wire _net_3793;
  wire _net_3794;
  wire _net_3795;
  wire _net_3796;
  wire _net_3797;
  wire _net_3798;
  wire _net_3799;
  wire _net_3800;
  wire _net_3801;
  wire _net_3802;
  wire _net_3803;
  wire _net_3804;
  wire _net_3805;
  wire _net_3806;
  wire _net_3807;
  wire _net_3808;
  wire _net_3809;
  wire _net_3810;
  wire _net_3811;
  wire _net_3812;
  wire _net_3813;
  wire _net_3814;
  wire _net_3815;
  wire _net_3816;
  wire _net_3817;
  wire _net_3818;
  wire _net_3819;
  wire _net_3820;
  wire _net_3821;
  wire _net_3822;
  wire _net_3823;
  wire _net_3824;
  wire _net_3825;
  wire _net_3826;
  wire _net_3827;
  wire _net_3828;
  wire _net_3829;
  wire _net_3830;
  wire _net_3831;
  wire _net_3832;
  wire _net_3833;
  wire _net_3834;
  wire _net_3835;
  wire _net_3836;
  wire _net_3837;
  wire _net_3838;
  wire _net_3839;
  wire _net_3840;
  wire _net_3841;
  wire _net_3842;
  wire _net_3843;
  wire _net_3844;
  wire _net_3845;
  wire _net_3846;
  wire _net_3847;
  wire _net_3848;
  wire _net_3849;
  wire _net_3850;
  wire _net_3851;
  wire _net_3852;
  wire _net_3853;
  wire _net_3854;
  wire _net_3855;
  wire _net_3856;
  wire _net_3857;
  wire _net_3858;
  wire _net_3859;
  wire _net_3860;
  wire _net_3861;
  wire _net_3862;
  wire _net_3863;
  wire _net_3864;
  wire _net_3865;
  wire _net_3866;
  wire _net_3867;
  wire _net_3868;
  wire _net_3869;
  wire _net_3870;
  wire _net_3871;
  wire _net_3872;
  wire _net_3873;
  wire _net_3874;
  wire _net_3875;
  wire _net_3876;
  wire _net_3877;
  wire _net_3878;
  wire _net_3879;
  wire _net_3880;
  wire _net_3881;
  wire _net_3882;
  wire _net_3883;
  wire _net_3884;
  wire _net_3885;
  wire _net_3886;
  wire _net_3887;
  wire _net_3888;
  wire _net_3889;
  wire _net_3890;
  wire _net_3891;
  wire _net_3892;
  wire _net_3893;
  wire _net_3894;
  wire _net_3895;
  wire _net_3896;
  wire _net_3897;
  wire _net_3898;
  wire _net_3899;
  wire _net_3900;
  wire _net_3901;
  wire _net_3902;
  wire _net_3903;
  wire _net_3904;
  wire _net_3905;
  wire _net_3906;
  wire _net_3907;
  wire _net_3908;
  wire _net_3909;
  wire _net_3910;
  wire _net_3911;
  wire _net_3912;
  wire _net_3913;
  wire _net_3914;
  wire _net_3915;
  wire _net_3916;
  wire _net_3917;
  wire _net_3918;
  wire _net_3919;
  wire _net_3920;
  wire _net_3921;
  wire _net_3922;
  wire _net_3923;
  wire _net_3924;
  wire _net_3925;
  wire _net_3926;
  wire _net_3927;
  wire _net_3928;
  wire _net_3929;
  wire _net_3930;
  wire _net_3931;
  wire _net_3932;
  wire _net_3933;
  wire _net_3934;
  wire _net_3935;
  wire _net_3936;
  wire _net_3937;
  wire _net_3938;
  wire _net_3939;
  wire _net_3940;
  wire _net_3941;
  wire _net_3942;
  wire _net_3943;
  wire _net_3944;
  wire _net_3945;
  wire _net_3946;
  wire _net_3947;
  wire _net_3948;
  wire _net_3949;
  wire _net_3950;
  wire _net_3951;
  wire _net_3952;
  wire _net_3953;
  wire _net_3954;
  wire _net_3955;
  wire _net_3956;
  wire _net_3957;
  wire _net_3958;
  wire _net_3959;
  wire _net_3960;
  wire _net_3961;
  wire _net_3962;
  wire _net_3963;
  wire _net_3964;
  wire _net_3965;
  wire _net_3966;
  wire _net_3967;
  wire _net_3968;
  wire _net_3969;
  wire _net_3970;
  wire _net_3971;
  wire _net_3972;
  wire _net_3973;
  wire _net_3974;
  wire _net_3975;
  wire _net_3976;
  wire _net_3977;
  wire _net_3978;
  wire _net_3979;
  wire _net_3980;
  wire _net_3981;
  wire _net_3982;
  wire _net_3983;
  wire _net_3984;
  wire _net_3985;
  wire _net_3986;
  wire _net_3987;
  wire _net_3988;
  wire _net_3989;
  wire _net_3990;
  wire _net_3991;
  wire _net_3992;
  wire _net_3993;
  wire _net_3994;
  wire _net_3995;
  wire _net_3996;
  wire _net_3997;
  wire _net_3998;
  wire _net_3999;
  wire _net_4000;
  wire _net_4001;
  wire _net_4002;
  wire _net_4003;
  wire _net_4004;
  wire _net_4005;
  wire _net_4006;
  wire _net_4007;
  wire _net_4008;
  wire _net_4009;
  wire _net_4010;
  wire _net_4011;
  wire _net_4012;
  wire _net_4013;
  wire _net_4014;
  wire _net_4015;
  wire _net_4016;
  wire _net_4017;
  wire _net_4018;
  wire _net_4019;
  wire _net_4020;
  wire _net_4021;
  wire _net_4022;
  wire _net_4023;
  wire _net_4024;
  wire _net_4025;
  wire _net_4026;
  wire _net_4027;
  wire _net_4028;
  wire _net_4029;
  wire _net_4030;
  wire _net_4031;
  wire _net_4032;
  wire _net_4033;
  wire _net_4034;
  wire _net_4035;
  wire _net_4036;
  wire _net_4037;
  wire _net_4038;
  wire _net_4039;
  wire _net_4040;
  wire _net_4041;
  wire _net_4042;
  wire _net_4043;
  wire _net_4044;
  wire _net_4045;
  wire _net_4046;
  wire _net_4047;
  wire _net_4048;
  wire _net_4049;
  wire _net_4050;
  wire _net_4051;
  wire _net_4052;
  wire _net_4053;
  wire _net_4054;
  wire _net_4055;
  wire _net_4056;
  wire _net_4057;
  wire _net_4058;
  wire _net_4059;
  wire _net_4060;
  wire _net_4061;
  wire _net_4062;
  wire _net_4063;
  wire _net_4064;
  wire _net_4065;
  wire _net_4066;
  wire _net_4067;
  wire _net_4068;
  wire _net_4069;
  wire _net_4070;
  wire _net_4071;
  wire _net_4072;
  wire _net_4073;
  wire _net_4074;
  wire _net_4075;
  wire _net_4076;
  wire _net_4077;
  wire _net_4078;
  wire _net_4079;
  wire _net_4080;
  wire _net_4081;
  wire _net_4082;
  wire _net_4083;
  wire _net_4084;
  wire _net_4085;
  wire _net_4086;
  wire _net_4087;
  wire _net_4088;
  wire _net_4089;
  wire _net_4090;
  wire _net_4091;
  wire _net_4092;
  wire _net_4093;
  wire _net_4094;
  wire _net_4095;
  wire _net_4096;
  wire _net_4097;
  wire _net_4098;
  wire _net_4099;
  wire _net_4100;
  wire _net_4101;
  wire _net_4102;
  wire _net_4103;
  wire _net_4104;
  wire _net_4105;
  wire _net_4106;
  wire _net_4107;
  wire _net_4108;
  wire _net_4109;
  wire _net_4110;
  wire _net_4111;
  wire _net_4112;
  wire _net_4113;
  wire _net_4114;
  wire _net_4115;
  wire _net_4116;
  wire _net_4117;
  wire _net_4118;
  wire _net_4119;
  wire _net_4120;
  wire _net_4121;
  wire _net_4122;
  wire _net_4123;
  wire _net_4124;
  wire _net_4125;
  wire _net_4126;
  wire _net_4127;
  wire _net_4128;
  wire _net_4129;
  wire _net_4130;
  wire _net_4131;
  wire _net_4132;
  wire _net_4133;
  wire _net_4134;
  wire _net_4135;
  wire _net_4136;
  wire _net_4137;
  wire _net_4138;
  wire _net_4139;
  wire _net_4140;
  wire _net_4141;
  wire _net_4142;
  wire _net_4143;
  wire _net_4144;
  wire _net_4145;
  wire _net_4146;
  wire _net_4147;
  wire _net_4148;
  wire _net_4149;
  wire _net_4150;
  wire _net_4151;
  wire _net_4152;
  wire _net_4153;
  wire _net_4154;
  wire _net_4155;
  wire _net_4156;
  wire _net_4157;
  wire _net_4158;
  wire _net_4159;
  wire _net_4160;
  wire _net_4161;
  wire _net_4162;
  wire _net_4163;
  wire _net_4164;
  wire _net_4165;
  wire _net_4166;
  wire _net_4167;
  wire _net_4168;
  wire _net_4169;
  wire _net_4170;
  wire _net_4171;
  wire _net_4172;
  wire _net_4173;
  wire _net_4174;
  wire _net_4175;
  wire _net_4176;
  wire _net_4177;
  wire _net_4178;
  wire _net_4179;
  wire _net_4180;
  wire _net_4181;
  wire _net_4182;
  wire _net_4183;
  wire _net_4184;
  wire _net_4185;
  wire _net_4186;
  wire _net_4187;
  wire _net_4188;
  wire _net_4189;
  wire _net_4190;
  wire _net_4191;
  wire _net_4192;
  wire _net_4193;
  wire _net_4194;
  wire _net_4195;
  wire _net_4196;
  wire _net_4197;
  wire _net_4198;
  wire _net_4199;
  wire _net_4200;
  wire _net_4201;
  wire _net_4202;
  wire _net_4203;
  wire _net_4204;
  wire _net_4205;
  wire _net_4206;
  wire _net_4207;
  wire _net_4208;
  wire _net_4209;
  wire _net_4210;
  wire _net_4211;
  wire _net_4212;
  wire _net_4213;
  wire _net_4214;
  wire _net_4215;
  wire _net_4216;
  wire _net_4217;
  wire _net_4218;
  wire _net_4219;
  wire _net_4220;
  wire _net_4221;
  wire _net_4222;
  wire _net_4223;
  wire _net_4224;
  wire _net_4225;
  wire _net_4226;
  wire _net_4227;
  wire _net_4228;
  wire _net_4229;
  wire _net_4230;
  wire _net_4231;
  wire _net_4232;
  wire _net_4233;
  wire _net_4234;
  wire _net_4235;
  wire _net_4236;
  wire _net_4237;
  wire _net_4238;
  wire _net_4239;
  wire _net_4240;
  wire _net_4241;
  wire _net_4242;
  wire _net_4243;
  wire _net_4244;
  wire _net_4245;
  wire _net_4246;
  wire _net_4247;
  wire _net_4248;
  wire _net_4249;
  wire _net_4250;
  wire _net_4251;
  wire _net_4252;
  wire _net_4253;
  wire _net_4254;
  wire _net_4255;
  wire _net_4256;
  wire _net_4257;
  wire _net_4258;
  wire _net_4259;
  wire _net_4260;
  wire _net_4261;
  wire _net_4262;
  wire _net_4263;
  wire _net_4264;
  wire _net_4265;
  wire _net_4266;
  wire _net_4267;
  wire _net_4268;
  wire _net_4269;
  wire _net_4270;
  wire _net_4271;
  wire _net_4272;
  wire _net_4273;
  wire _net_4274;
  wire _net_4275;
  wire _net_4276;
  wire _net_4277;
  wire _net_4278;
  wire _net_4279;
  wire _net_4280;
  wire _net_4281;
  wire _net_4282;
  wire _net_4283;
  wire _net_4284;
  wire _net_4285;
  wire _net_4286;
  wire _net_4287;
  wire _net_4288;
  wire _net_4289;
  wire _net_4290;
  wire _net_4291;
  wire _net_4292;
  wire _net_4293;
  wire _net_4294;
  wire _net_4295;
  wire _net_4296;
  wire _net_4297;
  wire _net_4298;
  wire _net_4299;
  wire _net_4300;
  wire _net_4301;
  wire _net_4302;
  wire _net_4303;
  wire _net_4304;
  wire _net_4305;
  wire _net_4306;
  wire _net_4307;
  wire _net_4308;
  wire _net_4309;
  wire _net_4310;
  wire _net_4311;
  wire _net_4312;
  wire _net_4313;
  wire _net_4314;
  wire _net_4315;
  wire _net_4316;
  wire _net_4317;
  wire _net_4318;
  wire _net_4319;
  wire _net_4320;
  wire _net_4321;
  wire _net_4322;
  wire _net_4323;
  wire _net_4324;
  wire _net_4325;
  wire _net_4326;
  wire _net_4327;
  wire _net_4328;
  wire _net_4329;
  wire _net_4330;
  wire _net_4331;
  wire _net_4332;
  wire _net_4333;
  wire _net_4334;
  wire _net_4335;
  wire _net_4336;
  wire _net_4337;
  wire _net_4338;
  wire _net_4339;
  wire _net_4340;
  wire _net_4341;
  wire _net_4342;
  wire _net_4343;
  wire _net_4344;
  wire _net_4345;
  wire _net_4346;
  wire _net_4347;
  wire _net_4348;
  wire _net_4349;
  wire _net_4350;
  wire _net_4351;
  wire _net_4352;
  wire _net_4353;
  wire _net_4354;
  wire _net_4355;
  wire _net_4356;
  wire _net_4357;
  wire _net_4358;
  wire _net_4359;
  wire _net_4360;
  wire _net_4361;
  wire _net_4362;
  wire _net_4363;
  wire _net_4364;
  wire _net_4365;
  wire _net_4366;
  wire _net_4367;
  wire _net_4368;
  wire _net_4369;
  wire _net_4370;
  wire _net_4371;
  wire _net_4372;
  wire _net_4373;
  wire _net_4374;
  wire _net_4375;
  wire _net_4376;
  wire _net_4377;
  wire _net_4378;
  wire _net_4379;
  wire _net_4380;
  wire _net_4381;
  wire _net_4382;
  wire _net_4383;
  wire _net_4384;
  wire _net_4385;
  wire _net_4386;
  wire _net_4387;
  wire _net_4388;
  wire _net_4389;
  wire _net_4390;
  wire _net_4391;
  wire _net_4392;
  wire _net_4393;
  wire _net_4394;
  wire _net_4395;
  wire _net_4396;
  wire _net_4397;
  wire _net_4398;
  wire _net_4399;
  wire _net_4400;
  wire _net_4401;
  wire _net_4402;
  wire _net_4403;
  wire _net_4404;
  wire _net_4405;
  wire _net_4406;
  wire _net_4407;
  wire _net_4408;
  wire _net_4409;
  wire _net_4410;
  wire _net_4411;
  wire _net_4412;
  wire _net_4413;
  wire _net_4414;
  wire _net_4415;
  wire _net_4416;
  wire _net_4417;
  wire _net_4418;
  wire _net_4419;
  wire _net_4420;
  wire _net_4421;
  wire _net_4422;
  wire _net_4423;
  wire _net_4424;
  wire _net_4425;
  wire _net_4426;
  wire _net_4427;
  wire _net_4428;
  wire _net_4429;
  wire _net_4430;
  wire _net_4431;
  wire _net_4432;
  wire _net_4433;
  wire _net_4434;
  wire _net_4435;
  wire _net_4436;
  wire _net_4437;
  wire _net_4438;
  wire _net_4439;
  wire _net_4440;
  wire _net_4441;
  wire _net_4442;
  wire _net_4443;
  wire _net_4444;
  wire _net_4445;
  wire _net_4446;
  wire _net_4447;
  wire _net_4448;
  wire _net_4449;
  wire _net_4450;
  wire _net_4451;
  wire _net_4452;
  wire _net_4453;
  wire _net_4454;
  wire _net_4455;
  wire _net_4456;
  wire _net_4457;
  wire _net_4458;
  wire _net_4459;
  wire _net_4460;
  wire _net_4461;
  wire _net_4462;
  wire _net_4463;
  wire _net_4464;
  wire _net_4465;
  wire _net_4466;
  wire _net_4467;
  wire _net_4468;
  wire _net_4469;
  wire _net_4470;
  wire _net_4471;
  wire _net_4472;
  wire _net_4473;
  wire _net_4474;
  wire _net_4475;
  wire _net_4476;
  wire _net_4477;
  wire _net_4478;
  wire _net_4479;
  wire _net_4480;
  wire _net_4481;
  wire _net_4482;
  wire _net_4483;
  wire _net_4484;
  wire _net_4485;
  wire _net_4486;
  wire _net_4487;
  wire _net_4488;
  wire _net_4489;
  wire _net_4490;
  wire _net_4491;
  wire _net_4492;
  wire _net_4493;
  wire _net_4494;
  wire _net_4495;
  wire _net_4496;
  wire _net_4497;
  wire _net_4498;
  wire _net_4499;
  wire _net_4500;
  wire _net_4501;
  wire _net_4502;
  wire _net_4503;
  wire _net_4504;
  wire _net_4505;
  wire _net_4506;
  wire _net_4507;
  wire _net_4508;
  wire _net_4509;
  wire _net_4510;
  wire _net_4511;
  wire _net_4512;
  wire _net_4513;
  wire _net_4514;
  wire _net_4515;
  wire _net_4516;
  wire _net_4517;
  wire _net_4518;
  wire _net_4519;
  wire _net_4520;
  wire _net_4521;
  wire _net_4522;
  wire _net_4523;
  wire _net_4524;
  wire _net_4525;
  wire _net_4526;
  wire _net_4527;
  wire _net_4528;
  wire _net_4529;
  wire _net_4530;
  wire _net_4531;
  wire _net_4532;
  wire _net_4533;
  wire _net_4534;
  wire _net_4535;
  wire _net_4536;
  wire _net_4537;
  wire _net_4538;
  wire _net_4539;
  wire _net_4540;
  wire _net_4541;
  wire _net_4542;
  wire _net_4543;
  wire _net_4544;
  wire _net_4545;
  wire _net_4546;
  wire _net_4547;
  wire _net_4548;
  wire _net_4549;
  wire _net_4550;
  wire _net_4551;
  wire _net_4552;
  wire _net_4553;
  wire _net_4554;
  wire _net_4555;
  wire _net_4556;
  wire _net_4557;
  wire _net_4558;
  wire _net_4559;
  wire _net_4560;
  wire _net_4561;
  wire _net_4562;
  wire _net_4563;
  wire _net_4564;
  wire _net_4565;
  wire _net_4566;
  wire _net_4567;
  wire _net_4568;
  wire _net_4569;
  wire _net_4570;
  wire _net_4571;
  wire _net_4572;
  wire _net_4573;
  wire _net_4574;
  wire _net_4575;
  wire _net_4576;
  wire _net_4577;
  wire _net_4578;
  wire _net_4579;
  wire _net_4580;
  wire _net_4581;
  wire _net_4582;
  wire _net_4583;
  wire _net_4584;
  wire _net_4585;
  wire _net_4586;
  wire _net_4587;
  wire _net_4588;
  wire _net_4589;
  wire _net_4590;
  wire _net_4591;
  wire _net_4592;
  wire _net_4593;
  wire _net_4594;
  wire _net_4595;
  wire _net_4596;
  wire _net_4597;
  wire _net_4598;
  wire _net_4599;
  wire _net_4600;
  wire _net_4601;
  wire _net_4602;
  wire _net_4603;
  wire _net_4604;
  wire _net_4605;
  wire _net_4606;
  wire _net_4607;
  wire _net_4608;
  wire _net_4609;
  wire _net_4610;
  wire _net_4611;
  wire _net_4612;
  wire _net_4613;
  wire _net_4614;
  wire _net_4615;
  wire _net_4616;
  wire _net_4617;
  wire _net_4618;
  wire _net_4619;
  wire _net_4620;
  wire _net_4621;
  wire _net_4622;
  wire _net_4623;
  wire _net_4624;
  wire _net_4625;
  wire _net_4626;
  wire _net_4627;
  wire _net_4628;
  wire _net_4629;
  wire _net_4630;
  wire _net_4631;
  wire _net_4632;
  wire _net_4633;
  wire _net_4634;
  wire _net_4635;
  wire _net_4636;
  wire _net_4637;
  wire _net_4638;
  wire _net_4639;
  wire _net_4640;
  wire _net_4641;
  wire _net_4642;
  wire _net_4643;
  wire _net_4644;
  wire _net_4645;
  wire _net_4646;
  wire _net_4647;
  wire _net_4648;
  wire _net_4649;
  wire _net_4650;
  wire _net_4651;
  wire _net_4652;
  wire _net_4653;
  wire _net_4654;
  wire _net_4655;
  wire _net_4656;
  wire _net_4657;
  wire _net_4658;
  wire _net_4659;
  wire _net_4660;
  wire _net_4661;
  wire _net_4662;
  wire _net_4663;
  wire _net_4664;
  wire _net_4665;
  wire _net_4666;
  wire _net_4667;
  wire _net_4668;
  wire _net_4669;
  wire _net_4670;
  wire _net_4671;
  wire _net_4672;
  wire _net_4673;
  wire _net_4674;
  wire _net_4675;
  wire _net_4676;
  wire _net_4677;
  wire _net_4678;
  wire _net_4679;
  wire _net_4680;
  wire _net_4681;
  wire _net_4682;
  wire _net_4683;
  wire _net_4684;
  wire _net_4685;
  wire _net_4686;
  wire _net_4687;
  wire _net_4688;
  wire _net_4689;
  wire _net_4690;
  wire _net_4691;
  wire _net_4692;
  wire _net_4693;
  wire _net_4694;
  wire _net_4695;
  wire _net_4696;
  wire _net_4697;
  wire _net_4698;
  wire _net_4699;
  wire _net_4700;
  wire _net_4701;
  wire _net_4702;
  wire _net_4703;
  wire _net_4704;
  wire _net_4705;
  wire _net_4706;
  wire _net_4707;
  wire _net_4708;
  wire _net_4709;
  wire _net_4710;
  wire _net_4711;
  wire _net_4712;
  wire _net_4713;
  wire _net_4714;
  wire _net_4715;
  wire _net_4716;
  wire _net_4717;
  wire _net_4718;
  wire _net_4719;
  wire _net_4720;
  wire _net_4721;
  wire _net_4722;
  wire _net_4723;
  wire _net_4724;
  wire _net_4725;
  wire _net_4726;
  wire _net_4727;
  wire _net_4728;
  wire _net_4729;
  wire _net_4730;
  wire _net_4731;
  wire _net_4732;
  wire _net_4733;
  wire _net_4734;
  wire _net_4735;
  wire _net_4736;
  wire _net_4737;
  wire _net_4738;
  wire _net_4739;
  wire _net_4740;
  wire _net_4741;
  wire _net_4742;
  wire _net_4743;
  wire _net_4744;
  wire _net_4745;
  wire _net_4746;
  wire _net_4747;
  wire _net_4748;
  wire _net_4749;
  wire _net_4750;
  wire _net_4751;
  wire _net_4752;
  wire _net_4753;
  wire _net_4754;
  wire _net_4755;
  wire _net_4756;
  wire _net_4757;
  wire _net_4758;
  wire _net_4759;
  wire _net_4760;
  wire _net_4761;
  wire _net_4762;
  wire _net_4763;
  wire _net_4764;
  wire _net_4765;
  wire _net_4766;
  wire _net_4767;
  wire _net_4768;
  wire _net_4769;
  wire _net_4770;
  wire _net_4771;
  wire _net_4772;
  wire _net_4773;
  wire _net_4774;
  wire _net_4775;
  wire _net_4776;
  wire _net_4777;
  wire _net_4778;
  wire _net_4779;
  wire _net_4780;
  wire _net_4781;
  wire _net_4782;
  wire _net_4783;
  wire _net_4784;
  wire _net_4785;
  wire _net_4786;
  wire _net_4787;
  wire _net_4788;
  wire _net_4789;
  wire _net_4790;
  wire _net_4791;
  wire _net_4792;
  wire _net_4793;
  wire _net_4794;
  wire _net_4795;
  wire _net_4796;
  wire _net_4797;
  wire _net_4798;
  wire _net_4799;
  wire _net_4800;
  wire _net_4801;
  wire _net_4802;
  wire _net_4803;
  wire _net_4804;
  wire _net_4805;
  wire _net_4806;
  wire _net_4807;
  wire _net_4808;
  wire _net_4809;
  wire _net_4810;
  wire _net_4811;
  wire _net_4812;
  wire _net_4813;
  wire _net_4814;
  wire _net_4815;
  wire _net_4816;
  wire _net_4817;
  wire _net_4818;
  wire _net_4819;
  wire _net_4820;
  wire _net_4821;
  wire _net_4822;
  wire _net_4823;
  wire _net_4824;
  wire _net_4825;
  wire _net_4826;
  wire _net_4827;
  wire _net_4828;
  wire _net_4829;
  wire _net_4830;
  wire _net_4831;
  wire _net_4832;
  wire _net_4833;
  wire _net_4834;
  wire _net_4835;
  wire _net_4836;
  wire _net_4837;
  wire _net_4838;
  wire _net_4839;
  wire _net_4840;
  wire _net_4841;
  wire _net_4842;
  wire _net_4843;
  wire _net_4844;
  wire _net_4845;
  wire _net_4846;
  wire _net_4847;
  wire _net_4848;
  wire _net_4849;
  wire _net_4850;
  wire _net_4851;
  wire _net_4852;
  wire _net_4853;
  wire _net_4854;
  wire _net_4855;
  wire _net_4856;
  wire _net_4857;
  wire _net_4858;
  wire _net_4859;
  wire _net_4860;
  wire _net_4861;
  wire _net_4862;
  wire _net_4863;
  wire _net_4864;
  wire _net_4865;
  wire _net_4866;
  wire _net_4867;
  wire _net_4868;
  wire _net_4869;
  wire _net_4870;
  wire _net_4871;
  wire _net_4872;
  wire _net_4873;
  wire _net_4874;
  wire _net_4875;
  wire _net_4876;
  wire _net_4877;
  wire _net_4878;
  wire _net_4879;
  wire _net_4880;
  wire _net_4881;
  wire _net_4882;
  wire _net_4883;
  wire _net_4884;
  wire _net_4885;
  wire _net_4886;
  wire _net_4887;
  wire _net_4888;
  wire _net_4889;
  wire _net_4890;
  wire _net_4891;
  wire _net_4892;
  wire _net_4893;
  wire _net_4894;
  wire _net_4895;
  wire _net_4896;
  wire _net_4897;
  wire _net_4898;
  wire _net_4899;
  wire _net_4900;
  wire _net_4901;
  wire _net_4902;
  wire _net_4903;
  wire _net_4904;
  wire _net_4905;
  wire _net_4906;
  wire _net_4907;
  wire _net_4908;
  wire _net_4909;
  wire _net_4910;
  wire _net_4911;
  wire _net_4912;
  wire _net_4913;
  wire _net_4914;
  wire _net_4915;
  wire _net_4916;
  wire _net_4917;
  wire _net_4918;
  wire _net_4919;
  wire _net_4920;
  wire _net_4921;
  wire _net_4922;
  wire _net_4923;
  wire _net_4924;
  wire _net_4925;
  wire _net_4926;
  wire _net_4927;
  wire _net_4928;
  wire _net_4929;
  wire _net_4930;
  wire _net_4931;
  wire _net_4932;
  wire _net_4933;
  wire _net_4934;
  wire _net_4935;
  wire _net_4936;
  wire _net_4937;
  wire _net_4938;
  wire _net_4939;
  wire _net_4940;
  wire _net_4941;
  wire _net_4942;
  wire _net_4943;
  wire _net_4944;
  wire _net_4945;
  wire _net_4946;
  wire _net_4947;
  wire _net_4948;
  wire _net_4949;
  wire _net_4950;
  wire _net_4951;
  wire _net_4952;
  wire _net_4953;
  wire _net_4954;
  wire _net_4955;
  wire _net_4956;
  wire _net_4957;
  wire _net_4958;
  wire _net_4959;
  wire _net_4960;
  wire _net_4961;
  wire _net_4962;
  wire _net_4963;
  wire _net_4964;
  wire _net_4965;
  wire _net_4966;
  wire _net_4967;
  wire _net_4968;
  wire _net_4969;
  wire _net_4970;
  wire _net_4971;
  wire _net_4972;
  wire _net_4973;
  wire _net_4974;
  wire _net_4975;
  wire _net_4976;
  wire _net_4977;
  wire _net_4978;
  wire _net_4979;
  wire _net_4980;
  wire _net_4981;
  wire _net_4982;
  wire _net_4983;
  wire _net_4984;
  wire _net_4985;
  wire _net_4986;
  wire _net_4987;
  wire _net_4988;
  wire _net_4989;
  wire _net_4990;
  wire _net_4991;
  wire _net_4992;
  wire _net_4993;
  wire _net_4994;
  wire _net_4995;
  wire _net_4996;
  wire _net_4997;
  wire _net_4998;
  wire _net_4999;
  wire _net_5000;
  wire _net_5001;
  wire _net_5002;
  wire _net_5003;
  wire _net_5004;
  wire _net_5005;
  wire _net_5006;
  wire _net_5007;
  wire _net_5008;
  wire _net_5009;
  wire _net_5010;
  wire _net_5011;
  wire _net_5012;
  wire _net_5013;
  wire _net_5014;
  wire _net_5015;
  wire _net_5016;
  wire _net_5017;
  wire _net_5018;
  wire _net_5019;
  wire _net_5020;
  wire _net_5021;
  wire _net_5022;
  wire _net_5023;
  wire _net_5024;
  wire _net_5025;
  wire _net_5026;
  wire _net_5027;
  wire _net_5028;
  wire _net_5029;
  wire _net_5030;
  wire _net_5031;
  wire _net_5032;
  wire _net_5033;
  wire _net_5034;
  wire _net_5035;
  wire _net_5036;
  wire _net_5037;
  wire _net_5038;
  wire _net_5039;
  wire _net_5040;
  wire _net_5041;
  wire _net_5042;
  wire _net_5043;
  wire _net_5044;
  wire _net_5045;
  wire _net_5046;
  wire _net_5047;
  wire _net_5048;
  wire _net_5049;
  wire _net_5050;
  wire _net_5051;
  wire _net_5052;
  wire _net_5053;
  wire _net_5054;
  wire _net_5055;
  wire _net_5056;
  wire _net_5057;
  wire _net_5058;
  wire _net_5059;
  wire _net_5060;
  wire _net_5061;
  wire _net_5062;
  wire _net_5063;
  wire _net_5064;
  wire _net_5065;
  wire _net_5066;
  wire _net_5067;
  wire _net_5068;
  wire _net_5069;
  wire _net_5070;
  wire _net_5071;
  wire _net_5072;
  wire _net_5073;
  wire _net_5074;
  wire _net_5075;
  wire _net_5076;
  wire _net_5077;
  wire _net_5078;
  wire _net_5079;
  wire _net_5080;
  wire _net_5081;
  wire _net_5082;
  wire _net_5083;
  wire _net_5084;
  wire _net_5085;
  wire _net_5086;
  wire _net_5087;
  wire _net_5088;
  wire _net_5089;
  wire _net_5090;
  wire _net_5091;
  wire _net_5092;
  wire _net_5093;
  wire _net_5094;
  wire _net_5095;
  wire _net_5096;
  wire _net_5097;
  wire _net_5098;
  wire _net_5099;
  wire _net_5100;
  wire _net_5101;
  wire _net_5102;
  wire _net_5103;
  wire _net_5104;
  wire _net_5105;
  wire _net_5106;
  wire _net_5107;
  wire _net_5108;
  wire _net_5109;
  wire _net_5110;
  wire _net_5111;
  wire _net_5112;
  wire _net_5113;
  wire _net_5114;
  wire _net_5115;
  wire _net_5116;
  wire _net_5117;
  wire _net_5118;
  wire _net_5119;
  wire _net_5120;
  wire _net_5121;
  wire _net_5122;
  wire _net_5123;
  wire _net_5124;
  wire _net_5125;
  wire _net_5126;
  wire _net_5127;
  wire _net_5128;
  wire _net_5129;
  wire _net_5130;
  wire _net_5131;
  wire _net_5132;
  wire _net_5133;
  wire _net_5134;
  wire _net_5135;
  wire _net_5136;
  wire _net_5137;
  wire _net_5138;
  wire _net_5139;
  wire _net_5140;
  wire _net_5141;
  wire _net_5142;
  wire _net_5143;
  wire _net_5144;
  wire _net_5145;
  wire _net_5146;
  wire _net_5147;
  wire _net_5148;
  wire _net_5149;
  wire _net_5150;
  wire _net_5151;
  wire _net_5152;
  wire _net_5153;
  wire _net_5154;
  wire _net_5155;
  wire _net_5156;
  wire _net_5157;
  wire _net_5158;
  wire _net_5159;
  wire _net_5160;
  wire _net_5161;
  wire _net_5162;
  wire _net_5163;
  wire _net_5164;
  wire _net_5165;
  wire _net_5166;
  wire _net_5167;
  wire _net_5168;
  wire _net_5169;
  wire _net_5170;
  wire _net_5171;
  wire _net_5172;
  wire _net_5173;
  wire _net_5174;
  wire _net_5175;
  wire _net_5176;
  wire _net_5177;
  wire _net_5178;
  wire _net_5179;
  wire _net_5180;
  wire _net_5181;
  wire _net_5182;
  wire _net_5183;
  wire _net_5184;
  wire _net_5185;
  wire _net_5186;
  wire _net_5187;
  wire _net_5188;
  wire _net_5189;
  wire _net_5190;
  wire _net_5191;
  wire _net_5192;
  wire _net_5193;
  wire _net_5194;
  wire _net_5195;
  wire _net_5196;
  wire _net_5197;
  wire _net_5198;
  wire _net_5199;
  wire _net_5200;
  wire _net_5201;
  wire _net_5202;
  wire _net_5203;
  wire _net_5204;
  wire _net_5205;
  wire _net_5206;
  wire _net_5207;
  wire _net_5208;
  wire _net_5209;
  wire _net_5210;
  wire _net_5211;
  wire _net_5212;
  wire _net_5213;
  wire _net_5214;
  wire _net_5215;
  wire _net_5216;
  wire _net_5217;
  wire _net_5218;
  wire _net_5219;
  wire _net_5220;
  wire _net_5221;
  wire _net_5222;
  wire _net_5223;
  wire _net_5224;
  wire _net_5225;
  wire _net_5226;
  wire _net_5227;
  wire _net_5228;
  wire _net_5229;
  wire _net_5230;
  wire _net_5231;
  wire _net_5232;
  wire _net_5233;
  wire _net_5234;
  wire _net_5235;
  wire _net_5236;
  wire _net_5237;
  wire _net_5238;
  wire _net_5239;
  wire _net_5240;
  wire _net_5241;
  wire _net_5242;
  wire _net_5243;
  wire _net_5244;
  wire _net_5245;
  wire _net_5246;
  wire _net_5247;
  wire _net_5248;
  wire _net_5249;
  wire _net_5250;
  wire _net_5251;
  wire _net_5252;
  wire _net_5253;
  wire _net_5254;
  wire _net_5255;
  wire _net_5256;
  wire _net_5257;
  wire _net_5258;
  wire _net_5259;
  wire _net_5260;
  wire _net_5261;
  wire _net_5262;
  wire _net_5263;
  wire _net_5264;
  wire _net_5265;
  wire _net_5266;
  wire _net_5267;
  wire _net_5268;
  wire _net_5269;
  wire _net_5270;
  wire _net_5271;
  wire _net_5272;
  wire _net_5273;
  wire _net_5274;
  wire _net_5275;
  wire _net_5276;
  wire _net_5277;
  wire _net_5278;
  wire _net_5279;
  wire _net_5280;
  wire _net_5281;
  wire _net_5282;
  wire _net_5283;
  wire _net_5284;
  wire _net_5285;
  wire _net_5286;
  wire _net_5287;
  wire _net_5288;
  wire _net_5289;
  wire _net_5290;
  wire _net_5291;
  wire _net_5292;
  wire _net_5293;
  wire _net_5294;
  wire _net_5295;
  wire _net_5296;
  wire _net_5297;
  wire _net_5298;
  wire _net_5299;
  wire _net_5300;
  wire _net_5301;
  wire _net_5302;
  wire _net_5303;
  wire _net_5304;
  wire _net_5305;
  wire _net_5306;
  wire _net_5307;
  wire _net_5308;
  wire _net_5309;
  wire _net_5310;
  wire _net_5311;
  wire _net_5312;
  wire _net_5313;
  wire _net_5314;
  wire _net_5315;
  wire _net_5316;
  wire _net_5317;
  wire _net_5318;
  wire _net_5319;
  wire _net_5320;
  wire _net_5321;
  wire _net_5322;
  wire _net_5323;
  wire _net_5324;
  wire _net_5325;
  wire _net_5326;
  wire _net_5327;
  wire _net_5328;
  wire _net_5329;
  wire _net_5330;
  wire _net_5331;
  wire _net_5332;
  wire _net_5333;
  wire _net_5334;
  wire _net_5335;
  wire _net_5336;
  wire _net_5337;
  wire _net_5338;
  wire _net_5339;
  wire _net_5340;
  wire _net_5341;
  wire _net_5342;
  wire _net_5343;
  wire _net_5344;
  wire _net_5345;
  wire _net_5346;
  wire _net_5347;
  wire _net_5348;
  wire _net_5349;
  wire _net_5350;
  wire _net_5351;
  wire _net_5352;
  wire _net_5353;
  wire _net_5354;
  wire _net_5355;
  wire _net_5356;
  wire _net_5357;
  wire _net_5358;
  wire _net_5359;
  wire _net_5360;
  wire _net_5361;
  wire _net_5362;
  wire _net_5363;
  wire _net_5364;
  wire _net_5365;
  wire _net_5366;
  wire _net_5367;
  wire _net_5368;
  wire _net_5369;
  wire _net_5370;
  wire _net_5371;
  wire _net_5372;
  wire _net_5373;
  wire _net_5374;
  wire _net_5375;
  wire _net_5376;
  wire _net_5377;
  wire _net_5378;
  wire _net_5379;
  wire _net_5380;
  wire _net_5381;
  wire _net_5382;
  wire _net_5383;
  wire _net_5384;
  wire _net_5385;
  wire _net_5386;
  wire _net_5387;
  wire _net_5388;
  wire _net_5389;
  wire _net_5390;
  wire _net_5391;
  wire _net_5392;
  wire _net_5393;
  wire _net_5394;
  wire _net_5395;
  wire _net_5396;
  wire _net_5397;
  wire _net_5398;
  wire _net_5399;
  wire _net_5400;
  wire _net_5401;
  wire _net_5402;
  wire _net_5403;
  wire _net_5404;
  wire _net_5405;
  wire _net_5406;
  wire _net_5407;
  wire _net_5408;
  wire _net_5409;
  wire _net_5410;
  wire _net_5411;
  wire _net_5412;
  wire _net_5413;
  wire _net_5414;
  wire _net_5415;
  wire _net_5416;
  wire _net_5417;
  wire _net_5418;
  wire _net_5419;
  wire _net_5420;
  wire _net_5421;
  wire _net_5422;
  wire _net_5423;
  wire _net_5424;
  wire _net_5425;
  wire _net_5426;
  wire _net_5427;
  wire _net_5428;
  wire _net_5429;
  wire _net_5430;
  wire _net_5431;
  wire _net_5432;
  wire _net_5433;
  wire _net_5434;
  wire _net_5435;
  wire _net_5436;
  wire _net_5437;
  wire _net_5438;
  wire _net_5439;
  wire _net_5440;
  wire _net_5441;
  wire _net_5442;
  wire _net_5443;
  wire _net_5444;
  wire _net_5445;
  wire _net_5446;
  wire _net_5447;
  wire _net_5448;
  wire _net_5449;
  wire _net_5450;
  wire _net_5451;
  wire _net_5452;
  wire _net_5453;
  wire _net_5454;
  wire _net_5455;
  wire _net_5456;
  wire _net_5457;
  wire _net_5458;
  wire _net_5459;
  wire _net_5460;
  wire _net_5461;
  wire _net_5462;
  wire _net_5463;
  wire _net_5464;
  wire _net_5465;
  wire _net_5466;
  wire _net_5467;
  wire _net_5468;
  wire _net_5469;
  wire _net_5470;
  wire _net_5471;
  wire _net_5472;
  wire _net_5473;
  wire _net_5474;
  wire _net_5475;
  wire _net_5476;
  wire _net_5477;
  wire _net_5478;
  wire _net_5479;
  wire _net_5480;
  wire _net_5481;
  wire _net_5482;
  wire _net_5483;
  wire _net_5484;
  wire _net_5485;
  wire _net_5486;
  wire _net_5487;
  wire _net_5488;
  wire _net_5489;
  wire _net_5490;
  wire _net_5491;
  wire _net_5492;
  wire _net_5493;
  wire _net_5494;
  wire _net_5495;
  wire _net_5496;
  wire _net_5497;
  wire _net_5498;
  wire _net_5499;
  wire _net_5500;
  wire _net_5501;
  wire _net_5502;
  wire _net_5503;
  wire _net_5504;
  wire _net_5505;
  wire _net_5506;
  wire _net_5507;
  wire _net_5508;
  wire _net_5509;
  wire _net_5510;
  wire _net_5511;
  wire _net_5512;
  wire _net_5513;
  wire _net_5514;
  wire _net_5515;
  wire _net_5516;
  wire _net_5517;
  wire _net_5518;
  wire _net_5519;
  wire _net_5520;
  wire _net_5521;
  wire _net_5522;
  wire _net_5523;
  wire _net_5524;
  wire _net_5525;
  wire _net_5526;
  wire _net_5527;
  wire _net_5528;
  wire _net_5529;
  wire _net_5530;
  wire _net_5531;
  wire _net_5532;
  wire _net_5533;
  wire _net_5534;
  wire _net_5535;
  wire _net_5536;
  wire _net_5537;
  wire _net_5538;
  wire _net_5539;
  wire _net_5540;
  wire _net_5541;
  wire _net_5542;
  wire _net_5543;
  wire _net_5544;
  wire _net_5545;
  wire _net_5546;
  wire _net_5547;
  wire _net_5548;
  wire _net_5549;
  wire _net_5550;
  wire _net_5551;
  wire _net_5552;
  wire _net_5553;
  wire _net_5554;
  wire _net_5555;
  wire _net_5556;
  wire _net_5557;
  wire _net_5558;
  wire _net_5559;
  wire _net_5560;
  wire _net_5561;
  wire _net_5562;
  wire _net_5563;
  wire _net_5564;
  wire _net_5565;
  wire _net_5566;
  wire _net_5567;
  wire _net_5568;
  wire _net_5569;
  wire _net_5570;
  wire _net_5571;
  wire _net_5572;
  wire _net_5573;
  wire _net_5574;
  wire _net_5575;
  wire _net_5576;
  wire _net_5577;
  wire _net_5578;
  wire _net_5579;
  wire _net_5580;
  wire _net_5581;
  wire _net_5582;
  wire _net_5583;
  wire _net_5584;
  wire _net_5585;
  wire _net_5586;
  wire _net_5587;
  wire _net_5588;
  wire _net_5589;
  wire _net_5590;
  wire _net_5591;
  wire _net_5592;
  wire _net_5593;
  wire _net_5594;
  wire _net_5595;
  wire _net_5596;
  wire _net_5597;
  wire _net_5598;
  wire _net_5599;
  wire _net_5600;
  wire _net_5601;
  wire _net_5602;
  wire _net_5603;
  wire _net_5604;
  wire _net_5605;
  wire _net_5606;
  wire _net_5607;
  wire _net_5608;
  wire _net_5609;
  wire _net_5610;
  wire _net_5611;
  wire _net_5612;
  wire _net_5613;
  wire _net_5614;
  wire _net_5615;
  wire _net_5616;
  wire _net_5617;
  wire _net_5618;
  wire _net_5619;
  wire _net_5620;
  wire _net_5621;
  wire _net_5622;
  wire _net_5623;
  wire _net_5624;
  wire _net_5625;
  wire _net_5626;
  wire _net_5627;
  wire _net_5628;
  wire _net_5629;
  wire _net_5630;
  wire _net_5631;
  wire _net_5632;
  wire _net_5633;
  wire _net_5634;
  wire _net_5635;
  wire _net_5636;
  wire _net_5637;
  wire _net_5638;
  wire _net_5639;
  wire _net_5640;
  wire _net_5641;
  wire _net_5642;
  wire _net_5643;
  wire _net_5644;
  wire _net_5645;
  wire _net_5646;
  wire _net_5647;
  wire _net_5648;
  wire _net_5649;
  wire _net_5650;
  wire _net_5651;
  wire _net_5652;
  wire _net_5653;
  wire _net_5654;
  wire _net_5655;
  wire _net_5656;
  wire _net_5657;
  wire _net_5658;
  wire _net_5659;
  wire _net_5660;
  wire _net_5661;
  wire _net_5662;
  wire _net_5663;
  wire _net_5664;
  wire _net_5665;
  wire _net_5666;
  wire _net_5667;
  wire _net_5668;
  wire _net_5669;
  wire _net_5670;
  wire _net_5671;
  wire _net_5672;
  wire _net_5673;
  wire _net_5674;
  wire _net_5675;
  wire _net_5676;
  wire _net_5677;
  wire _net_5678;
  wire _net_5679;
  wire _net_5680;
  wire _net_5681;
  wire _net_5682;
  wire _net_5683;
  wire _net_5684;
  wire _net_5685;
  wire _net_5686;
  wire _net_5687;
  wire _net_5688;
  wire _net_5689;
  wire _net_5690;
  wire _net_5691;
  wire _net_5692;
  wire _net_5693;
  wire _net_5694;
  wire _net_5695;
  wire _net_5696;
  wire _net_5697;
  wire _net_5698;
  wire _net_5699;
  wire _net_5700;
  wire _net_5701;
  wire _net_5702;
  wire _net_5703;
  wire _net_5704;
  wire _net_5705;
  wire _net_5706;
  wire _net_5707;
  wire _net_5708;
  wire _net_5709;
  wire _net_5710;
  wire _net_5711;
  wire _net_5712;
  wire _net_5713;
  wire _net_5714;
  wire _net_5715;
  wire _net_5716;
  wire _net_5717;
  wire _net_5718;
  wire _net_5719;
  wire _net_5720;
  wire _net_5721;
  wire _net_5722;
  wire _net_5723;
  wire _net_5724;
  wire _net_5725;
  wire _net_5726;
  wire _net_5727;
  wire _net_5728;
  wire _net_5729;
  wire _net_5730;
  wire _net_5731;
  wire _net_5732;
  wire _net_5733;
  wire _net_5734;
  wire _net_5735;
  wire _net_5736;
  wire _net_5737;
  wire _net_5738;
  wire _net_5739;
  wire _net_5740;
  wire _net_5741;
  wire _net_5742;
  wire _net_5743;
  wire _net_5744;
  wire _net_5745;
  wire _net_5746;
  wire _net_5747;
  wire _net_5748;
  wire _net_5749;
  wire _net_5750;
  wire _net_5751;
  wire _net_5752;
  wire _net_5753;
  wire _net_5754;
  wire _net_5755;
  wire _net_5756;
  wire _net_5757;
  wire _net_5758;
  wire _net_5759;
  wire _net_5760;
  wire _net_5761;
  wire _net_5762;
  wire _net_5763;
  wire _net_5764;
  wire _net_5765;
  wire _net_5766;
  wire _net_5767;
  wire _net_5768;
  wire _net_5769;
  wire _net_5770;
  wire _net_5771;
  wire _net_5772;
  wire _net_5773;
  wire _net_5774;
  wire _net_5775;
  wire _net_5776;
  wire _net_5777;
  wire _net_5778;
  wire _net_5779;
  wire _net_5780;
  wire _net_5781;
  wire _net_5782;
  wire _net_5783;
  wire _net_5784;
  wire _net_5785;
  wire _net_5786;
  wire _net_5787;
  wire _net_5788;
  wire _net_5789;
  wire _net_5790;
  wire _net_5791;
  wire _net_5792;
  wire _net_5793;
  wire _net_5794;
  wire _net_5795;
  wire _net_5796;
  wire _net_5797;
  wire _net_5798;
  wire _net_5799;
  wire _net_5800;
  wire _net_5801;
  wire _net_5802;
  wire _net_5803;
  wire _net_5804;
  wire _net_5805;
  wire _net_5806;
  wire _net_5807;
  wire _net_5808;
  wire _net_5809;
  wire _net_5810;
  wire _net_5811;
  wire _net_5812;
  wire _net_5813;
  wire _net_5814;
  wire _net_5815;
  wire _net_5816;
  wire _net_5817;
  wire _net_5818;
  wire _net_5819;
  wire _net_5820;
  wire _net_5821;
  wire _net_5822;
  wire _net_5823;
  wire _net_5824;
  wire _net_5825;
  wire _net_5826;
  wire _net_5827;
  wire _net_5828;
  wire _net_5829;
  wire _net_5830;
  wire _net_5831;
  wire _net_5832;
  wire _net_5833;
  wire _net_5834;
  wire _net_5835;
  wire _net_5836;
  wire _net_5837;
  wire _net_5838;
  wire _net_5839;
  wire _net_5840;
  wire _net_5841;
  wire _net_5842;
  wire _net_5843;
  wire _net_5844;
  wire _net_5845;
  wire _net_5846;
  wire _net_5847;
  wire _net_5848;
  wire _net_5849;
  wire _net_5850;
  wire _net_5851;
  wire _net_5852;
  wire _net_5853;
  wire _net_5854;
  wire _net_5855;
  wire _net_5856;
  wire _net_5857;
  wire _net_5858;
  wire _net_5859;
  wire _net_5860;
  wire _net_5861;
  wire _net_5862;
  wire _net_5863;
  wire _net_5864;
  wire _net_5865;
  wire _net_5866;
  wire _net_5867;
  wire _net_5868;
  wire _net_5869;
  wire _net_5870;
  wire _net_5871;
  wire _net_5872;
  wire _net_5873;
  wire _net_5874;
  wire _net_5875;
  wire _net_5876;
  wire _net_5877;
  wire _net_5878;
  wire _net_5879;
  wire _net_5880;
  wire _net_5881;
  wire _net_5882;
  wire _net_5883;
  wire _net_5884;
  wire _net_5885;
  wire _net_5886;
  wire _net_5887;
  wire _net_5888;
  wire _net_5889;
  wire _net_5890;
  wire _net_5891;
  wire _net_5892;
  wire _net_5893;
  wire _net_5894;
  wire _net_5895;
  wire _net_5896;
  wire _net_5897;
  wire _net_5898;
  wire _net_5899;
  wire _net_5900;
  wire _net_5901;
  wire _net_5902;
  wire _net_5903;
  wire _net_5904;
  wire _net_5905;
  wire _net_5906;
  wire _net_5907;
  wire _net_5908;
  wire _net_5909;
  wire _net_5910;
  wire _net_5911;
  wire _net_5912;
  wire _net_5913;
  wire _net_5914;
  wire _net_5915;
  wire _net_5916;
  wire _net_5917;
  wire _net_5918;
  wire _net_5919;
  wire _net_5920;
  wire _net_5921;
  wire _net_5922;
  wire _net_5923;
  wire _net_5924;
  wire _net_5925;
  wire _net_5926;
  wire _net_5927;
  wire _net_5928;
  wire _net_5929;
  wire _net_5930;
  wire _net_5931;
  wire _net_5932;
  wire _net_5933;
  wire _net_5934;
  wire _net_5935;
  wire _net_5936;
  wire _net_5937;
  wire _net_5938;
  wire _net_5939;
  wire _net_5940;
  wire _net_5941;
  wire _net_5942;
  wire _net_5943;
  wire _net_5944;
  wire _net_5945;
  wire _net_5946;
  wire _net_5947;
  wire _net_5948;
  wire _net_5949;
  wire _net_5950;
  wire _net_5951;
  wire _net_5952;
  wire _net_5953;
  wire _net_5954;
  wire _net_5955;
  wire _net_5956;
  wire _net_5957;
  wire _net_5958;
  wire _net_5959;
  wire _net_5960;
  wire _net_5961;
  wire _net_5962;
  wire _net_5963;
  wire _net_5964;
  wire _net_5965;
  wire _net_5966;
  wire _net_5967;
  wire _net_5968;
  wire _net_5969;
  wire _net_5970;
  wire _net_5971;
  wire _net_5972;
  wire _net_5973;
  wire _net_5974;
  wire _net_5975;
  wire _net_5976;
  wire _net_5977;
  wire _net_5978;
  wire _net_5979;
  wire _net_5980;
  wire _net_5981;
  wire _net_5982;
  wire _net_5983;
  wire _net_5984;
  wire _net_5985;
  wire _net_5986;
  wire _net_5987;
  wire _net_5988;
  wire _net_5989;
  wire _net_5990;
  wire _net_5991;
  wire _net_5992;
  wire _net_5993;
  wire _net_5994;
  wire _net_5995;
  wire _net_5996;
  wire _net_5997;
  wire _net_5998;
  wire _net_5999;
  wire _net_6000;
  wire _net_6001;
  wire _net_6002;
  wire _net_6003;
  wire _net_6004;
  wire _net_6005;
  wire _net_6006;
  wire _net_6007;
  wire _net_6008;
  wire _net_6009;
  wire _net_6010;
  wire _net_6011;
  wire _net_6012;
  wire _net_6013;
  wire _net_6014;
  wire _net_6015;
  wire _net_6016;
  wire _net_6017;
  wire _net_6018;
  wire _net_6019;
  wire _net_6020;
  wire _net_6021;
  wire _net_6022;
  wire _net_6023;
  wire _net_6024;
  wire _net_6025;
  wire _net_6026;
  wire _net_6027;
  wire _net_6028;
  wire _net_6029;
  wire _net_6030;
  wire _net_6031;
  wire _net_6032;
  wire _net_6033;
  wire _net_6034;
  wire _net_6035;
  wire _net_6036;
  wire _net_6037;
  wire _net_6038;
  wire _net_6039;
  wire _net_6040;
  wire _net_6041;
  wire _net_6042;
  wire _net_6043;
  wire _net_6044;
  wire _net_6045;
  wire _net_6046;
  wire _net_6047;
  wire _net_6048;
  wire _net_6049;
  wire _net_6050;
  wire _net_6051;
  wire _net_6052;
  wire _net_6053;
  wire _net_6054;
  wire _net_6055;
  wire _net_6056;
  wire _net_6057;
  wire _net_6058;
  wire _net_6059;
  wire _net_6060;
  wire _net_6061;
  wire _net_6062;
  wire _net_6063;
  wire _net_6064;
  wire _net_6065;
  wire _net_6066;
  wire _net_6067;
  wire _net_6068;
  wire _net_6069;
  wire _net_6070;
  wire _net_6071;
  wire _net_6072;
  wire _net_6073;
  wire _net_6074;
  wire _net_6075;
  wire _net_6076;
  wire _net_6077;
  wire _net_6078;
  wire _net_6079;
  wire _net_6080;
  wire _net_6081;
  wire _net_6082;
  wire _net_6083;
  wire _net_6084;
  wire _net_6085;
  wire _net_6086;
  wire _net_6087;
  wire _net_6088;
  wire _net_6089;
  wire _net_6090;
  wire _net_6091;
  wire _net_6092;
  wire _net_6093;
  wire _net_6094;
  wire _net_6095;
  wire _net_6096;
  wire _net_6097;
  wire _net_6098;
  wire _net_6099;
  wire _net_6100;
  wire _net_6101;
  wire _net_6102;
  wire _net_6103;
  wire _net_6104;
  wire _net_6105;
  wire _net_6106;
  wire _net_6107;
  wire _net_6108;
  wire _net_6109;
  wire _net_6110;
  wire _net_6111;
  wire _net_6112;
  wire _net_6113;
  wire _net_6114;
  wire _net_6115;
  wire _net_6116;
  wire _net_6117;
  wire _net_6118;
  wire _net_6119;
  wire _net_6120;
  wire _net_6121;
  wire _net_6122;
  wire _net_6123;
  wire _net_6124;
  wire _net_6125;
  wire _net_6126;
  wire _net_6127;
  wire _net_6128;
  wire _net_6129;
  wire _net_6130;
  wire _net_6131;
  wire _net_6132;
  wire _net_6133;
  wire _net_6134;
  wire _net_6135;
  wire _net_6136;
  wire _net_6137;
  wire _net_6138;
  wire _net_6139;
  wire _net_6140;
  wire _net_6141;
  wire _net_6142;
  wire _net_6143;
  wire _net_6144;
  wire _net_6145;
  wire _net_6146;
  wire _net_6147;
  wire _net_6148;
  wire _net_6149;
  wire _net_6150;
  wire _net_6151;
  wire _net_6152;
  wire _net_6153;
  wire _net_6154;
  wire _net_6155;
  wire _net_6156;
  wire _net_6157;
  wire _net_6158;
  wire _net_6159;
  wire _net_6160;
  wire _net_6161;
  wire _net_6162;
  wire _net_6163;
  wire _net_6164;
  wire _net_6165;
  wire _net_6166;
  wire _net_6167;
  wire _net_6168;
  wire _net_6169;
  wire _net_6170;
  wire _net_6171;
  wire _net_6172;
  wire _net_6173;
  wire _net_6174;
  wire _net_6175;
  wire _net_6176;
  wire _net_6177;
  wire _net_6178;
  wire _net_6179;
  wire _net_6180;
  wire _net_6181;
  wire _net_6182;
  wire _net_6183;
  wire _net_6184;
  wire _net_6185;
  wire _net_6186;
  wire _net_6187;
  wire _net_6188;
  wire _net_6189;
  wire _net_6190;
  wire _net_6191;
  wire _net_6192;
  wire _net_6193;
  wire _net_6194;
  wire _net_6195;
  wire _net_6196;
  wire _net_6197;
  wire _net_6198;
  wire _net_6199;
  wire _net_6200;
  wire _net_6201;
  wire _net_6202;
  wire _net_6203;
  wire _net_6204;
  wire _net_6205;
  wire _net_6206;
  wire _net_6207;
  wire _net_6208;
  wire _net_6209;
  wire _net_6210;
  wire _net_6211;
  wire _net_6212;
  wire _net_6213;
  wire _net_6214;
  wire _net_6215;
  wire _net_6216;
  wire _net_6217;
  wire _net_6218;
  wire _net_6219;
  wire _net_6220;
  wire _net_6221;
  wire _net_6222;
  wire _net_6223;
  wire _net_6224;
  wire _net_6225;
  wire _net_6226;
  wire _net_6227;
  wire _net_6228;
  wire _net_6229;
  wire _net_6230;
  wire _net_6231;
  wire _net_6232;
  wire _net_6233;
  wire _net_6234;
  wire _net_6235;
  wire _net_6236;
  wire _net_6237;
  wire _net_6238;
  wire _net_6239;
  wire _net_6240;
  wire _net_6241;
  wire _net_6242;
  wire _net_6243;
  wire _net_6244;
  wire _net_6245;
  wire _net_6246;
  wire _net_6247;
  wire _net_6248;
  wire _net_6249;
  wire _net_6250;
  wire _net_6251;
  wire _net_6252;
  wire _net_6253;
  wire _net_6254;
  wire _net_6255;
  wire _net_6256;
  wire _net_6257;
  wire _net_6258;
  wire _net_6259;
  wire _net_6260;
  wire _net_6261;
  wire _net_6262;
  wire _net_6263;
  wire _net_6264;
  wire _net_6265;
  wire _net_6266;
  wire _net_6267;
  wire _net_6268;
  wire _net_6269;
  wire _net_6270;
  wire _net_6271;
  wire _net_6272;
  wire _net_6273;
  wire _net_6274;
  wire _net_6275;
  wire _net_6276;
  wire _net_6277;
  wire _net_6278;
  wire _net_6279;
  wire _net_6280;
  wire _net_6281;
  wire _net_6282;
  wire _net_6283;
  wire _net_6284;
  wire _net_6285;
  wire _net_6286;
  wire _net_6287;
  wire _net_6288;
  wire _net_6289;
  wire _net_6290;
  wire _net_6291;
  wire _net_6292;
  wire _net_6293;
  wire _net_6294;
  wire _net_6295;
  wire _net_6296;
  wire _net_6297;
  wire _net_6298;
  wire _net_6299;
  wire _net_6300;
  wire _net_6301;
  wire _net_6302;
  wire _net_6303;
  wire _net_6304;
  wire _net_6305;
  wire _net_6306;
  wire _net_6307;
  wire _net_6308;
  wire _net_6309;
  wire _net_6310;
  wire _net_6311;
  wire _net_6312;
  wire _net_6313;
  wire _net_6314;
  wire _net_6315;
  wire _net_6316;
  wire _net_6317;
  wire _net_6318;
  wire _net_6319;
  wire _net_6320;
  wire _net_6321;
  wire _net_6322;
  wire _net_6323;
  wire _net_6324;
  wire _net_6325;
  wire _net_6326;
  wire _net_6327;
  wire _net_6328;
  wire _net_6329;
  wire _net_6330;
  wire _net_6331;
  wire _net_6332;
  wire _net_6333;
  wire _net_6334;
  wire _net_6335;
  wire _net_6336;
  wire _net_6337;
  wire _net_6338;
  wire _net_6339;
  wire _net_6340;
  wire _net_6341;
  wire _net_6342;
  wire _net_6343;
  wire _net_6344;
  wire _net_6345;
  wire _net_6346;
  wire _net_6347;
  wire _net_6348;
  wire _net_6349;
  wire _net_6350;
  wire _net_6351;
  wire _net_6352;
  wire _net_6353;
  wire _net_6354;
  wire _net_6355;
  wire _net_6356;
  wire _net_6357;
  wire _net_6358;
  wire _net_6359;
  wire _net_6360;
  wire _net_6361;
  wire _net_6362;
  wire _net_6363;
  wire _net_6364;
  wire _net_6365;
  wire _net_6366;
  wire _net_6367;
  wire _net_6368;
  wire _net_6369;
  wire _net_6370;
  wire _net_6371;
  wire _net_6372;
  wire _net_6373;
  wire _net_6374;
  wire _net_6375;
  wire _net_6376;
  wire _net_6377;
  wire _net_6378;
  wire _net_6379;
  wire _net_6380;
  wire _net_6381;
  wire _net_6382;
  wire _net_6383;
  wire _net_6384;
  wire _net_6385;
  wire _net_6386;
  wire _net_6387;
  wire _net_6388;
  wire _net_6389;
  wire _net_6390;
  wire _net_6391;
  wire _net_6392;
  wire _net_6393;
  wire _net_6394;
  wire _net_6395;
  wire _net_6396;
  wire _net_6397;
  wire _net_6398;
  wire _net_6399;
  wire _net_6400;
  wire _net_6401;
  wire _net_6402;
  wire _net_6403;
  wire _net_6404;
  wire _net_6405;
  wire _net_6406;
  wire _net_6407;
  wire _net_6408;
  wire _net_6409;
  wire _net_6410;
  wire _net_6411;
  wire _net_6412;
  wire _net_6413;
  wire _net_6414;
  wire _net_6415;
  wire _net_6416;
  wire _net_6417;
  wire _net_6418;
  wire _net_6419;
  wire _net_6420;
  wire _net_6421;
  wire _net_6422;
  wire _net_6423;
  wire _net_6424;
  wire _net_6425;
  wire _net_6426;
  wire _net_6427;
  wire _net_6428;
  wire _net_6429;
  wire _net_6430;
  wire _net_6431;
  wire _net_6432;
  wire _net_6433;
  wire _net_6434;
  wire _net_6435;
  wire _net_6436;
  wire _net_6437;
  wire _net_6438;
  wire _net_6439;
  wire _net_6440;
  wire _net_6441;
  wire _net_6442;
  wire _net_6443;
  wire _net_6444;
  wire _net_6445;
  wire _net_6446;
  wire _net_6447;
  wire _net_6448;
  wire _net_6449;
  wire _net_6450;
  wire _net_6451;
  wire _net_6452;
  wire _net_6453;
  wire _net_6454;
  wire _net_6455;
  wire _net_6456;
  wire _net_6457;
  wire _net_6458;
  wire _net_6459;
  wire _net_6460;
  wire _net_6461;
  wire _net_6462;
  wire _net_6463;
  wire _net_6464;
  wire _net_6465;
  wire _net_6466;
  wire _net_6467;
  wire _net_6468;
  wire _net_6469;
  wire _net_6470;
  wire _net_6471;
  wire _net_6472;
  wire _net_6473;
  wire _net_6474;
  wire _net_6475;
  wire _net_6476;
  wire _net_6477;
  wire _net_6478;
  wire _net_6479;
  wire _net_6480;
  wire _net_6481;
  wire _net_6482;
  wire _net_6483;
  wire _net_6484;
  wire _net_6485;
  wire _net_6486;
  wire _net_6487;
  wire _net_6488;
  wire _net_6489;
  wire _net_6490;
  wire _net_6491;
  wire _net_6492;
  wire _net_6493;
  wire _net_6494;
  wire _net_6495;
  wire _net_6496;
  wire _net_6497;
  wire _net_6498;
  wire _net_6499;
  wire _net_6500;
  wire _net_6501;
  wire _net_6502;
  wire _net_6503;
  wire _net_6504;
  wire _net_6505;
  wire _net_6506;
  wire _net_6507;
  wire _net_6508;
  wire _net_6509;
  wire _net_6510;
  wire _net_6511;
  wire _net_6512;
  wire _net_6513;
  wire _net_6514;
  wire _net_6515;
  wire _net_6516;
  wire _net_6517;
  wire _net_6518;
  wire _net_6519;
  wire _net_6520;
  wire _net_6521;
  wire _net_6522;
  wire _net_6523;
  wire _net_6524;
  wire _net_6525;
  wire _net_6526;
  wire _net_6527;
  wire _net_6528;
  wire _net_6529;
  wire _net_6530;
  wire _net_6531;
  wire _net_6532;
  wire _net_6533;
  wire _net_6534;
  wire _net_6535;
  wire _net_6536;
  wire _net_6537;
  wire _net_6538;
  wire _net_6539;
  wire _net_6540;
  wire _net_6541;
  wire _net_6542;
  wire _net_6543;
  wire _net_6544;
  wire _net_6545;
  wire _net_6546;
  wire _net_6547;
  wire _net_6548;
  wire _net_6549;
  wire _net_6550;
  wire _net_6551;
  wire _net_6552;
  wire _net_6553;
  wire _net_6554;
  wire _net_6555;
  wire _net_6556;
  wire _net_6557;
  wire _net_6558;
  wire _net_6559;
  wire _net_6560;
  wire _net_6561;
  wire _net_6562;
  wire _net_6563;
  wire _net_6564;
  wire _net_6565;
  wire _net_6566;
  wire _net_6567;
  wire _net_6568;
  wire _net_6569;
  wire _net_6570;
  wire _net_6571;
  wire _net_6572;
  wire _net_6573;
  wire _net_6574;
  wire _net_6575;
  wire _net_6576;
  wire _net_6577;
  wire _net_6578;
  wire _net_6579;
  wire _net_6580;
  wire _net_6581;
  wire _net_6582;
  wire _net_6583;
  wire _net_6584;
  wire _net_6585;
  wire _net_6586;
  wire _net_6587;
  wire _net_6588;
  wire _net_6589;
  wire _net_6590;
  wire _net_6591;
  wire _net_6592;
  wire _net_6593;
  wire _net_6594;
  wire _net_6595;
  wire _net_6596;
  wire _net_6597;
  wire _net_6598;
  wire _net_6599;
  wire _net_6600;
  wire _net_6601;
  wire _net_6602;
  wire _net_6603;
  wire _net_6604;
  wire _net_6605;
  wire _net_6606;
  wire _net_6607;
  wire _net_6608;
  wire _net_6609;
  wire _net_6610;
  wire _net_6611;
  wire _net_6612;
  wire _net_6613;
  wire _net_6614;
  wire _net_6615;
  wire _net_6616;
  wire _net_6617;
  wire _net_6618;
  wire _net_6619;
  wire _net_6620;
  wire _net_6621;
  wire _net_6622;
  wire _net_6623;
  wire _net_6624;
  wire _net_6625;
  wire _net_6626;
  wire _net_6627;
  wire _net_6628;
  wire _net_6629;
  wire _net_6630;
  wire _net_6631;
  wire _net_6632;
  wire _net_6633;
  wire _net_6634;
  wire _net_6635;
  wire _net_6636;
  wire _net_6637;
  wire _net_6638;
  wire _net_6639;
  wire _net_6640;
  wire _net_6641;
  wire _net_6642;
  wire _net_6643;
  wire _net_6644;
  wire _net_6645;
  wire _net_6646;
  wire _net_6647;
  wire _net_6648;
  wire _net_6649;
  wire _net_6650;
  wire _net_6651;
  wire _net_6652;
  wire _net_6653;
  wire _net_6654;
  wire _net_6655;
  wire _net_6656;
  wire _net_6657;
  wire _net_6658;
  wire _net_6659;
  wire _net_6660;
  wire _net_6661;
  wire _net_6662;
  wire _net_6663;
  wire _net_6664;
  wire _net_6665;
  wire _net_6666;
  wire _net_6667;
  wire _net_6668;
  wire _net_6669;
  wire _net_6670;
  wire _net_6671;
  wire _net_6672;
  wire _net_6673;
  wire _net_6674;
  wire _net_6675;
  wire _net_6676;
  wire _net_6677;
  wire _net_6678;
  wire _net_6679;
  wire _net_6680;
  wire _net_6681;
  wire _net_6682;
  wire _net_6683;
  wire _net_6684;
  wire _net_6685;
  wire _net_6686;
  wire _net_6687;
  wire _net_6688;
  wire _net_6689;
  wire _net_6690;
  wire _net_6691;
  wire _net_6692;
  wire _net_6693;
  wire _net_6694;
  wire _net_6695;
  wire _net_6696;
  wire _net_6697;
  wire _net_6698;
  wire _net_6699;
  wire _net_6700;
  wire _net_6701;
  wire _net_6702;
  wire _net_6703;
  wire _net_6704;
  wire _net_6705;
  wire _net_6706;
  wire _net_6707;
  wire _net_6708;
  wire _net_6709;
  wire _net_6710;
  wire _net_6711;
  wire _net_6712;
  wire _net_6713;
  wire _net_6714;
  wire _net_6715;
  wire _net_6716;
  wire _net_6717;
  wire _net_6718;
  wire _net_6719;
  wire _net_6720;
  wire _net_6721;
  wire _net_6722;
  wire _net_6723;
  wire _net_6724;
  wire _net_6725;
  wire _net_6726;
  wire _net_6727;
  wire _net_6728;
  wire _net_6729;
  wire _net_6730;
  wire _net_6731;
  wire _net_6732;
  wire _net_6733;
  wire _net_6734;
  wire _net_6735;
  wire _net_6736;
  wire _net_6737;
  wire _net_6738;
  wire _net_6739;
  wire _net_6740;
  wire _net_6741;
  wire _net_6742;
  wire _net_6743;
  wire _net_6744;
  wire _net_6745;
  wire _net_6746;
  wire _net_6747;
  wire _net_6748;
  wire _net_6749;
  wire _net_6750;
  wire _net_6751;
  wire _net_6752;
  wire _net_6753;
  wire _net_6754;
  wire _net_6755;
  wire _net_6756;
  wire _net_6757;
  wire _net_6758;
  wire _net_6759;
  wire _net_6760;
  wire _net_6761;
  wire _net_6762;
  wire _net_6763;
  wire _net_6764;
  wire _net_6765;
  wire _net_6766;
  wire _net_6767;
  wire _net_6768;
  wire _net_6769;
  wire _net_6770;
  wire _net_6771;
  wire _net_6772;
  wire _net_6773;
  wire _net_6774;
  wire _net_6775;
  wire _net_6776;
  wire _net_6777;
  wire _net_6778;
  wire _net_6779;
  wire _net_6780;
  wire _net_6781;
  wire _net_6782;
  wire _net_6783;
  wire _net_6784;
  wire _net_6785;
  wire _net_6786;
  wire _net_6787;
  wire _net_6788;
  wire _net_6789;
  wire _net_6790;
  wire _net_6791;
  wire _net_6792;
  wire _net_6793;
  wire _net_6794;
  wire _net_6795;
  wire _net_6796;
  wire _net_6797;
  wire _net_6798;
  wire _net_6799;
  wire _net_6800;
  wire _net_6801;
  wire _net_6802;
  wire _net_6803;
  wire _net_6804;
  wire _net_6805;
  wire _net_6806;
  wire _net_6807;
  wire _net_6808;
  wire _net_6809;
  wire _net_6810;
  wire _net_6811;
  wire _net_6812;
  wire _net_6813;
  wire _net_6814;
  wire _net_6815;
  wire _net_6816;
  wire _net_6817;
  wire _net_6818;
  wire _net_6819;
  wire _net_6820;
  wire _net_6821;
  wire _net_6822;
  wire _net_6823;
  wire _net_6824;
  wire _net_6825;
  wire _net_6826;
  wire _net_6827;
  wire _net_6828;
  wire _net_6829;
  wire _net_6830;
  wire _net_6831;
  wire _net_6832;
  wire _net_6833;
  wire _net_6834;
  wire _net_6835;
  wire _net_6836;
  wire _net_6837;
  wire _net_6838;
  wire _net_6839;
  wire _net_6840;
  wire _net_6841;
  wire _net_6842;
  wire _net_6843;
  wire _net_6844;
  wire _net_6845;
  wire _net_6846;
  wire _net_6847;
  wire _net_6848;
  wire _net_6849;
  wire _net_6850;
  wire _net_6851;
  wire _net_6852;
  wire _net_6853;
  wire _net_6854;
  wire _net_6855;
  wire _net_6856;
  wire _net_6857;
  wire _net_6858;
  wire _net_6859;
  wire _net_6860;
  wire _net_6861;
  wire _net_6862;
  wire _net_6863;
  wire _net_6864;
  wire _net_6865;
  wire _net_6866;
  wire _net_6867;
  wire _net_6868;
  wire _net_6869;
  wire _net_6870;
  wire _net_6871;
  wire _net_6872;
  wire _net_6873;
  wire _net_6874;
  wire _net_6875;
  wire _net_6876;
  wire _net_6877;
  wire _net_6878;
  wire _net_6879;
  wire _net_6880;
  wire _net_6881;
  wire _net_6882;
  wire _net_6883;
  wire _net_6884;
  wire _net_6885;
  wire _net_6886;
  wire _net_6887;
  wire _net_6888;
  wire _net_6889;
  wire _net_6890;
  wire _net_6891;
  wire _net_6892;
  wire _net_6893;
  wire _net_6894;
  wire _net_6895;
  wire _net_6896;
  wire _net_6897;
  wire _net_6898;
  wire _net_6899;
  wire _net_6900;
  wire _net_6901;
  wire _net_6902;
  wire _net_6903;
  wire _net_6904;
  wire _net_6905;
  wire _net_6906;
  wire _net_6907;
  wire _net_6908;
  wire _net_6909;
  wire _net_6910;
  wire _net_6911;
  wire _net_6912;
  wire _net_6913;
  wire _net_6914;
  wire _net_6915;
  wire _net_6916;
  wire _net_6917;
  wire _net_6918;
  wire _net_6919;
  wire _net_6920;
  wire _net_6921;
  wire _net_6922;
  wire _net_6923;
  wire _net_6924;
  wire _net_6925;
  wire _net_6926;
  wire _net_6927;
  wire _net_6928;
  wire _net_6929;
  wire _net_6930;
  wire _net_6931;
  wire _net_6932;
  wire _net_6933;
  wire _net_6934;
  wire _net_6935;
  wire _net_6936;
  wire _net_6937;
  wire _net_6938;
  wire _net_6939;
  wire _net_6940;
  wire _net_6941;
  wire _net_6942;
  wire _net_6943;
  wire _net_6944;
  wire _net_6945;
  wire _net_6946;
  wire _net_6947;
  wire _net_6948;
  wire _net_6949;
  wire _net_6950;
  wire _net_6951;
  wire _net_6952;
  wire _net_6953;
  wire _net_6954;
  wire _net_6955;
  wire _net_6956;
  wire _net_6957;
  wire _net_6958;
  wire _net_6959;
  wire _net_6960;
  wire _net_6961;
  wire _net_6962;
  wire _net_6963;
  wire _net_6964;
  wire _net_6965;
  wire _net_6966;
  wire _net_6967;
  wire _net_6968;
  wire _net_6969;
  wire _net_6970;
  wire _net_6971;
  wire _net_6972;
  wire _net_6973;
  wire _net_6974;
  wire _net_6975;
  wire _net_6976;
  wire _net_6977;
  wire _net_6978;
  wire _net_6979;
  wire _net_6980;
  wire _net_6981;
  wire _net_6982;
  wire _net_6983;
  wire _net_6984;
  wire _net_6985;
  wire _net_6986;
  wire _net_6987;
  wire _net_6988;
  wire _net_6989;
  wire _net_6990;
  wire _net_6991;
  wire _net_6992;
  wire _net_6993;
  wire _net_6994;
  wire _net_6995;
  wire _net_6996;
  wire _net_6997;
  wire _net_6998;
  wire _net_6999;
  wire _net_7000;
  wire _net_7001;
  wire _net_7002;
  wire _net_7003;
  wire _net_7004;
  wire _net_7005;
  wire _net_7006;
  wire _net_7007;
  wire _net_7008;
  wire _net_7009;
  wire _net_7010;
  wire _net_7011;
  wire _net_7012;
  wire _net_7013;
  wire _net_7014;
  wire _net_7015;
  wire _net_7016;
  wire _net_7017;
  wire _net_7018;
  wire _net_7019;
  wire _net_7020;
  wire _net_7021;
  wire _net_7022;
  wire _net_7023;
  wire _net_7024;
  wire _net_7025;
  wire _net_7026;
  wire _net_7027;
  wire _net_7028;
  wire _net_7029;
  wire _net_7030;
  wire _net_7031;
  wire _net_7032;
  wire _net_7033;
  wire _net_7034;
  wire _net_7035;
  wire _net_7036;
  wire _net_7037;
  wire _net_7038;
  wire _net_7039;
  wire _net_7040;
  wire _net_7041;
  wire _net_7042;
  wire _net_7043;
  wire _net_7044;
  wire _net_7045;
  wire _net_7046;
  wire _net_7047;
  wire _net_7048;
  wire _net_7049;
  wire _net_7050;
  wire _net_7051;
  wire _net_7052;
  wire _net_7053;
  wire _net_7054;
  wire _net_7055;
  wire _net_7056;
  wire _net_7057;
  wire _net_7058;
  wire _net_7059;
  wire _net_7060;
  wire _net_7061;
  wire _net_7062;
  wire _net_7063;
  wire _net_7064;
  wire _net_7065;
  wire _net_7066;
  wire _net_7067;
  wire _net_7068;
  wire _net_7069;
  wire _net_7070;
  wire _net_7071;
  wire _net_7072;
  wire _net_7073;
  wire _net_7074;
  wire _net_7075;
  wire _net_7076;
  wire _net_7077;
  wire _net_7078;
  wire _net_7079;
  wire _net_7080;
  wire _net_7081;
  wire _net_7082;
  wire _net_7083;
  wire _net_7084;
  wire _net_7085;
  wire _net_7086;
  wire _net_7087;
  wire _net_7088;
  wire _net_7089;
  wire _net_7090;
  wire _net_7091;
  wire _net_7092;
  wire _net_7093;
  wire _net_7094;
  wire _net_7095;
  wire _net_7096;
  wire _net_7097;
  wire _net_7098;
  wire _net_7099;
  wire _net_7100;
  wire _net_7101;
  wire _net_7102;
  wire _net_7103;
  wire _net_7104;
  wire _net_7105;
  wire _net_7106;
  wire _net_7107;
  wire _net_7108;
  wire _net_7109;
  wire _net_7110;
  wire _net_7111;
  wire _net_7112;
  wire _net_7113;
  wire _net_7114;
  wire _net_7115;
  wire _net_7116;
  wire _net_7117;
  wire _net_7118;
  wire _net_7119;
  wire _net_7120;
  wire _net_7121;
  wire _net_7122;
  wire _net_7123;
  wire _net_7124;
  wire _net_7125;
  wire _net_7126;
  wire _net_7127;
  wire _net_7128;
  wire _net_7129;
  wire _net_7130;
  wire _net_7131;
  wire _net_7132;
  wire _net_7133;
  wire _net_7134;
  wire _net_7135;
  wire _net_7136;
  wire _net_7137;
  wire _net_7138;
  wire _net_7139;
  wire _net_7140;
  wire _net_7141;
  wire _net_7142;
  wire _net_7143;
  wire _net_7144;
  wire _net_7145;
  wire _net_7146;
  wire _net_7147;
  wire _net_7148;
  wire _net_7149;
  wire _net_7150;
  wire _net_7151;
  wire _net_7152;
  wire _net_7153;
  wire _net_7154;
  wire _net_7155;
  wire _net_7156;
  wire _net_7157;
  wire _net_7158;
  wire _net_7159;
  wire _net_7160;
  wire _net_7161;
  wire _net_7162;
  wire _net_7163;
  wire _net_7164;
  wire _net_7165;
  wire _net_7166;
  wire _net_7167;
  wire _net_7168;
  wire _net_7169;
  wire _net_7170;
  wire _net_7171;
  wire _net_7172;
  wire _net_7173;
  wire _net_7174;
  wire _net_7175;
  wire _net_7176;
  wire _net_7177;
  wire _net_7178;
  wire _net_7179;
  wire _net_7180;
  wire _net_7181;
  wire _net_7182;
  wire _net_7183;
  wire _net_7184;
  wire _net_7185;
  wire _net_7186;
  wire _net_7187;
  wire _net_7188;
  wire _net_7189;
  wire _net_7190;
  wire _net_7191;
  wire _net_7192;
  wire _net_7193;
  wire _net_7194;
  wire _net_7195;
  wire _net_7196;
  wire _net_7197;
  wire _net_7198;
  wire _net_7199;
  wire _net_7200;
  wire _net_7201;
  wire _net_7202;
  wire _net_7203;
  wire _net_7204;
  wire _net_7205;
  wire _net_7206;
  wire _net_7207;
  wire _net_7208;
  wire _net_7209;
  wire _net_7210;
  wire _net_7211;
  wire _net_7212;
  wire _net_7213;
  wire _net_7214;
  wire _net_7215;
  wire _net_7216;
  wire _net_7217;
  wire _net_7218;
  wire _net_7219;
  wire _net_7220;
  wire _net_7221;
  wire _net_7222;
  wire _net_7223;
  wire _net_7224;
  wire _net_7225;
  wire _net_7226;
  wire _net_7227;
  wire _net_7228;
  wire _net_7229;
  wire _net_7230;
  wire _net_7231;
  wire _net_7232;
  wire _net_7233;
  wire _net_7234;
  wire _net_7235;
  wire _net_7236;
  wire _net_7237;
  wire _net_7238;
  wire _net_7239;
  wire _net_7240;
  wire _net_7241;
  wire _net_7242;
  wire _net_7243;
  wire _net_7244;
  wire _net_7245;
  wire _net_7246;
  wire _net_7247;
  wire _net_7248;
  wire _net_7249;
  wire _net_7250;
  wire _net_7251;
  wire _net_7252;
  wire _net_7253;
  wire _net_7254;
  wire _net_7255;
  wire _net_7256;
  wire _net_7257;
  wire _net_7258;
  wire _net_7259;
  wire _net_7260;
  wire _net_7261;
  wire _net_7262;
  wire _net_7263;
  wire _net_7264;
  wire _net_7265;
  wire _net_7266;
  wire _net_7267;
  wire _net_7268;
  wire _net_7269;
  wire _net_7270;
  wire _net_7271;
  wire _net_7272;
  wire _net_7273;
  wire _net_7274;
  wire _net_7275;
  wire _net_7276;
  wire _net_7277;
  wire _net_7278;
  wire _net_7279;
  wire _net_7280;
  wire _net_7281;
  wire _net_7282;
  wire _net_7283;
  wire _net_7284;
  wire _net_7285;
  wire _net_7286;
  wire _net_7287;
  wire _net_7288;
  wire _net_7289;
  wire _net_7290;
  wire _net_7291;
  wire _net_7292;
  wire _net_7293;
  wire _net_7294;
  wire _net_7295;
  wire _net_7296;
  wire _net_7297;
  wire _net_7298;
  wire _net_7299;
  wire _net_7300;
  wire _net_7301;
  wire _net_7302;
  wire _net_7303;
  wire _net_7304;
  wire _net_7305;
  wire _net_7306;
  wire _net_7307;
  wire _net_7308;
  wire _net_7309;
  wire _net_7310;
  wire _net_7311;
  wire _net_7312;
  wire _net_7313;
  wire _net_7314;
  wire _net_7315;
  wire _net_7316;
  wire _net_7317;
  wire _net_7318;
  wire _net_7319;
  wire _net_7320;
  wire _net_7321;
  wire _net_7322;
  wire _net_7323;
  wire _net_7324;
  wire _net_7325;
  wire _net_7326;
  wire _net_7327;
  wire _net_7328;
  wire _net_7329;
  wire _net_7330;
  wire _net_7331;
  wire _net_7332;
  wire _net_7333;
  wire _net_7334;
  wire _net_7335;
  wire _net_7336;
  wire _net_7337;
  wire _net_7338;
  wire _net_7339;
  wire _net_7340;
  wire _net_7341;
  wire _net_7342;
  wire _net_7343;
  wire _net_7344;
  wire _net_7345;
  wire _net_7346;
  wire _net_7347;
  wire _net_7348;
  wire _net_7349;
  wire _net_7350;
  wire _net_7351;
  wire _net_7352;
  wire _net_7353;
  wire _net_7354;
  wire _net_7355;
  wire _net_7356;
  wire _net_7357;
  wire _net_7358;
  wire _net_7359;
  wire _net_7360;
  wire _net_7361;
  wire _net_7362;
  wire _net_7363;
  wire _net_7364;
  wire _net_7365;
  wire _net_7366;
  wire _net_7367;
  wire _net_7368;
  wire _net_7369;
  wire _net_7370;
  wire _net_7371;
  wire _net_7372;
  wire _net_7373;
  wire _net_7374;
  wire _net_7375;
  wire _net_7376;
  wire _net_7377;
  wire _net_7378;
  wire _net_7379;
  wire _net_7380;
  wire _net_7381;
  wire _net_7382;
  wire _net_7383;
  wire _net_7384;
  wire _net_7385;
  wire _net_7386;
  wire _net_7387;
  wire _net_7388;
  wire _net_7389;
  wire _net_7390;
  wire _net_7391;
  wire _net_7392;
  wire _net_7393;
  wire _net_7394;
  wire _net_7395;
  wire _net_7396;
  wire _net_7397;
  wire _net_7398;
  wire _net_7399;
  wire _net_7400;
  wire _net_7401;
  wire _net_7402;
  wire _net_7403;
  wire _net_7404;
  wire _net_7405;
  wire _net_7406;
  wire _net_7407;
  wire _net_7408;
  wire _net_7409;
  wire _net_7410;
  wire _net_7411;
  wire _net_7412;
  wire _net_7413;
  wire _net_7414;
  wire _net_7415;
  wire _net_7416;
  wire _net_7417;
  wire _net_7418;
  wire _net_7419;
  wire _net_7420;
  wire _net_7421;
  wire _net_7422;
  wire _net_7423;
  wire _net_7424;
  wire _net_7425;
  wire _net_7426;
  wire _net_7427;
  wire _net_7428;
  wire _net_7429;
  wire _net_7430;
  wire _net_7431;
  wire _net_7432;
  wire _net_7433;
  wire _net_7434;
  wire _net_7435;
  wire _net_7436;
  wire _net_7437;
  wire _net_7438;
  wire _net_7439;
  wire _net_7440;
  wire _net_7441;
  wire _net_7442;
  wire _net_7443;
  wire _net_7444;
  wire _net_7445;
  wire _net_7446;
  wire _net_7447;
  wire _net_7448;
  wire _net_7449;
  wire _net_7450;
  wire _net_7451;
  wire _net_7452;
  wire _net_7453;
  wire _net_7454;
  wire _net_7455;
  wire _net_7456;
  wire _net_7457;
  wire _net_7458;
  wire _net_7459;
  wire _net_7460;
  wire _net_7461;
  wire _net_7462;
  wire _net_7463;
  wire _net_7464;
  wire _net_7465;
  wire _net_7466;
  wire _net_7467;
  wire _net_7468;
  wire _net_7469;
  wire _net_7470;
  wire _net_7471;
  wire _net_7472;
  wire _net_7473;
  wire _net_7474;
  wire _net_7475;
  wire _net_7476;
  wire _net_7477;
  wire _net_7478;
  wire _net_7479;
  wire _net_7480;
  wire _net_7481;
  wire _net_7482;
  wire _net_7483;
  wire _net_7484;
  wire _net_7485;
  wire _net_7486;
  wire _net_7487;
  wire _net_7488;
  wire _net_7489;
  wire _net_7490;
  wire _net_7491;
  wire _net_7492;
  wire _net_7493;
  wire _net_7494;
  wire _net_7495;
  wire _net_7496;
  wire _net_7497;
  wire _net_7498;
  wire _net_7499;
  wire _net_7500;
  wire _net_7501;
  wire _net_7502;
  wire _net_7503;
  wire _net_7504;
  wire _net_7505;
  wire _net_7506;
  wire _net_7507;
  wire _net_7508;
  wire _net_7509;
  wire _net_7510;
  wire _net_7511;
  wire _net_7512;
  wire _net_7513;
  wire _net_7514;
  wire _net_7515;
  wire _net_7516;
  wire _net_7517;
  wire _net_7518;
  wire _net_7519;
  wire _net_7520;
  wire _net_7521;
  wire _net_7522;
  wire _net_7523;
  wire _net_7524;
  wire _net_7525;
  wire _net_7526;
  wire _net_7527;
  wire _net_7528;
  wire _net_7529;
  wire _net_7530;
  wire _net_7531;
  wire _net_7532;
  wire _net_7533;
  wire _net_7534;
  wire _net_7535;
  wire _net_7536;
  wire _net_7537;
  wire _net_7538;
  wire _net_7539;
  wire _net_7540;
  wire _net_7541;
  wire _net_7542;
  wire _net_7543;
  wire _net_7544;
  wire _net_7545;
  wire _net_7546;
  wire _net_7547;
  wire _net_7548;
  wire _net_7549;
  wire _net_7550;
  wire _net_7551;
  wire _net_7552;
  wire _net_7553;
  wire _net_7554;
  wire _net_7555;
  wire _net_7556;
  wire _net_7557;
  wire _net_7558;
  wire _net_7559;
  wire _net_7560;
  wire _net_7561;
  wire _net_7562;
  wire _net_7563;
  wire _net_7564;
  wire _net_7565;
  wire _net_7566;
  wire _net_7567;
  wire _net_7568;
  wire _net_7569;
  wire _net_7570;
  wire _net_7571;
  wire _net_7572;
  wire _net_7573;
  wire _net_7574;
  wire _net_7575;
  wire _net_7576;
  wire _net_7577;
  wire _net_7578;
  wire _net_7579;
  wire _net_7580;
  wire _net_7581;
  wire _net_7582;
  wire _net_7583;
  wire _net_7584;
  wire _net_7585;
  wire _net_7586;
  wire _net_7587;
  wire _net_7588;
  wire _net_7589;
  wire _net_7590;
  wire _net_7591;
  wire _net_7592;
  wire _net_7593;
  wire _net_7594;
  wire _net_7595;
  wire _net_7596;
  wire _net_7597;
  wire _net_7598;
  wire _net_7599;
  wire _net_7600;
  wire _net_7601;
  wire _net_7602;
  wire _net_7603;
  wire _net_7604;
  wire _net_7605;
  wire _net_7606;
  wire _net_7607;
  wire _net_7608;
  wire _net_7609;
  wire _net_7610;
  wire _net_7611;
  wire _net_7612;
  wire _net_7613;
  wire _net_7614;
  wire _net_7615;
  wire _net_7616;
  wire _net_7617;
  wire _net_7618;
  wire _net_7619;
  wire _net_7620;
  wire _net_7621;
  wire _net_7622;
  wire _net_7623;
  wire _net_7624;
  wire _net_7625;
  wire _net_7626;
  wire _net_7627;
  wire _net_7628;
  wire _net_7629;
  wire _net_7630;
  wire _net_7631;
  wire _net_7632;
  wire _net_7633;
  wire _net_7634;
  wire _net_7635;
  wire _net_7636;
  wire _net_7637;
  wire _net_7638;
  wire _net_7639;
  wire _net_7640;
  wire _net_7641;
  wire _net_7642;
  wire _net_7643;
  wire _net_7644;
  wire _net_7645;
  wire _net_7646;
  wire _net_7647;
  wire _net_7648;
  wire _net_7649;
  wire _net_7650;
  wire _net_7651;
  wire _net_7652;
  wire _net_7653;
  wire _net_7654;
  wire _net_7655;
  wire _net_7656;
  wire _net_7657;
  wire _net_7658;
  wire _net_7659;
  wire _net_7660;
  wire _net_7661;
  wire _net_7662;
  wire _net_7663;
  wire _net_7664;
  wire _net_7665;
  wire _net_7666;
  wire _net_7667;
  wire _net_7668;
  wire _net_7669;
  wire _net_7670;
  wire _net_7671;
  wire _net_7672;
  wire _net_7673;
  wire _net_7674;
  wire _net_7675;
  wire _net_7676;
  wire _net_7677;
  wire _net_7678;
  wire _net_7679;
  wire _net_7680;
  wire _net_7681;
  wire _net_7682;
  wire _net_7683;
  wire _net_7684;
  wire _net_7685;
  wire _net_7686;
  wire _net_7687;
  wire _net_7688;
  wire _net_7689;
  wire _net_7690;
  wire _net_7691;
  wire _net_7692;
  wire _net_7693;
  wire _net_7694;
  wire _net_7695;
  wire _net_7696;
  wire _net_7697;
  wire _net_7698;
  wire _net_7699;
  wire _net_7700;
  wire _net_7701;
  wire _net_7702;
  wire _net_7703;
  wire _net_7704;
  wire _net_7705;
  wire _net_7706;
  wire _net_7707;
  wire _net_7708;
  wire _net_7709;
  wire _net_7710;
  wire _net_7711;
  wire _net_7712;
  wire _net_7713;
  wire _net_7714;
  wire _net_7715;
  wire _net_7716;
  wire _net_7717;
  wire _net_7718;
  wire _net_7719;
  wire _net_7720;
  wire _net_7721;
  wire _net_7722;
  wire _net_7723;
  wire _net_7724;
  wire _net_7725;
  wire _net_7726;
  wire _net_7727;
  wire _net_7728;
  wire _net_7729;
  wire _net_7730;
  wire _net_7731;
  wire _net_7732;
  wire _net_7733;
  wire _net_7734;
  wire _net_7735;
  wire _net_7736;
  wire _net_7737;
  wire _net_7738;
  wire _net_7739;
  wire _net_7740;
  wire _net_7741;
  wire _net_7742;
  wire _net_7743;
  wire _net_7744;
  wire _net_7745;
  wire _net_7746;
  wire _net_7747;
  wire _net_7748;
  wire _net_7749;
  wire _net_7750;
  wire _net_7751;
  wire _net_7752;
  wire _net_7753;
  wire _net_7754;
  wire _net_7755;
  wire _net_7756;
  wire _net_7757;
  wire _net_7758;
  wire _net_7759;
  wire _net_7760;
  wire _net_7761;
  wire _net_7762;
  wire _net_7763;
  wire _net_7764;
  wire _net_7765;
  wire _net_7766;
  wire _net_7767;
  wire _net_7768;
  wire _net_7769;
  wire _net_7770;
  wire _net_7771;
  wire _net_7772;
  wire _net_7773;
  wire _net_7774;
  wire _net_7775;
  wire _net_7776;
  wire _net_7777;
  wire _net_7778;
  wire _net_7779;
  wire _net_7780;
  wire _net_7781;
  wire _net_7782;
  wire _net_7783;
  wire _net_7784;
  wire _net_7785;
  wire _net_7786;
  wire _net_7787;
  wire _net_7788;
  wire _net_7789;
  wire _net_7790;
  wire _net_7791;
  wire _net_7792;
  wire _net_7793;
  wire _net_7794;
  wire _net_7795;
  wire _net_7796;
  wire _net_7797;
  wire _net_7798;
  wire _net_7799;
  wire _net_7800;
  wire _net_7801;
  wire _net_7802;
  wire _net_7803;
  wire _net_7804;
  wire _net_7805;
  wire _net_7806;
  wire _net_7807;
  wire _net_7808;
  wire _net_7809;
  wire _net_7810;
  wire _net_7811;
  wire _net_7812;
  wire _net_7813;
  wire _net_7814;
  wire _net_7815;
  wire _net_7816;
  wire _net_7817;
  wire _net_7818;
  wire _net_7819;
  wire _net_7820;
  wire _net_7821;
  wire _net_7822;
  wire _net_7823;
  wire _net_7824;
  wire _net_7825;
  wire _net_7826;
  wire _net_7827;
  wire _net_7828;
  wire _net_7829;
  wire _net_7830;
  wire _net_7831;
  wire _net_7832;
  wire _net_7833;
  wire _net_7834;
  wire _net_7835;
  wire _net_7836;
  wire _net_7837;
  wire _net_7838;
  wire _net_7839;
  wire _net_7840;
  wire _net_7841;
  wire _net_7842;
  wire _net_7843;
  wire _net_7844;
  wire _net_7845;
  wire _net_7846;
  wire _net_7847;
  wire _net_7848;
  wire _net_7849;
  wire _net_7850;
  wire _net_7851;
  wire _net_7852;
  wire _net_7853;
  wire _net_7854;
  wire _net_7855;
  wire _net_7856;
  wire _net_7857;
  wire _net_7858;
  wire _net_7859;
  wire _net_7860;
  wire _net_7861;
  wire _net_7862;
  wire _net_7863;
  wire _net_7864;
  wire _net_7865;
  wire _net_7866;
  wire _net_7867;
  wire _net_7868;
  wire _net_7869;
  wire _net_7870;
  wire _net_7871;
  wire _net_7872;
  wire _net_7873;
  wire _net_7874;
  wire _net_7875;
  wire _net_7876;
  wire _net_7877;
  wire _net_7878;
  wire _net_7879;
  wire _net_7880;
  wire _net_7881;
  wire _net_7882;
  wire _net_7883;
  wire _net_7884;
  wire _net_7885;
  wire _net_7886;
  wire _net_7887;
  wire _net_7888;
  wire _net_7889;
  wire _net_7890;
  wire _net_7891;
  wire _net_7892;
  wire _net_7893;
  wire _net_7894;
  wire _net_7895;
  wire _net_7896;
  wire _net_7897;
  wire _net_7898;
  wire _net_7899;
  wire _net_7900;
  wire _net_7901;
  wire _net_7902;
  wire _net_7903;
  wire _net_7904;
  wire _net_7905;
  wire _net_7906;
  wire _net_7907;
  wire _net_7908;
  wire _net_7909;
  wire _net_7910;
  wire _net_7911;
  wire _net_7912;
  wire _net_7913;
  wire _net_7914;
  wire _net_7915;
  wire _net_7916;
  wire _net_7917;
  wire _net_7918;
  wire _net_7919;
  wire _net_7920;
  wire _net_7921;
  wire _net_7922;
  wire _net_7923;
  wire _net_7924;
  wire _net_7925;
  wire _net_7926;
  wire _net_7927;
  wire _net_7928;
  wire _net_7929;
  wire _net_7930;
  wire _net_7931;
  wire _net_7932;
  wire _net_7933;
  wire _net_7934;
  wire _net_7935;
  wire _net_7936;
  wire _net_7937;
  wire _net_7938;
  wire _net_7939;
  wire _net_7940;
  wire _net_7941;
  wire _net_7942;
  wire _net_7943;
  wire _net_7944;
  wire _net_7945;
  wire _net_7946;
  wire _net_7947;
  wire _net_7948;
  wire _net_7949;
  wire _net_7950;
  wire _net_7951;
  wire _net_7952;
  wire _net_7953;
  wire _net_7954;
  wire _net_7955;
  wire _net_7956;
  wire _net_7957;
  wire _net_7958;
  wire _net_7959;
  wire _net_7960;
  wire _net_7961;
  wire _net_7962;
  wire _net_7963;
  wire _net_7964;
  wire _net_7965;
  wire _net_7966;
  wire _net_7967;
  wire _net_7968;
  wire _net_7969;
  wire _net_7970;
  wire _net_7971;
  wire _net_7972;
  wire _net_7973;
  wire _net_7974;
  wire _net_7975;
  wire _net_7976;
  wire _net_7977;
  wire _net_7978;
  wire _net_7979;
  wire _net_7980;
  wire _net_7981;
  wire _net_7982;
  wire _net_7983;
  wire _net_7984;
  wire _net_7985;
add_map add_map_x (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_add_exe), .data_out(_add_map_x_data_out), .data_out_index(_add_map_x_data_out_index), .data_near(_add_map_x_data_near), .wall_t_out(_add_map_x_wall_t_out), .data_org(_add_map_x_data_org), .data_org_near(_add_map_x_data_org_near), .s_g(_add_map_x_s_g), .s_g_near(_add_map_x_s_g_near), .moto_org_near(_add_map_x_moto_org_near), .moto_org_near1(_add_map_x_moto_org_near1), .moto_org_near2(_add_map_x_moto_org_near2), .moto_org_near3(_add_map_x_moto_org_near3), .moto_org(_add_map_x_moto_org), .sg_up(_add_map_x_sg_up), .sg_down(_add_map_x_sg_down), .sg_left(_add_map_x_sg_left), .sg_right(_add_map_x_sg_right), .wall_t_in(_add_map_x_wall_t_in), .moto(_add_map_x_moto), .up(_add_map_x_up), .right(_add_map_x_right), .down(_add_map_x_down), .left(_add_map_x_left), .start(_add_map_x_start), .goal(_add_map_x_goal), .now(_add_map_x_now));
add_map add_map_x_209 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_209_add_exe), .data_out(_add_map_x_209_data_out), .data_out_index(_add_map_x_209_data_out_index), .data_near(_add_map_x_209_data_near), .wall_t_out(_add_map_x_209_wall_t_out), .data_org(_add_map_x_209_data_org), .data_org_near(_add_map_x_209_data_org_near), .s_g(_add_map_x_209_s_g), .s_g_near(_add_map_x_209_s_g_near), .moto_org_near(_add_map_x_209_moto_org_near), .moto_org_near1(_add_map_x_209_moto_org_near1), .moto_org_near2(_add_map_x_209_moto_org_near2), .moto_org_near3(_add_map_x_209_moto_org_near3), .moto_org(_add_map_x_209_moto_org), .sg_up(_add_map_x_209_sg_up), .sg_down(_add_map_x_209_sg_down), .sg_left(_add_map_x_209_sg_left), .sg_right(_add_map_x_209_sg_right), .wall_t_in(_add_map_x_209_wall_t_in), .moto(_add_map_x_209_moto), .up(_add_map_x_209_up), .right(_add_map_x_209_right), .down(_add_map_x_209_down), .left(_add_map_x_209_left), .start(_add_map_x_209_start), .goal(_add_map_x_209_goal), .now(_add_map_x_209_now));
add_map add_map_x_208 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_208_add_exe), .data_out(_add_map_x_208_data_out), .data_out_index(_add_map_x_208_data_out_index), .data_near(_add_map_x_208_data_near), .wall_t_out(_add_map_x_208_wall_t_out), .data_org(_add_map_x_208_data_org), .data_org_near(_add_map_x_208_data_org_near), .s_g(_add_map_x_208_s_g), .s_g_near(_add_map_x_208_s_g_near), .moto_org_near(_add_map_x_208_moto_org_near), .moto_org_near1(_add_map_x_208_moto_org_near1), .moto_org_near2(_add_map_x_208_moto_org_near2), .moto_org_near3(_add_map_x_208_moto_org_near3), .moto_org(_add_map_x_208_moto_org), .sg_up(_add_map_x_208_sg_up), .sg_down(_add_map_x_208_sg_down), .sg_left(_add_map_x_208_sg_left), .sg_right(_add_map_x_208_sg_right), .wall_t_in(_add_map_x_208_wall_t_in), .moto(_add_map_x_208_moto), .up(_add_map_x_208_up), .right(_add_map_x_208_right), .down(_add_map_x_208_down), .left(_add_map_x_208_left), .start(_add_map_x_208_start), .goal(_add_map_x_208_goal), .now(_add_map_x_208_now));
add_map add_map_x_207 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_207_add_exe), .data_out(_add_map_x_207_data_out), .data_out_index(_add_map_x_207_data_out_index), .data_near(_add_map_x_207_data_near), .wall_t_out(_add_map_x_207_wall_t_out), .data_org(_add_map_x_207_data_org), .data_org_near(_add_map_x_207_data_org_near), .s_g(_add_map_x_207_s_g), .s_g_near(_add_map_x_207_s_g_near), .moto_org_near(_add_map_x_207_moto_org_near), .moto_org_near1(_add_map_x_207_moto_org_near1), .moto_org_near2(_add_map_x_207_moto_org_near2), .moto_org_near3(_add_map_x_207_moto_org_near3), .moto_org(_add_map_x_207_moto_org), .sg_up(_add_map_x_207_sg_up), .sg_down(_add_map_x_207_sg_down), .sg_left(_add_map_x_207_sg_left), .sg_right(_add_map_x_207_sg_right), .wall_t_in(_add_map_x_207_wall_t_in), .moto(_add_map_x_207_moto), .up(_add_map_x_207_up), .right(_add_map_x_207_right), .down(_add_map_x_207_down), .left(_add_map_x_207_left), .start(_add_map_x_207_start), .goal(_add_map_x_207_goal), .now(_add_map_x_207_now));
add_map add_map_x_206 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_206_add_exe), .data_out(_add_map_x_206_data_out), .data_out_index(_add_map_x_206_data_out_index), .data_near(_add_map_x_206_data_near), .wall_t_out(_add_map_x_206_wall_t_out), .data_org(_add_map_x_206_data_org), .data_org_near(_add_map_x_206_data_org_near), .s_g(_add_map_x_206_s_g), .s_g_near(_add_map_x_206_s_g_near), .moto_org_near(_add_map_x_206_moto_org_near), .moto_org_near1(_add_map_x_206_moto_org_near1), .moto_org_near2(_add_map_x_206_moto_org_near2), .moto_org_near3(_add_map_x_206_moto_org_near3), .moto_org(_add_map_x_206_moto_org), .sg_up(_add_map_x_206_sg_up), .sg_down(_add_map_x_206_sg_down), .sg_left(_add_map_x_206_sg_left), .sg_right(_add_map_x_206_sg_right), .wall_t_in(_add_map_x_206_wall_t_in), .moto(_add_map_x_206_moto), .up(_add_map_x_206_up), .right(_add_map_x_206_right), .down(_add_map_x_206_down), .left(_add_map_x_206_left), .start(_add_map_x_206_start), .goal(_add_map_x_206_goal), .now(_add_map_x_206_now));
add_map add_map_x_205 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_205_add_exe), .data_out(_add_map_x_205_data_out), .data_out_index(_add_map_x_205_data_out_index), .data_near(_add_map_x_205_data_near), .wall_t_out(_add_map_x_205_wall_t_out), .data_org(_add_map_x_205_data_org), .data_org_near(_add_map_x_205_data_org_near), .s_g(_add_map_x_205_s_g), .s_g_near(_add_map_x_205_s_g_near), .moto_org_near(_add_map_x_205_moto_org_near), .moto_org_near1(_add_map_x_205_moto_org_near1), .moto_org_near2(_add_map_x_205_moto_org_near2), .moto_org_near3(_add_map_x_205_moto_org_near3), .moto_org(_add_map_x_205_moto_org), .sg_up(_add_map_x_205_sg_up), .sg_down(_add_map_x_205_sg_down), .sg_left(_add_map_x_205_sg_left), .sg_right(_add_map_x_205_sg_right), .wall_t_in(_add_map_x_205_wall_t_in), .moto(_add_map_x_205_moto), .up(_add_map_x_205_up), .right(_add_map_x_205_right), .down(_add_map_x_205_down), .left(_add_map_x_205_left), .start(_add_map_x_205_start), .goal(_add_map_x_205_goal), .now(_add_map_x_205_now));
add_map add_map_x_204 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_204_add_exe), .data_out(_add_map_x_204_data_out), .data_out_index(_add_map_x_204_data_out_index), .data_near(_add_map_x_204_data_near), .wall_t_out(_add_map_x_204_wall_t_out), .data_org(_add_map_x_204_data_org), .data_org_near(_add_map_x_204_data_org_near), .s_g(_add_map_x_204_s_g), .s_g_near(_add_map_x_204_s_g_near), .moto_org_near(_add_map_x_204_moto_org_near), .moto_org_near1(_add_map_x_204_moto_org_near1), .moto_org_near2(_add_map_x_204_moto_org_near2), .moto_org_near3(_add_map_x_204_moto_org_near3), .moto_org(_add_map_x_204_moto_org), .sg_up(_add_map_x_204_sg_up), .sg_down(_add_map_x_204_sg_down), .sg_left(_add_map_x_204_sg_left), .sg_right(_add_map_x_204_sg_right), .wall_t_in(_add_map_x_204_wall_t_in), .moto(_add_map_x_204_moto), .up(_add_map_x_204_up), .right(_add_map_x_204_right), .down(_add_map_x_204_down), .left(_add_map_x_204_left), .start(_add_map_x_204_start), .goal(_add_map_x_204_goal), .now(_add_map_x_204_now));
add_map add_map_x_203 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_203_add_exe), .data_out(_add_map_x_203_data_out), .data_out_index(_add_map_x_203_data_out_index), .data_near(_add_map_x_203_data_near), .wall_t_out(_add_map_x_203_wall_t_out), .data_org(_add_map_x_203_data_org), .data_org_near(_add_map_x_203_data_org_near), .s_g(_add_map_x_203_s_g), .s_g_near(_add_map_x_203_s_g_near), .moto_org_near(_add_map_x_203_moto_org_near), .moto_org_near1(_add_map_x_203_moto_org_near1), .moto_org_near2(_add_map_x_203_moto_org_near2), .moto_org_near3(_add_map_x_203_moto_org_near3), .moto_org(_add_map_x_203_moto_org), .sg_up(_add_map_x_203_sg_up), .sg_down(_add_map_x_203_sg_down), .sg_left(_add_map_x_203_sg_left), .sg_right(_add_map_x_203_sg_right), .wall_t_in(_add_map_x_203_wall_t_in), .moto(_add_map_x_203_moto), .up(_add_map_x_203_up), .right(_add_map_x_203_right), .down(_add_map_x_203_down), .left(_add_map_x_203_left), .start(_add_map_x_203_start), .goal(_add_map_x_203_goal), .now(_add_map_x_203_now));
add_map add_map_x_202 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_202_add_exe), .data_out(_add_map_x_202_data_out), .data_out_index(_add_map_x_202_data_out_index), .data_near(_add_map_x_202_data_near), .wall_t_out(_add_map_x_202_wall_t_out), .data_org(_add_map_x_202_data_org), .data_org_near(_add_map_x_202_data_org_near), .s_g(_add_map_x_202_s_g), .s_g_near(_add_map_x_202_s_g_near), .moto_org_near(_add_map_x_202_moto_org_near), .moto_org_near1(_add_map_x_202_moto_org_near1), .moto_org_near2(_add_map_x_202_moto_org_near2), .moto_org_near3(_add_map_x_202_moto_org_near3), .moto_org(_add_map_x_202_moto_org), .sg_up(_add_map_x_202_sg_up), .sg_down(_add_map_x_202_sg_down), .sg_left(_add_map_x_202_sg_left), .sg_right(_add_map_x_202_sg_right), .wall_t_in(_add_map_x_202_wall_t_in), .moto(_add_map_x_202_moto), .up(_add_map_x_202_up), .right(_add_map_x_202_right), .down(_add_map_x_202_down), .left(_add_map_x_202_left), .start(_add_map_x_202_start), .goal(_add_map_x_202_goal), .now(_add_map_x_202_now));
add_map add_map_x_201 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_201_add_exe), .data_out(_add_map_x_201_data_out), .data_out_index(_add_map_x_201_data_out_index), .data_near(_add_map_x_201_data_near), .wall_t_out(_add_map_x_201_wall_t_out), .data_org(_add_map_x_201_data_org), .data_org_near(_add_map_x_201_data_org_near), .s_g(_add_map_x_201_s_g), .s_g_near(_add_map_x_201_s_g_near), .moto_org_near(_add_map_x_201_moto_org_near), .moto_org_near1(_add_map_x_201_moto_org_near1), .moto_org_near2(_add_map_x_201_moto_org_near2), .moto_org_near3(_add_map_x_201_moto_org_near3), .moto_org(_add_map_x_201_moto_org), .sg_up(_add_map_x_201_sg_up), .sg_down(_add_map_x_201_sg_down), .sg_left(_add_map_x_201_sg_left), .sg_right(_add_map_x_201_sg_right), .wall_t_in(_add_map_x_201_wall_t_in), .moto(_add_map_x_201_moto), .up(_add_map_x_201_up), .right(_add_map_x_201_right), .down(_add_map_x_201_down), .left(_add_map_x_201_left), .start(_add_map_x_201_start), .goal(_add_map_x_201_goal), .now(_add_map_x_201_now));
add_map add_map_x_200 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_200_add_exe), .data_out(_add_map_x_200_data_out), .data_out_index(_add_map_x_200_data_out_index), .data_near(_add_map_x_200_data_near), .wall_t_out(_add_map_x_200_wall_t_out), .data_org(_add_map_x_200_data_org), .data_org_near(_add_map_x_200_data_org_near), .s_g(_add_map_x_200_s_g), .s_g_near(_add_map_x_200_s_g_near), .moto_org_near(_add_map_x_200_moto_org_near), .moto_org_near1(_add_map_x_200_moto_org_near1), .moto_org_near2(_add_map_x_200_moto_org_near2), .moto_org_near3(_add_map_x_200_moto_org_near3), .moto_org(_add_map_x_200_moto_org), .sg_up(_add_map_x_200_sg_up), .sg_down(_add_map_x_200_sg_down), .sg_left(_add_map_x_200_sg_left), .sg_right(_add_map_x_200_sg_right), .wall_t_in(_add_map_x_200_wall_t_in), .moto(_add_map_x_200_moto), .up(_add_map_x_200_up), .right(_add_map_x_200_right), .down(_add_map_x_200_down), .left(_add_map_x_200_left), .start(_add_map_x_200_start), .goal(_add_map_x_200_goal), .now(_add_map_x_200_now));
add_map add_map_x_199 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_199_add_exe), .data_out(_add_map_x_199_data_out), .data_out_index(_add_map_x_199_data_out_index), .data_near(_add_map_x_199_data_near), .wall_t_out(_add_map_x_199_wall_t_out), .data_org(_add_map_x_199_data_org), .data_org_near(_add_map_x_199_data_org_near), .s_g(_add_map_x_199_s_g), .s_g_near(_add_map_x_199_s_g_near), .moto_org_near(_add_map_x_199_moto_org_near), .moto_org_near1(_add_map_x_199_moto_org_near1), .moto_org_near2(_add_map_x_199_moto_org_near2), .moto_org_near3(_add_map_x_199_moto_org_near3), .moto_org(_add_map_x_199_moto_org), .sg_up(_add_map_x_199_sg_up), .sg_down(_add_map_x_199_sg_down), .sg_left(_add_map_x_199_sg_left), .sg_right(_add_map_x_199_sg_right), .wall_t_in(_add_map_x_199_wall_t_in), .moto(_add_map_x_199_moto), .up(_add_map_x_199_up), .right(_add_map_x_199_right), .down(_add_map_x_199_down), .left(_add_map_x_199_left), .start(_add_map_x_199_start), .goal(_add_map_x_199_goal), .now(_add_map_x_199_now));
add_map add_map_x_198 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_198_add_exe), .data_out(_add_map_x_198_data_out), .data_out_index(_add_map_x_198_data_out_index), .data_near(_add_map_x_198_data_near), .wall_t_out(_add_map_x_198_wall_t_out), .data_org(_add_map_x_198_data_org), .data_org_near(_add_map_x_198_data_org_near), .s_g(_add_map_x_198_s_g), .s_g_near(_add_map_x_198_s_g_near), .moto_org_near(_add_map_x_198_moto_org_near), .moto_org_near1(_add_map_x_198_moto_org_near1), .moto_org_near2(_add_map_x_198_moto_org_near2), .moto_org_near3(_add_map_x_198_moto_org_near3), .moto_org(_add_map_x_198_moto_org), .sg_up(_add_map_x_198_sg_up), .sg_down(_add_map_x_198_sg_down), .sg_left(_add_map_x_198_sg_left), .sg_right(_add_map_x_198_sg_right), .wall_t_in(_add_map_x_198_wall_t_in), .moto(_add_map_x_198_moto), .up(_add_map_x_198_up), .right(_add_map_x_198_right), .down(_add_map_x_198_down), .left(_add_map_x_198_left), .start(_add_map_x_198_start), .goal(_add_map_x_198_goal), .now(_add_map_x_198_now));
add_map add_map_x_197 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_197_add_exe), .data_out(_add_map_x_197_data_out), .data_out_index(_add_map_x_197_data_out_index), .data_near(_add_map_x_197_data_near), .wall_t_out(_add_map_x_197_wall_t_out), .data_org(_add_map_x_197_data_org), .data_org_near(_add_map_x_197_data_org_near), .s_g(_add_map_x_197_s_g), .s_g_near(_add_map_x_197_s_g_near), .moto_org_near(_add_map_x_197_moto_org_near), .moto_org_near1(_add_map_x_197_moto_org_near1), .moto_org_near2(_add_map_x_197_moto_org_near2), .moto_org_near3(_add_map_x_197_moto_org_near3), .moto_org(_add_map_x_197_moto_org), .sg_up(_add_map_x_197_sg_up), .sg_down(_add_map_x_197_sg_down), .sg_left(_add_map_x_197_sg_left), .sg_right(_add_map_x_197_sg_right), .wall_t_in(_add_map_x_197_wall_t_in), .moto(_add_map_x_197_moto), .up(_add_map_x_197_up), .right(_add_map_x_197_right), .down(_add_map_x_197_down), .left(_add_map_x_197_left), .start(_add_map_x_197_start), .goal(_add_map_x_197_goal), .now(_add_map_x_197_now));
add_map add_map_x_196 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_196_add_exe), .data_out(_add_map_x_196_data_out), .data_out_index(_add_map_x_196_data_out_index), .data_near(_add_map_x_196_data_near), .wall_t_out(_add_map_x_196_wall_t_out), .data_org(_add_map_x_196_data_org), .data_org_near(_add_map_x_196_data_org_near), .s_g(_add_map_x_196_s_g), .s_g_near(_add_map_x_196_s_g_near), .moto_org_near(_add_map_x_196_moto_org_near), .moto_org_near1(_add_map_x_196_moto_org_near1), .moto_org_near2(_add_map_x_196_moto_org_near2), .moto_org_near3(_add_map_x_196_moto_org_near3), .moto_org(_add_map_x_196_moto_org), .sg_up(_add_map_x_196_sg_up), .sg_down(_add_map_x_196_sg_down), .sg_left(_add_map_x_196_sg_left), .sg_right(_add_map_x_196_sg_right), .wall_t_in(_add_map_x_196_wall_t_in), .moto(_add_map_x_196_moto), .up(_add_map_x_196_up), .right(_add_map_x_196_right), .down(_add_map_x_196_down), .left(_add_map_x_196_left), .start(_add_map_x_196_start), .goal(_add_map_x_196_goal), .now(_add_map_x_196_now));
add_map add_map_x_195 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_195_add_exe), .data_out(_add_map_x_195_data_out), .data_out_index(_add_map_x_195_data_out_index), .data_near(_add_map_x_195_data_near), .wall_t_out(_add_map_x_195_wall_t_out), .data_org(_add_map_x_195_data_org), .data_org_near(_add_map_x_195_data_org_near), .s_g(_add_map_x_195_s_g), .s_g_near(_add_map_x_195_s_g_near), .moto_org_near(_add_map_x_195_moto_org_near), .moto_org_near1(_add_map_x_195_moto_org_near1), .moto_org_near2(_add_map_x_195_moto_org_near2), .moto_org_near3(_add_map_x_195_moto_org_near3), .moto_org(_add_map_x_195_moto_org), .sg_up(_add_map_x_195_sg_up), .sg_down(_add_map_x_195_sg_down), .sg_left(_add_map_x_195_sg_left), .sg_right(_add_map_x_195_sg_right), .wall_t_in(_add_map_x_195_wall_t_in), .moto(_add_map_x_195_moto), .up(_add_map_x_195_up), .right(_add_map_x_195_right), .down(_add_map_x_195_down), .left(_add_map_x_195_left), .start(_add_map_x_195_start), .goal(_add_map_x_195_goal), .now(_add_map_x_195_now));
add_map add_map_x_194 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_194_add_exe), .data_out(_add_map_x_194_data_out), .data_out_index(_add_map_x_194_data_out_index), .data_near(_add_map_x_194_data_near), .wall_t_out(_add_map_x_194_wall_t_out), .data_org(_add_map_x_194_data_org), .data_org_near(_add_map_x_194_data_org_near), .s_g(_add_map_x_194_s_g), .s_g_near(_add_map_x_194_s_g_near), .moto_org_near(_add_map_x_194_moto_org_near), .moto_org_near1(_add_map_x_194_moto_org_near1), .moto_org_near2(_add_map_x_194_moto_org_near2), .moto_org_near3(_add_map_x_194_moto_org_near3), .moto_org(_add_map_x_194_moto_org), .sg_up(_add_map_x_194_sg_up), .sg_down(_add_map_x_194_sg_down), .sg_left(_add_map_x_194_sg_left), .sg_right(_add_map_x_194_sg_right), .wall_t_in(_add_map_x_194_wall_t_in), .moto(_add_map_x_194_moto), .up(_add_map_x_194_up), .right(_add_map_x_194_right), .down(_add_map_x_194_down), .left(_add_map_x_194_left), .start(_add_map_x_194_start), .goal(_add_map_x_194_goal), .now(_add_map_x_194_now));
add_map add_map_x_193 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_193_add_exe), .data_out(_add_map_x_193_data_out), .data_out_index(_add_map_x_193_data_out_index), .data_near(_add_map_x_193_data_near), .wall_t_out(_add_map_x_193_wall_t_out), .data_org(_add_map_x_193_data_org), .data_org_near(_add_map_x_193_data_org_near), .s_g(_add_map_x_193_s_g), .s_g_near(_add_map_x_193_s_g_near), .moto_org_near(_add_map_x_193_moto_org_near), .moto_org_near1(_add_map_x_193_moto_org_near1), .moto_org_near2(_add_map_x_193_moto_org_near2), .moto_org_near3(_add_map_x_193_moto_org_near3), .moto_org(_add_map_x_193_moto_org), .sg_up(_add_map_x_193_sg_up), .sg_down(_add_map_x_193_sg_down), .sg_left(_add_map_x_193_sg_left), .sg_right(_add_map_x_193_sg_right), .wall_t_in(_add_map_x_193_wall_t_in), .moto(_add_map_x_193_moto), .up(_add_map_x_193_up), .right(_add_map_x_193_right), .down(_add_map_x_193_down), .left(_add_map_x_193_left), .start(_add_map_x_193_start), .goal(_add_map_x_193_goal), .now(_add_map_x_193_now));
add_map add_map_x_192 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_192_add_exe), .data_out(_add_map_x_192_data_out), .data_out_index(_add_map_x_192_data_out_index), .data_near(_add_map_x_192_data_near), .wall_t_out(_add_map_x_192_wall_t_out), .data_org(_add_map_x_192_data_org), .data_org_near(_add_map_x_192_data_org_near), .s_g(_add_map_x_192_s_g), .s_g_near(_add_map_x_192_s_g_near), .moto_org_near(_add_map_x_192_moto_org_near), .moto_org_near1(_add_map_x_192_moto_org_near1), .moto_org_near2(_add_map_x_192_moto_org_near2), .moto_org_near3(_add_map_x_192_moto_org_near3), .moto_org(_add_map_x_192_moto_org), .sg_up(_add_map_x_192_sg_up), .sg_down(_add_map_x_192_sg_down), .sg_left(_add_map_x_192_sg_left), .sg_right(_add_map_x_192_sg_right), .wall_t_in(_add_map_x_192_wall_t_in), .moto(_add_map_x_192_moto), .up(_add_map_x_192_up), .right(_add_map_x_192_right), .down(_add_map_x_192_down), .left(_add_map_x_192_left), .start(_add_map_x_192_start), .goal(_add_map_x_192_goal), .now(_add_map_x_192_now));
add_map add_map_x_191 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_191_add_exe), .data_out(_add_map_x_191_data_out), .data_out_index(_add_map_x_191_data_out_index), .data_near(_add_map_x_191_data_near), .wall_t_out(_add_map_x_191_wall_t_out), .data_org(_add_map_x_191_data_org), .data_org_near(_add_map_x_191_data_org_near), .s_g(_add_map_x_191_s_g), .s_g_near(_add_map_x_191_s_g_near), .moto_org_near(_add_map_x_191_moto_org_near), .moto_org_near1(_add_map_x_191_moto_org_near1), .moto_org_near2(_add_map_x_191_moto_org_near2), .moto_org_near3(_add_map_x_191_moto_org_near3), .moto_org(_add_map_x_191_moto_org), .sg_up(_add_map_x_191_sg_up), .sg_down(_add_map_x_191_sg_down), .sg_left(_add_map_x_191_sg_left), .sg_right(_add_map_x_191_sg_right), .wall_t_in(_add_map_x_191_wall_t_in), .moto(_add_map_x_191_moto), .up(_add_map_x_191_up), .right(_add_map_x_191_right), .down(_add_map_x_191_down), .left(_add_map_x_191_left), .start(_add_map_x_191_start), .goal(_add_map_x_191_goal), .now(_add_map_x_191_now));
add_map add_map_x_190 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_190_add_exe), .data_out(_add_map_x_190_data_out), .data_out_index(_add_map_x_190_data_out_index), .data_near(_add_map_x_190_data_near), .wall_t_out(_add_map_x_190_wall_t_out), .data_org(_add_map_x_190_data_org), .data_org_near(_add_map_x_190_data_org_near), .s_g(_add_map_x_190_s_g), .s_g_near(_add_map_x_190_s_g_near), .moto_org_near(_add_map_x_190_moto_org_near), .moto_org_near1(_add_map_x_190_moto_org_near1), .moto_org_near2(_add_map_x_190_moto_org_near2), .moto_org_near3(_add_map_x_190_moto_org_near3), .moto_org(_add_map_x_190_moto_org), .sg_up(_add_map_x_190_sg_up), .sg_down(_add_map_x_190_sg_down), .sg_left(_add_map_x_190_sg_left), .sg_right(_add_map_x_190_sg_right), .wall_t_in(_add_map_x_190_wall_t_in), .moto(_add_map_x_190_moto), .up(_add_map_x_190_up), .right(_add_map_x_190_right), .down(_add_map_x_190_down), .left(_add_map_x_190_left), .start(_add_map_x_190_start), .goal(_add_map_x_190_goal), .now(_add_map_x_190_now));
add_map add_map_x_189 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_189_add_exe), .data_out(_add_map_x_189_data_out), .data_out_index(_add_map_x_189_data_out_index), .data_near(_add_map_x_189_data_near), .wall_t_out(_add_map_x_189_wall_t_out), .data_org(_add_map_x_189_data_org), .data_org_near(_add_map_x_189_data_org_near), .s_g(_add_map_x_189_s_g), .s_g_near(_add_map_x_189_s_g_near), .moto_org_near(_add_map_x_189_moto_org_near), .moto_org_near1(_add_map_x_189_moto_org_near1), .moto_org_near2(_add_map_x_189_moto_org_near2), .moto_org_near3(_add_map_x_189_moto_org_near3), .moto_org(_add_map_x_189_moto_org), .sg_up(_add_map_x_189_sg_up), .sg_down(_add_map_x_189_sg_down), .sg_left(_add_map_x_189_sg_left), .sg_right(_add_map_x_189_sg_right), .wall_t_in(_add_map_x_189_wall_t_in), .moto(_add_map_x_189_moto), .up(_add_map_x_189_up), .right(_add_map_x_189_right), .down(_add_map_x_189_down), .left(_add_map_x_189_left), .start(_add_map_x_189_start), .goal(_add_map_x_189_goal), .now(_add_map_x_189_now));
add_map add_map_x_188 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_188_add_exe), .data_out(_add_map_x_188_data_out), .data_out_index(_add_map_x_188_data_out_index), .data_near(_add_map_x_188_data_near), .wall_t_out(_add_map_x_188_wall_t_out), .data_org(_add_map_x_188_data_org), .data_org_near(_add_map_x_188_data_org_near), .s_g(_add_map_x_188_s_g), .s_g_near(_add_map_x_188_s_g_near), .moto_org_near(_add_map_x_188_moto_org_near), .moto_org_near1(_add_map_x_188_moto_org_near1), .moto_org_near2(_add_map_x_188_moto_org_near2), .moto_org_near3(_add_map_x_188_moto_org_near3), .moto_org(_add_map_x_188_moto_org), .sg_up(_add_map_x_188_sg_up), .sg_down(_add_map_x_188_sg_down), .sg_left(_add_map_x_188_sg_left), .sg_right(_add_map_x_188_sg_right), .wall_t_in(_add_map_x_188_wall_t_in), .moto(_add_map_x_188_moto), .up(_add_map_x_188_up), .right(_add_map_x_188_right), .down(_add_map_x_188_down), .left(_add_map_x_188_left), .start(_add_map_x_188_start), .goal(_add_map_x_188_goal), .now(_add_map_x_188_now));
add_map add_map_x_187 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_187_add_exe), .data_out(_add_map_x_187_data_out), .data_out_index(_add_map_x_187_data_out_index), .data_near(_add_map_x_187_data_near), .wall_t_out(_add_map_x_187_wall_t_out), .data_org(_add_map_x_187_data_org), .data_org_near(_add_map_x_187_data_org_near), .s_g(_add_map_x_187_s_g), .s_g_near(_add_map_x_187_s_g_near), .moto_org_near(_add_map_x_187_moto_org_near), .moto_org_near1(_add_map_x_187_moto_org_near1), .moto_org_near2(_add_map_x_187_moto_org_near2), .moto_org_near3(_add_map_x_187_moto_org_near3), .moto_org(_add_map_x_187_moto_org), .sg_up(_add_map_x_187_sg_up), .sg_down(_add_map_x_187_sg_down), .sg_left(_add_map_x_187_sg_left), .sg_right(_add_map_x_187_sg_right), .wall_t_in(_add_map_x_187_wall_t_in), .moto(_add_map_x_187_moto), .up(_add_map_x_187_up), .right(_add_map_x_187_right), .down(_add_map_x_187_down), .left(_add_map_x_187_left), .start(_add_map_x_187_start), .goal(_add_map_x_187_goal), .now(_add_map_x_187_now));
add_map add_map_x_186 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_186_add_exe), .data_out(_add_map_x_186_data_out), .data_out_index(_add_map_x_186_data_out_index), .data_near(_add_map_x_186_data_near), .wall_t_out(_add_map_x_186_wall_t_out), .data_org(_add_map_x_186_data_org), .data_org_near(_add_map_x_186_data_org_near), .s_g(_add_map_x_186_s_g), .s_g_near(_add_map_x_186_s_g_near), .moto_org_near(_add_map_x_186_moto_org_near), .moto_org_near1(_add_map_x_186_moto_org_near1), .moto_org_near2(_add_map_x_186_moto_org_near2), .moto_org_near3(_add_map_x_186_moto_org_near3), .moto_org(_add_map_x_186_moto_org), .sg_up(_add_map_x_186_sg_up), .sg_down(_add_map_x_186_sg_down), .sg_left(_add_map_x_186_sg_left), .sg_right(_add_map_x_186_sg_right), .wall_t_in(_add_map_x_186_wall_t_in), .moto(_add_map_x_186_moto), .up(_add_map_x_186_up), .right(_add_map_x_186_right), .down(_add_map_x_186_down), .left(_add_map_x_186_left), .start(_add_map_x_186_start), .goal(_add_map_x_186_goal), .now(_add_map_x_186_now));
add_map add_map_x_185 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_185_add_exe), .data_out(_add_map_x_185_data_out), .data_out_index(_add_map_x_185_data_out_index), .data_near(_add_map_x_185_data_near), .wall_t_out(_add_map_x_185_wall_t_out), .data_org(_add_map_x_185_data_org), .data_org_near(_add_map_x_185_data_org_near), .s_g(_add_map_x_185_s_g), .s_g_near(_add_map_x_185_s_g_near), .moto_org_near(_add_map_x_185_moto_org_near), .moto_org_near1(_add_map_x_185_moto_org_near1), .moto_org_near2(_add_map_x_185_moto_org_near2), .moto_org_near3(_add_map_x_185_moto_org_near3), .moto_org(_add_map_x_185_moto_org), .sg_up(_add_map_x_185_sg_up), .sg_down(_add_map_x_185_sg_down), .sg_left(_add_map_x_185_sg_left), .sg_right(_add_map_x_185_sg_right), .wall_t_in(_add_map_x_185_wall_t_in), .moto(_add_map_x_185_moto), .up(_add_map_x_185_up), .right(_add_map_x_185_right), .down(_add_map_x_185_down), .left(_add_map_x_185_left), .start(_add_map_x_185_start), .goal(_add_map_x_185_goal), .now(_add_map_x_185_now));
add_map add_map_x_184 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_184_add_exe), .data_out(_add_map_x_184_data_out), .data_out_index(_add_map_x_184_data_out_index), .data_near(_add_map_x_184_data_near), .wall_t_out(_add_map_x_184_wall_t_out), .data_org(_add_map_x_184_data_org), .data_org_near(_add_map_x_184_data_org_near), .s_g(_add_map_x_184_s_g), .s_g_near(_add_map_x_184_s_g_near), .moto_org_near(_add_map_x_184_moto_org_near), .moto_org_near1(_add_map_x_184_moto_org_near1), .moto_org_near2(_add_map_x_184_moto_org_near2), .moto_org_near3(_add_map_x_184_moto_org_near3), .moto_org(_add_map_x_184_moto_org), .sg_up(_add_map_x_184_sg_up), .sg_down(_add_map_x_184_sg_down), .sg_left(_add_map_x_184_sg_left), .sg_right(_add_map_x_184_sg_right), .wall_t_in(_add_map_x_184_wall_t_in), .moto(_add_map_x_184_moto), .up(_add_map_x_184_up), .right(_add_map_x_184_right), .down(_add_map_x_184_down), .left(_add_map_x_184_left), .start(_add_map_x_184_start), .goal(_add_map_x_184_goal), .now(_add_map_x_184_now));
add_map add_map_x_183 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_183_add_exe), .data_out(_add_map_x_183_data_out), .data_out_index(_add_map_x_183_data_out_index), .data_near(_add_map_x_183_data_near), .wall_t_out(_add_map_x_183_wall_t_out), .data_org(_add_map_x_183_data_org), .data_org_near(_add_map_x_183_data_org_near), .s_g(_add_map_x_183_s_g), .s_g_near(_add_map_x_183_s_g_near), .moto_org_near(_add_map_x_183_moto_org_near), .moto_org_near1(_add_map_x_183_moto_org_near1), .moto_org_near2(_add_map_x_183_moto_org_near2), .moto_org_near3(_add_map_x_183_moto_org_near3), .moto_org(_add_map_x_183_moto_org), .sg_up(_add_map_x_183_sg_up), .sg_down(_add_map_x_183_sg_down), .sg_left(_add_map_x_183_sg_left), .sg_right(_add_map_x_183_sg_right), .wall_t_in(_add_map_x_183_wall_t_in), .moto(_add_map_x_183_moto), .up(_add_map_x_183_up), .right(_add_map_x_183_right), .down(_add_map_x_183_down), .left(_add_map_x_183_left), .start(_add_map_x_183_start), .goal(_add_map_x_183_goal), .now(_add_map_x_183_now));
add_map add_map_x_182 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_182_add_exe), .data_out(_add_map_x_182_data_out), .data_out_index(_add_map_x_182_data_out_index), .data_near(_add_map_x_182_data_near), .wall_t_out(_add_map_x_182_wall_t_out), .data_org(_add_map_x_182_data_org), .data_org_near(_add_map_x_182_data_org_near), .s_g(_add_map_x_182_s_g), .s_g_near(_add_map_x_182_s_g_near), .moto_org_near(_add_map_x_182_moto_org_near), .moto_org_near1(_add_map_x_182_moto_org_near1), .moto_org_near2(_add_map_x_182_moto_org_near2), .moto_org_near3(_add_map_x_182_moto_org_near3), .moto_org(_add_map_x_182_moto_org), .sg_up(_add_map_x_182_sg_up), .sg_down(_add_map_x_182_sg_down), .sg_left(_add_map_x_182_sg_left), .sg_right(_add_map_x_182_sg_right), .wall_t_in(_add_map_x_182_wall_t_in), .moto(_add_map_x_182_moto), .up(_add_map_x_182_up), .right(_add_map_x_182_right), .down(_add_map_x_182_down), .left(_add_map_x_182_left), .start(_add_map_x_182_start), .goal(_add_map_x_182_goal), .now(_add_map_x_182_now));
add_map add_map_x_181 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_181_add_exe), .data_out(_add_map_x_181_data_out), .data_out_index(_add_map_x_181_data_out_index), .data_near(_add_map_x_181_data_near), .wall_t_out(_add_map_x_181_wall_t_out), .data_org(_add_map_x_181_data_org), .data_org_near(_add_map_x_181_data_org_near), .s_g(_add_map_x_181_s_g), .s_g_near(_add_map_x_181_s_g_near), .moto_org_near(_add_map_x_181_moto_org_near), .moto_org_near1(_add_map_x_181_moto_org_near1), .moto_org_near2(_add_map_x_181_moto_org_near2), .moto_org_near3(_add_map_x_181_moto_org_near3), .moto_org(_add_map_x_181_moto_org), .sg_up(_add_map_x_181_sg_up), .sg_down(_add_map_x_181_sg_down), .sg_left(_add_map_x_181_sg_left), .sg_right(_add_map_x_181_sg_right), .wall_t_in(_add_map_x_181_wall_t_in), .moto(_add_map_x_181_moto), .up(_add_map_x_181_up), .right(_add_map_x_181_right), .down(_add_map_x_181_down), .left(_add_map_x_181_left), .start(_add_map_x_181_start), .goal(_add_map_x_181_goal), .now(_add_map_x_181_now));
add_map add_map_x_180 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_180_add_exe), .data_out(_add_map_x_180_data_out), .data_out_index(_add_map_x_180_data_out_index), .data_near(_add_map_x_180_data_near), .wall_t_out(_add_map_x_180_wall_t_out), .data_org(_add_map_x_180_data_org), .data_org_near(_add_map_x_180_data_org_near), .s_g(_add_map_x_180_s_g), .s_g_near(_add_map_x_180_s_g_near), .moto_org_near(_add_map_x_180_moto_org_near), .moto_org_near1(_add_map_x_180_moto_org_near1), .moto_org_near2(_add_map_x_180_moto_org_near2), .moto_org_near3(_add_map_x_180_moto_org_near3), .moto_org(_add_map_x_180_moto_org), .sg_up(_add_map_x_180_sg_up), .sg_down(_add_map_x_180_sg_down), .sg_left(_add_map_x_180_sg_left), .sg_right(_add_map_x_180_sg_right), .wall_t_in(_add_map_x_180_wall_t_in), .moto(_add_map_x_180_moto), .up(_add_map_x_180_up), .right(_add_map_x_180_right), .down(_add_map_x_180_down), .left(_add_map_x_180_left), .start(_add_map_x_180_start), .goal(_add_map_x_180_goal), .now(_add_map_x_180_now));
add_map add_map_x_179 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_179_add_exe), .data_out(_add_map_x_179_data_out), .data_out_index(_add_map_x_179_data_out_index), .data_near(_add_map_x_179_data_near), .wall_t_out(_add_map_x_179_wall_t_out), .data_org(_add_map_x_179_data_org), .data_org_near(_add_map_x_179_data_org_near), .s_g(_add_map_x_179_s_g), .s_g_near(_add_map_x_179_s_g_near), .moto_org_near(_add_map_x_179_moto_org_near), .moto_org_near1(_add_map_x_179_moto_org_near1), .moto_org_near2(_add_map_x_179_moto_org_near2), .moto_org_near3(_add_map_x_179_moto_org_near3), .moto_org(_add_map_x_179_moto_org), .sg_up(_add_map_x_179_sg_up), .sg_down(_add_map_x_179_sg_down), .sg_left(_add_map_x_179_sg_left), .sg_right(_add_map_x_179_sg_right), .wall_t_in(_add_map_x_179_wall_t_in), .moto(_add_map_x_179_moto), .up(_add_map_x_179_up), .right(_add_map_x_179_right), .down(_add_map_x_179_down), .left(_add_map_x_179_left), .start(_add_map_x_179_start), .goal(_add_map_x_179_goal), .now(_add_map_x_179_now));
add_map add_map_x_178 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_178_add_exe), .data_out(_add_map_x_178_data_out), .data_out_index(_add_map_x_178_data_out_index), .data_near(_add_map_x_178_data_near), .wall_t_out(_add_map_x_178_wall_t_out), .data_org(_add_map_x_178_data_org), .data_org_near(_add_map_x_178_data_org_near), .s_g(_add_map_x_178_s_g), .s_g_near(_add_map_x_178_s_g_near), .moto_org_near(_add_map_x_178_moto_org_near), .moto_org_near1(_add_map_x_178_moto_org_near1), .moto_org_near2(_add_map_x_178_moto_org_near2), .moto_org_near3(_add_map_x_178_moto_org_near3), .moto_org(_add_map_x_178_moto_org), .sg_up(_add_map_x_178_sg_up), .sg_down(_add_map_x_178_sg_down), .sg_left(_add_map_x_178_sg_left), .sg_right(_add_map_x_178_sg_right), .wall_t_in(_add_map_x_178_wall_t_in), .moto(_add_map_x_178_moto), .up(_add_map_x_178_up), .right(_add_map_x_178_right), .down(_add_map_x_178_down), .left(_add_map_x_178_left), .start(_add_map_x_178_start), .goal(_add_map_x_178_goal), .now(_add_map_x_178_now));
add_map add_map_x_177 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_177_add_exe), .data_out(_add_map_x_177_data_out), .data_out_index(_add_map_x_177_data_out_index), .data_near(_add_map_x_177_data_near), .wall_t_out(_add_map_x_177_wall_t_out), .data_org(_add_map_x_177_data_org), .data_org_near(_add_map_x_177_data_org_near), .s_g(_add_map_x_177_s_g), .s_g_near(_add_map_x_177_s_g_near), .moto_org_near(_add_map_x_177_moto_org_near), .moto_org_near1(_add_map_x_177_moto_org_near1), .moto_org_near2(_add_map_x_177_moto_org_near2), .moto_org_near3(_add_map_x_177_moto_org_near3), .moto_org(_add_map_x_177_moto_org), .sg_up(_add_map_x_177_sg_up), .sg_down(_add_map_x_177_sg_down), .sg_left(_add_map_x_177_sg_left), .sg_right(_add_map_x_177_sg_right), .wall_t_in(_add_map_x_177_wall_t_in), .moto(_add_map_x_177_moto), .up(_add_map_x_177_up), .right(_add_map_x_177_right), .down(_add_map_x_177_down), .left(_add_map_x_177_left), .start(_add_map_x_177_start), .goal(_add_map_x_177_goal), .now(_add_map_x_177_now));
add_map add_map_x_176 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_176_add_exe), .data_out(_add_map_x_176_data_out), .data_out_index(_add_map_x_176_data_out_index), .data_near(_add_map_x_176_data_near), .wall_t_out(_add_map_x_176_wall_t_out), .data_org(_add_map_x_176_data_org), .data_org_near(_add_map_x_176_data_org_near), .s_g(_add_map_x_176_s_g), .s_g_near(_add_map_x_176_s_g_near), .moto_org_near(_add_map_x_176_moto_org_near), .moto_org_near1(_add_map_x_176_moto_org_near1), .moto_org_near2(_add_map_x_176_moto_org_near2), .moto_org_near3(_add_map_x_176_moto_org_near3), .moto_org(_add_map_x_176_moto_org), .sg_up(_add_map_x_176_sg_up), .sg_down(_add_map_x_176_sg_down), .sg_left(_add_map_x_176_sg_left), .sg_right(_add_map_x_176_sg_right), .wall_t_in(_add_map_x_176_wall_t_in), .moto(_add_map_x_176_moto), .up(_add_map_x_176_up), .right(_add_map_x_176_right), .down(_add_map_x_176_down), .left(_add_map_x_176_left), .start(_add_map_x_176_start), .goal(_add_map_x_176_goal), .now(_add_map_x_176_now));
add_map add_map_x_175 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_175_add_exe), .data_out(_add_map_x_175_data_out), .data_out_index(_add_map_x_175_data_out_index), .data_near(_add_map_x_175_data_near), .wall_t_out(_add_map_x_175_wall_t_out), .data_org(_add_map_x_175_data_org), .data_org_near(_add_map_x_175_data_org_near), .s_g(_add_map_x_175_s_g), .s_g_near(_add_map_x_175_s_g_near), .moto_org_near(_add_map_x_175_moto_org_near), .moto_org_near1(_add_map_x_175_moto_org_near1), .moto_org_near2(_add_map_x_175_moto_org_near2), .moto_org_near3(_add_map_x_175_moto_org_near3), .moto_org(_add_map_x_175_moto_org), .sg_up(_add_map_x_175_sg_up), .sg_down(_add_map_x_175_sg_down), .sg_left(_add_map_x_175_sg_left), .sg_right(_add_map_x_175_sg_right), .wall_t_in(_add_map_x_175_wall_t_in), .moto(_add_map_x_175_moto), .up(_add_map_x_175_up), .right(_add_map_x_175_right), .down(_add_map_x_175_down), .left(_add_map_x_175_left), .start(_add_map_x_175_start), .goal(_add_map_x_175_goal), .now(_add_map_x_175_now));
add_map add_map_x_174 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_174_add_exe), .data_out(_add_map_x_174_data_out), .data_out_index(_add_map_x_174_data_out_index), .data_near(_add_map_x_174_data_near), .wall_t_out(_add_map_x_174_wall_t_out), .data_org(_add_map_x_174_data_org), .data_org_near(_add_map_x_174_data_org_near), .s_g(_add_map_x_174_s_g), .s_g_near(_add_map_x_174_s_g_near), .moto_org_near(_add_map_x_174_moto_org_near), .moto_org_near1(_add_map_x_174_moto_org_near1), .moto_org_near2(_add_map_x_174_moto_org_near2), .moto_org_near3(_add_map_x_174_moto_org_near3), .moto_org(_add_map_x_174_moto_org), .sg_up(_add_map_x_174_sg_up), .sg_down(_add_map_x_174_sg_down), .sg_left(_add_map_x_174_sg_left), .sg_right(_add_map_x_174_sg_right), .wall_t_in(_add_map_x_174_wall_t_in), .moto(_add_map_x_174_moto), .up(_add_map_x_174_up), .right(_add_map_x_174_right), .down(_add_map_x_174_down), .left(_add_map_x_174_left), .start(_add_map_x_174_start), .goal(_add_map_x_174_goal), .now(_add_map_x_174_now));
add_map add_map_x_173 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_173_add_exe), .data_out(_add_map_x_173_data_out), .data_out_index(_add_map_x_173_data_out_index), .data_near(_add_map_x_173_data_near), .wall_t_out(_add_map_x_173_wall_t_out), .data_org(_add_map_x_173_data_org), .data_org_near(_add_map_x_173_data_org_near), .s_g(_add_map_x_173_s_g), .s_g_near(_add_map_x_173_s_g_near), .moto_org_near(_add_map_x_173_moto_org_near), .moto_org_near1(_add_map_x_173_moto_org_near1), .moto_org_near2(_add_map_x_173_moto_org_near2), .moto_org_near3(_add_map_x_173_moto_org_near3), .moto_org(_add_map_x_173_moto_org), .sg_up(_add_map_x_173_sg_up), .sg_down(_add_map_x_173_sg_down), .sg_left(_add_map_x_173_sg_left), .sg_right(_add_map_x_173_sg_right), .wall_t_in(_add_map_x_173_wall_t_in), .moto(_add_map_x_173_moto), .up(_add_map_x_173_up), .right(_add_map_x_173_right), .down(_add_map_x_173_down), .left(_add_map_x_173_left), .start(_add_map_x_173_start), .goal(_add_map_x_173_goal), .now(_add_map_x_173_now));
add_map add_map_x_172 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_172_add_exe), .data_out(_add_map_x_172_data_out), .data_out_index(_add_map_x_172_data_out_index), .data_near(_add_map_x_172_data_near), .wall_t_out(_add_map_x_172_wall_t_out), .data_org(_add_map_x_172_data_org), .data_org_near(_add_map_x_172_data_org_near), .s_g(_add_map_x_172_s_g), .s_g_near(_add_map_x_172_s_g_near), .moto_org_near(_add_map_x_172_moto_org_near), .moto_org_near1(_add_map_x_172_moto_org_near1), .moto_org_near2(_add_map_x_172_moto_org_near2), .moto_org_near3(_add_map_x_172_moto_org_near3), .moto_org(_add_map_x_172_moto_org), .sg_up(_add_map_x_172_sg_up), .sg_down(_add_map_x_172_sg_down), .sg_left(_add_map_x_172_sg_left), .sg_right(_add_map_x_172_sg_right), .wall_t_in(_add_map_x_172_wall_t_in), .moto(_add_map_x_172_moto), .up(_add_map_x_172_up), .right(_add_map_x_172_right), .down(_add_map_x_172_down), .left(_add_map_x_172_left), .start(_add_map_x_172_start), .goal(_add_map_x_172_goal), .now(_add_map_x_172_now));
add_map add_map_x_171 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_171_add_exe), .data_out(_add_map_x_171_data_out), .data_out_index(_add_map_x_171_data_out_index), .data_near(_add_map_x_171_data_near), .wall_t_out(_add_map_x_171_wall_t_out), .data_org(_add_map_x_171_data_org), .data_org_near(_add_map_x_171_data_org_near), .s_g(_add_map_x_171_s_g), .s_g_near(_add_map_x_171_s_g_near), .moto_org_near(_add_map_x_171_moto_org_near), .moto_org_near1(_add_map_x_171_moto_org_near1), .moto_org_near2(_add_map_x_171_moto_org_near2), .moto_org_near3(_add_map_x_171_moto_org_near3), .moto_org(_add_map_x_171_moto_org), .sg_up(_add_map_x_171_sg_up), .sg_down(_add_map_x_171_sg_down), .sg_left(_add_map_x_171_sg_left), .sg_right(_add_map_x_171_sg_right), .wall_t_in(_add_map_x_171_wall_t_in), .moto(_add_map_x_171_moto), .up(_add_map_x_171_up), .right(_add_map_x_171_right), .down(_add_map_x_171_down), .left(_add_map_x_171_left), .start(_add_map_x_171_start), .goal(_add_map_x_171_goal), .now(_add_map_x_171_now));
add_map add_map_x_170 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_170_add_exe), .data_out(_add_map_x_170_data_out), .data_out_index(_add_map_x_170_data_out_index), .data_near(_add_map_x_170_data_near), .wall_t_out(_add_map_x_170_wall_t_out), .data_org(_add_map_x_170_data_org), .data_org_near(_add_map_x_170_data_org_near), .s_g(_add_map_x_170_s_g), .s_g_near(_add_map_x_170_s_g_near), .moto_org_near(_add_map_x_170_moto_org_near), .moto_org_near1(_add_map_x_170_moto_org_near1), .moto_org_near2(_add_map_x_170_moto_org_near2), .moto_org_near3(_add_map_x_170_moto_org_near3), .moto_org(_add_map_x_170_moto_org), .sg_up(_add_map_x_170_sg_up), .sg_down(_add_map_x_170_sg_down), .sg_left(_add_map_x_170_sg_left), .sg_right(_add_map_x_170_sg_right), .wall_t_in(_add_map_x_170_wall_t_in), .moto(_add_map_x_170_moto), .up(_add_map_x_170_up), .right(_add_map_x_170_right), .down(_add_map_x_170_down), .left(_add_map_x_170_left), .start(_add_map_x_170_start), .goal(_add_map_x_170_goal), .now(_add_map_x_170_now));
add_map add_map_x_169 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_169_add_exe), .data_out(_add_map_x_169_data_out), .data_out_index(_add_map_x_169_data_out_index), .data_near(_add_map_x_169_data_near), .wall_t_out(_add_map_x_169_wall_t_out), .data_org(_add_map_x_169_data_org), .data_org_near(_add_map_x_169_data_org_near), .s_g(_add_map_x_169_s_g), .s_g_near(_add_map_x_169_s_g_near), .moto_org_near(_add_map_x_169_moto_org_near), .moto_org_near1(_add_map_x_169_moto_org_near1), .moto_org_near2(_add_map_x_169_moto_org_near2), .moto_org_near3(_add_map_x_169_moto_org_near3), .moto_org(_add_map_x_169_moto_org), .sg_up(_add_map_x_169_sg_up), .sg_down(_add_map_x_169_sg_down), .sg_left(_add_map_x_169_sg_left), .sg_right(_add_map_x_169_sg_right), .wall_t_in(_add_map_x_169_wall_t_in), .moto(_add_map_x_169_moto), .up(_add_map_x_169_up), .right(_add_map_x_169_right), .down(_add_map_x_169_down), .left(_add_map_x_169_left), .start(_add_map_x_169_start), .goal(_add_map_x_169_goal), .now(_add_map_x_169_now));
add_map add_map_x_168 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_168_add_exe), .data_out(_add_map_x_168_data_out), .data_out_index(_add_map_x_168_data_out_index), .data_near(_add_map_x_168_data_near), .wall_t_out(_add_map_x_168_wall_t_out), .data_org(_add_map_x_168_data_org), .data_org_near(_add_map_x_168_data_org_near), .s_g(_add_map_x_168_s_g), .s_g_near(_add_map_x_168_s_g_near), .moto_org_near(_add_map_x_168_moto_org_near), .moto_org_near1(_add_map_x_168_moto_org_near1), .moto_org_near2(_add_map_x_168_moto_org_near2), .moto_org_near3(_add_map_x_168_moto_org_near3), .moto_org(_add_map_x_168_moto_org), .sg_up(_add_map_x_168_sg_up), .sg_down(_add_map_x_168_sg_down), .sg_left(_add_map_x_168_sg_left), .sg_right(_add_map_x_168_sg_right), .wall_t_in(_add_map_x_168_wall_t_in), .moto(_add_map_x_168_moto), .up(_add_map_x_168_up), .right(_add_map_x_168_right), .down(_add_map_x_168_down), .left(_add_map_x_168_left), .start(_add_map_x_168_start), .goal(_add_map_x_168_goal), .now(_add_map_x_168_now));
add_map add_map_x_167 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_167_add_exe), .data_out(_add_map_x_167_data_out), .data_out_index(_add_map_x_167_data_out_index), .data_near(_add_map_x_167_data_near), .wall_t_out(_add_map_x_167_wall_t_out), .data_org(_add_map_x_167_data_org), .data_org_near(_add_map_x_167_data_org_near), .s_g(_add_map_x_167_s_g), .s_g_near(_add_map_x_167_s_g_near), .moto_org_near(_add_map_x_167_moto_org_near), .moto_org_near1(_add_map_x_167_moto_org_near1), .moto_org_near2(_add_map_x_167_moto_org_near2), .moto_org_near3(_add_map_x_167_moto_org_near3), .moto_org(_add_map_x_167_moto_org), .sg_up(_add_map_x_167_sg_up), .sg_down(_add_map_x_167_sg_down), .sg_left(_add_map_x_167_sg_left), .sg_right(_add_map_x_167_sg_right), .wall_t_in(_add_map_x_167_wall_t_in), .moto(_add_map_x_167_moto), .up(_add_map_x_167_up), .right(_add_map_x_167_right), .down(_add_map_x_167_down), .left(_add_map_x_167_left), .start(_add_map_x_167_start), .goal(_add_map_x_167_goal), .now(_add_map_x_167_now));
add_map add_map_x_166 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_166_add_exe), .data_out(_add_map_x_166_data_out), .data_out_index(_add_map_x_166_data_out_index), .data_near(_add_map_x_166_data_near), .wall_t_out(_add_map_x_166_wall_t_out), .data_org(_add_map_x_166_data_org), .data_org_near(_add_map_x_166_data_org_near), .s_g(_add_map_x_166_s_g), .s_g_near(_add_map_x_166_s_g_near), .moto_org_near(_add_map_x_166_moto_org_near), .moto_org_near1(_add_map_x_166_moto_org_near1), .moto_org_near2(_add_map_x_166_moto_org_near2), .moto_org_near3(_add_map_x_166_moto_org_near3), .moto_org(_add_map_x_166_moto_org), .sg_up(_add_map_x_166_sg_up), .sg_down(_add_map_x_166_sg_down), .sg_left(_add_map_x_166_sg_left), .sg_right(_add_map_x_166_sg_right), .wall_t_in(_add_map_x_166_wall_t_in), .moto(_add_map_x_166_moto), .up(_add_map_x_166_up), .right(_add_map_x_166_right), .down(_add_map_x_166_down), .left(_add_map_x_166_left), .start(_add_map_x_166_start), .goal(_add_map_x_166_goal), .now(_add_map_x_166_now));
add_map add_map_x_165 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_165_add_exe), .data_out(_add_map_x_165_data_out), .data_out_index(_add_map_x_165_data_out_index), .data_near(_add_map_x_165_data_near), .wall_t_out(_add_map_x_165_wall_t_out), .data_org(_add_map_x_165_data_org), .data_org_near(_add_map_x_165_data_org_near), .s_g(_add_map_x_165_s_g), .s_g_near(_add_map_x_165_s_g_near), .moto_org_near(_add_map_x_165_moto_org_near), .moto_org_near1(_add_map_x_165_moto_org_near1), .moto_org_near2(_add_map_x_165_moto_org_near2), .moto_org_near3(_add_map_x_165_moto_org_near3), .moto_org(_add_map_x_165_moto_org), .sg_up(_add_map_x_165_sg_up), .sg_down(_add_map_x_165_sg_down), .sg_left(_add_map_x_165_sg_left), .sg_right(_add_map_x_165_sg_right), .wall_t_in(_add_map_x_165_wall_t_in), .moto(_add_map_x_165_moto), .up(_add_map_x_165_up), .right(_add_map_x_165_right), .down(_add_map_x_165_down), .left(_add_map_x_165_left), .start(_add_map_x_165_start), .goal(_add_map_x_165_goal), .now(_add_map_x_165_now));
add_map add_map_x_164 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_164_add_exe), .data_out(_add_map_x_164_data_out), .data_out_index(_add_map_x_164_data_out_index), .data_near(_add_map_x_164_data_near), .wall_t_out(_add_map_x_164_wall_t_out), .data_org(_add_map_x_164_data_org), .data_org_near(_add_map_x_164_data_org_near), .s_g(_add_map_x_164_s_g), .s_g_near(_add_map_x_164_s_g_near), .moto_org_near(_add_map_x_164_moto_org_near), .moto_org_near1(_add_map_x_164_moto_org_near1), .moto_org_near2(_add_map_x_164_moto_org_near2), .moto_org_near3(_add_map_x_164_moto_org_near3), .moto_org(_add_map_x_164_moto_org), .sg_up(_add_map_x_164_sg_up), .sg_down(_add_map_x_164_sg_down), .sg_left(_add_map_x_164_sg_left), .sg_right(_add_map_x_164_sg_right), .wall_t_in(_add_map_x_164_wall_t_in), .moto(_add_map_x_164_moto), .up(_add_map_x_164_up), .right(_add_map_x_164_right), .down(_add_map_x_164_down), .left(_add_map_x_164_left), .start(_add_map_x_164_start), .goal(_add_map_x_164_goal), .now(_add_map_x_164_now));
add_map add_map_x_163 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_163_add_exe), .data_out(_add_map_x_163_data_out), .data_out_index(_add_map_x_163_data_out_index), .data_near(_add_map_x_163_data_near), .wall_t_out(_add_map_x_163_wall_t_out), .data_org(_add_map_x_163_data_org), .data_org_near(_add_map_x_163_data_org_near), .s_g(_add_map_x_163_s_g), .s_g_near(_add_map_x_163_s_g_near), .moto_org_near(_add_map_x_163_moto_org_near), .moto_org_near1(_add_map_x_163_moto_org_near1), .moto_org_near2(_add_map_x_163_moto_org_near2), .moto_org_near3(_add_map_x_163_moto_org_near3), .moto_org(_add_map_x_163_moto_org), .sg_up(_add_map_x_163_sg_up), .sg_down(_add_map_x_163_sg_down), .sg_left(_add_map_x_163_sg_left), .sg_right(_add_map_x_163_sg_right), .wall_t_in(_add_map_x_163_wall_t_in), .moto(_add_map_x_163_moto), .up(_add_map_x_163_up), .right(_add_map_x_163_right), .down(_add_map_x_163_down), .left(_add_map_x_163_left), .start(_add_map_x_163_start), .goal(_add_map_x_163_goal), .now(_add_map_x_163_now));
add_map add_map_x_162 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_162_add_exe), .data_out(_add_map_x_162_data_out), .data_out_index(_add_map_x_162_data_out_index), .data_near(_add_map_x_162_data_near), .wall_t_out(_add_map_x_162_wall_t_out), .data_org(_add_map_x_162_data_org), .data_org_near(_add_map_x_162_data_org_near), .s_g(_add_map_x_162_s_g), .s_g_near(_add_map_x_162_s_g_near), .moto_org_near(_add_map_x_162_moto_org_near), .moto_org_near1(_add_map_x_162_moto_org_near1), .moto_org_near2(_add_map_x_162_moto_org_near2), .moto_org_near3(_add_map_x_162_moto_org_near3), .moto_org(_add_map_x_162_moto_org), .sg_up(_add_map_x_162_sg_up), .sg_down(_add_map_x_162_sg_down), .sg_left(_add_map_x_162_sg_left), .sg_right(_add_map_x_162_sg_right), .wall_t_in(_add_map_x_162_wall_t_in), .moto(_add_map_x_162_moto), .up(_add_map_x_162_up), .right(_add_map_x_162_right), .down(_add_map_x_162_down), .left(_add_map_x_162_left), .start(_add_map_x_162_start), .goal(_add_map_x_162_goal), .now(_add_map_x_162_now));
add_map add_map_x_161 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_161_add_exe), .data_out(_add_map_x_161_data_out), .data_out_index(_add_map_x_161_data_out_index), .data_near(_add_map_x_161_data_near), .wall_t_out(_add_map_x_161_wall_t_out), .data_org(_add_map_x_161_data_org), .data_org_near(_add_map_x_161_data_org_near), .s_g(_add_map_x_161_s_g), .s_g_near(_add_map_x_161_s_g_near), .moto_org_near(_add_map_x_161_moto_org_near), .moto_org_near1(_add_map_x_161_moto_org_near1), .moto_org_near2(_add_map_x_161_moto_org_near2), .moto_org_near3(_add_map_x_161_moto_org_near3), .moto_org(_add_map_x_161_moto_org), .sg_up(_add_map_x_161_sg_up), .sg_down(_add_map_x_161_sg_down), .sg_left(_add_map_x_161_sg_left), .sg_right(_add_map_x_161_sg_right), .wall_t_in(_add_map_x_161_wall_t_in), .moto(_add_map_x_161_moto), .up(_add_map_x_161_up), .right(_add_map_x_161_right), .down(_add_map_x_161_down), .left(_add_map_x_161_left), .start(_add_map_x_161_start), .goal(_add_map_x_161_goal), .now(_add_map_x_161_now));
add_map add_map_x_160 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_160_add_exe), .data_out(_add_map_x_160_data_out), .data_out_index(_add_map_x_160_data_out_index), .data_near(_add_map_x_160_data_near), .wall_t_out(_add_map_x_160_wall_t_out), .data_org(_add_map_x_160_data_org), .data_org_near(_add_map_x_160_data_org_near), .s_g(_add_map_x_160_s_g), .s_g_near(_add_map_x_160_s_g_near), .moto_org_near(_add_map_x_160_moto_org_near), .moto_org_near1(_add_map_x_160_moto_org_near1), .moto_org_near2(_add_map_x_160_moto_org_near2), .moto_org_near3(_add_map_x_160_moto_org_near3), .moto_org(_add_map_x_160_moto_org), .sg_up(_add_map_x_160_sg_up), .sg_down(_add_map_x_160_sg_down), .sg_left(_add_map_x_160_sg_left), .sg_right(_add_map_x_160_sg_right), .wall_t_in(_add_map_x_160_wall_t_in), .moto(_add_map_x_160_moto), .up(_add_map_x_160_up), .right(_add_map_x_160_right), .down(_add_map_x_160_down), .left(_add_map_x_160_left), .start(_add_map_x_160_start), .goal(_add_map_x_160_goal), .now(_add_map_x_160_now));
add_map add_map_x_159 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_159_add_exe), .data_out(_add_map_x_159_data_out), .data_out_index(_add_map_x_159_data_out_index), .data_near(_add_map_x_159_data_near), .wall_t_out(_add_map_x_159_wall_t_out), .data_org(_add_map_x_159_data_org), .data_org_near(_add_map_x_159_data_org_near), .s_g(_add_map_x_159_s_g), .s_g_near(_add_map_x_159_s_g_near), .moto_org_near(_add_map_x_159_moto_org_near), .moto_org_near1(_add_map_x_159_moto_org_near1), .moto_org_near2(_add_map_x_159_moto_org_near2), .moto_org_near3(_add_map_x_159_moto_org_near3), .moto_org(_add_map_x_159_moto_org), .sg_up(_add_map_x_159_sg_up), .sg_down(_add_map_x_159_sg_down), .sg_left(_add_map_x_159_sg_left), .sg_right(_add_map_x_159_sg_right), .wall_t_in(_add_map_x_159_wall_t_in), .moto(_add_map_x_159_moto), .up(_add_map_x_159_up), .right(_add_map_x_159_right), .down(_add_map_x_159_down), .left(_add_map_x_159_left), .start(_add_map_x_159_start), .goal(_add_map_x_159_goal), .now(_add_map_x_159_now));
add_map add_map_x_158 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_158_add_exe), .data_out(_add_map_x_158_data_out), .data_out_index(_add_map_x_158_data_out_index), .data_near(_add_map_x_158_data_near), .wall_t_out(_add_map_x_158_wall_t_out), .data_org(_add_map_x_158_data_org), .data_org_near(_add_map_x_158_data_org_near), .s_g(_add_map_x_158_s_g), .s_g_near(_add_map_x_158_s_g_near), .moto_org_near(_add_map_x_158_moto_org_near), .moto_org_near1(_add_map_x_158_moto_org_near1), .moto_org_near2(_add_map_x_158_moto_org_near2), .moto_org_near3(_add_map_x_158_moto_org_near3), .moto_org(_add_map_x_158_moto_org), .sg_up(_add_map_x_158_sg_up), .sg_down(_add_map_x_158_sg_down), .sg_left(_add_map_x_158_sg_left), .sg_right(_add_map_x_158_sg_right), .wall_t_in(_add_map_x_158_wall_t_in), .moto(_add_map_x_158_moto), .up(_add_map_x_158_up), .right(_add_map_x_158_right), .down(_add_map_x_158_down), .left(_add_map_x_158_left), .start(_add_map_x_158_start), .goal(_add_map_x_158_goal), .now(_add_map_x_158_now));
add_map add_map_x_157 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_157_add_exe), .data_out(_add_map_x_157_data_out), .data_out_index(_add_map_x_157_data_out_index), .data_near(_add_map_x_157_data_near), .wall_t_out(_add_map_x_157_wall_t_out), .data_org(_add_map_x_157_data_org), .data_org_near(_add_map_x_157_data_org_near), .s_g(_add_map_x_157_s_g), .s_g_near(_add_map_x_157_s_g_near), .moto_org_near(_add_map_x_157_moto_org_near), .moto_org_near1(_add_map_x_157_moto_org_near1), .moto_org_near2(_add_map_x_157_moto_org_near2), .moto_org_near3(_add_map_x_157_moto_org_near3), .moto_org(_add_map_x_157_moto_org), .sg_up(_add_map_x_157_sg_up), .sg_down(_add_map_x_157_sg_down), .sg_left(_add_map_x_157_sg_left), .sg_right(_add_map_x_157_sg_right), .wall_t_in(_add_map_x_157_wall_t_in), .moto(_add_map_x_157_moto), .up(_add_map_x_157_up), .right(_add_map_x_157_right), .down(_add_map_x_157_down), .left(_add_map_x_157_left), .start(_add_map_x_157_start), .goal(_add_map_x_157_goal), .now(_add_map_x_157_now));
add_map add_map_x_156 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_156_add_exe), .data_out(_add_map_x_156_data_out), .data_out_index(_add_map_x_156_data_out_index), .data_near(_add_map_x_156_data_near), .wall_t_out(_add_map_x_156_wall_t_out), .data_org(_add_map_x_156_data_org), .data_org_near(_add_map_x_156_data_org_near), .s_g(_add_map_x_156_s_g), .s_g_near(_add_map_x_156_s_g_near), .moto_org_near(_add_map_x_156_moto_org_near), .moto_org_near1(_add_map_x_156_moto_org_near1), .moto_org_near2(_add_map_x_156_moto_org_near2), .moto_org_near3(_add_map_x_156_moto_org_near3), .moto_org(_add_map_x_156_moto_org), .sg_up(_add_map_x_156_sg_up), .sg_down(_add_map_x_156_sg_down), .sg_left(_add_map_x_156_sg_left), .sg_right(_add_map_x_156_sg_right), .wall_t_in(_add_map_x_156_wall_t_in), .moto(_add_map_x_156_moto), .up(_add_map_x_156_up), .right(_add_map_x_156_right), .down(_add_map_x_156_down), .left(_add_map_x_156_left), .start(_add_map_x_156_start), .goal(_add_map_x_156_goal), .now(_add_map_x_156_now));
add_map add_map_x_155 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_155_add_exe), .data_out(_add_map_x_155_data_out), .data_out_index(_add_map_x_155_data_out_index), .data_near(_add_map_x_155_data_near), .wall_t_out(_add_map_x_155_wall_t_out), .data_org(_add_map_x_155_data_org), .data_org_near(_add_map_x_155_data_org_near), .s_g(_add_map_x_155_s_g), .s_g_near(_add_map_x_155_s_g_near), .moto_org_near(_add_map_x_155_moto_org_near), .moto_org_near1(_add_map_x_155_moto_org_near1), .moto_org_near2(_add_map_x_155_moto_org_near2), .moto_org_near3(_add_map_x_155_moto_org_near3), .moto_org(_add_map_x_155_moto_org), .sg_up(_add_map_x_155_sg_up), .sg_down(_add_map_x_155_sg_down), .sg_left(_add_map_x_155_sg_left), .sg_right(_add_map_x_155_sg_right), .wall_t_in(_add_map_x_155_wall_t_in), .moto(_add_map_x_155_moto), .up(_add_map_x_155_up), .right(_add_map_x_155_right), .down(_add_map_x_155_down), .left(_add_map_x_155_left), .start(_add_map_x_155_start), .goal(_add_map_x_155_goal), .now(_add_map_x_155_now));
add_map add_map_x_154 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_154_add_exe), .data_out(_add_map_x_154_data_out), .data_out_index(_add_map_x_154_data_out_index), .data_near(_add_map_x_154_data_near), .wall_t_out(_add_map_x_154_wall_t_out), .data_org(_add_map_x_154_data_org), .data_org_near(_add_map_x_154_data_org_near), .s_g(_add_map_x_154_s_g), .s_g_near(_add_map_x_154_s_g_near), .moto_org_near(_add_map_x_154_moto_org_near), .moto_org_near1(_add_map_x_154_moto_org_near1), .moto_org_near2(_add_map_x_154_moto_org_near2), .moto_org_near3(_add_map_x_154_moto_org_near3), .moto_org(_add_map_x_154_moto_org), .sg_up(_add_map_x_154_sg_up), .sg_down(_add_map_x_154_sg_down), .sg_left(_add_map_x_154_sg_left), .sg_right(_add_map_x_154_sg_right), .wall_t_in(_add_map_x_154_wall_t_in), .moto(_add_map_x_154_moto), .up(_add_map_x_154_up), .right(_add_map_x_154_right), .down(_add_map_x_154_down), .left(_add_map_x_154_left), .start(_add_map_x_154_start), .goal(_add_map_x_154_goal), .now(_add_map_x_154_now));
add_map add_map_x_153 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_153_add_exe), .data_out(_add_map_x_153_data_out), .data_out_index(_add_map_x_153_data_out_index), .data_near(_add_map_x_153_data_near), .wall_t_out(_add_map_x_153_wall_t_out), .data_org(_add_map_x_153_data_org), .data_org_near(_add_map_x_153_data_org_near), .s_g(_add_map_x_153_s_g), .s_g_near(_add_map_x_153_s_g_near), .moto_org_near(_add_map_x_153_moto_org_near), .moto_org_near1(_add_map_x_153_moto_org_near1), .moto_org_near2(_add_map_x_153_moto_org_near2), .moto_org_near3(_add_map_x_153_moto_org_near3), .moto_org(_add_map_x_153_moto_org), .sg_up(_add_map_x_153_sg_up), .sg_down(_add_map_x_153_sg_down), .sg_left(_add_map_x_153_sg_left), .sg_right(_add_map_x_153_sg_right), .wall_t_in(_add_map_x_153_wall_t_in), .moto(_add_map_x_153_moto), .up(_add_map_x_153_up), .right(_add_map_x_153_right), .down(_add_map_x_153_down), .left(_add_map_x_153_left), .start(_add_map_x_153_start), .goal(_add_map_x_153_goal), .now(_add_map_x_153_now));
add_map add_map_x_152 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_152_add_exe), .data_out(_add_map_x_152_data_out), .data_out_index(_add_map_x_152_data_out_index), .data_near(_add_map_x_152_data_near), .wall_t_out(_add_map_x_152_wall_t_out), .data_org(_add_map_x_152_data_org), .data_org_near(_add_map_x_152_data_org_near), .s_g(_add_map_x_152_s_g), .s_g_near(_add_map_x_152_s_g_near), .moto_org_near(_add_map_x_152_moto_org_near), .moto_org_near1(_add_map_x_152_moto_org_near1), .moto_org_near2(_add_map_x_152_moto_org_near2), .moto_org_near3(_add_map_x_152_moto_org_near3), .moto_org(_add_map_x_152_moto_org), .sg_up(_add_map_x_152_sg_up), .sg_down(_add_map_x_152_sg_down), .sg_left(_add_map_x_152_sg_left), .sg_right(_add_map_x_152_sg_right), .wall_t_in(_add_map_x_152_wall_t_in), .moto(_add_map_x_152_moto), .up(_add_map_x_152_up), .right(_add_map_x_152_right), .down(_add_map_x_152_down), .left(_add_map_x_152_left), .start(_add_map_x_152_start), .goal(_add_map_x_152_goal), .now(_add_map_x_152_now));
add_map add_map_x_151 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_151_add_exe), .data_out(_add_map_x_151_data_out), .data_out_index(_add_map_x_151_data_out_index), .data_near(_add_map_x_151_data_near), .wall_t_out(_add_map_x_151_wall_t_out), .data_org(_add_map_x_151_data_org), .data_org_near(_add_map_x_151_data_org_near), .s_g(_add_map_x_151_s_g), .s_g_near(_add_map_x_151_s_g_near), .moto_org_near(_add_map_x_151_moto_org_near), .moto_org_near1(_add_map_x_151_moto_org_near1), .moto_org_near2(_add_map_x_151_moto_org_near2), .moto_org_near3(_add_map_x_151_moto_org_near3), .moto_org(_add_map_x_151_moto_org), .sg_up(_add_map_x_151_sg_up), .sg_down(_add_map_x_151_sg_down), .sg_left(_add_map_x_151_sg_left), .sg_right(_add_map_x_151_sg_right), .wall_t_in(_add_map_x_151_wall_t_in), .moto(_add_map_x_151_moto), .up(_add_map_x_151_up), .right(_add_map_x_151_right), .down(_add_map_x_151_down), .left(_add_map_x_151_left), .start(_add_map_x_151_start), .goal(_add_map_x_151_goal), .now(_add_map_x_151_now));
add_map add_map_x_150 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_150_add_exe), .data_out(_add_map_x_150_data_out), .data_out_index(_add_map_x_150_data_out_index), .data_near(_add_map_x_150_data_near), .wall_t_out(_add_map_x_150_wall_t_out), .data_org(_add_map_x_150_data_org), .data_org_near(_add_map_x_150_data_org_near), .s_g(_add_map_x_150_s_g), .s_g_near(_add_map_x_150_s_g_near), .moto_org_near(_add_map_x_150_moto_org_near), .moto_org_near1(_add_map_x_150_moto_org_near1), .moto_org_near2(_add_map_x_150_moto_org_near2), .moto_org_near3(_add_map_x_150_moto_org_near3), .moto_org(_add_map_x_150_moto_org), .sg_up(_add_map_x_150_sg_up), .sg_down(_add_map_x_150_sg_down), .sg_left(_add_map_x_150_sg_left), .sg_right(_add_map_x_150_sg_right), .wall_t_in(_add_map_x_150_wall_t_in), .moto(_add_map_x_150_moto), .up(_add_map_x_150_up), .right(_add_map_x_150_right), .down(_add_map_x_150_down), .left(_add_map_x_150_left), .start(_add_map_x_150_start), .goal(_add_map_x_150_goal), .now(_add_map_x_150_now));
add_map add_map_x_149 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_149_add_exe), .data_out(_add_map_x_149_data_out), .data_out_index(_add_map_x_149_data_out_index), .data_near(_add_map_x_149_data_near), .wall_t_out(_add_map_x_149_wall_t_out), .data_org(_add_map_x_149_data_org), .data_org_near(_add_map_x_149_data_org_near), .s_g(_add_map_x_149_s_g), .s_g_near(_add_map_x_149_s_g_near), .moto_org_near(_add_map_x_149_moto_org_near), .moto_org_near1(_add_map_x_149_moto_org_near1), .moto_org_near2(_add_map_x_149_moto_org_near2), .moto_org_near3(_add_map_x_149_moto_org_near3), .moto_org(_add_map_x_149_moto_org), .sg_up(_add_map_x_149_sg_up), .sg_down(_add_map_x_149_sg_down), .sg_left(_add_map_x_149_sg_left), .sg_right(_add_map_x_149_sg_right), .wall_t_in(_add_map_x_149_wall_t_in), .moto(_add_map_x_149_moto), .up(_add_map_x_149_up), .right(_add_map_x_149_right), .down(_add_map_x_149_down), .left(_add_map_x_149_left), .start(_add_map_x_149_start), .goal(_add_map_x_149_goal), .now(_add_map_x_149_now));
add_map add_map_x_148 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_148_add_exe), .data_out(_add_map_x_148_data_out), .data_out_index(_add_map_x_148_data_out_index), .data_near(_add_map_x_148_data_near), .wall_t_out(_add_map_x_148_wall_t_out), .data_org(_add_map_x_148_data_org), .data_org_near(_add_map_x_148_data_org_near), .s_g(_add_map_x_148_s_g), .s_g_near(_add_map_x_148_s_g_near), .moto_org_near(_add_map_x_148_moto_org_near), .moto_org_near1(_add_map_x_148_moto_org_near1), .moto_org_near2(_add_map_x_148_moto_org_near2), .moto_org_near3(_add_map_x_148_moto_org_near3), .moto_org(_add_map_x_148_moto_org), .sg_up(_add_map_x_148_sg_up), .sg_down(_add_map_x_148_sg_down), .sg_left(_add_map_x_148_sg_left), .sg_right(_add_map_x_148_sg_right), .wall_t_in(_add_map_x_148_wall_t_in), .moto(_add_map_x_148_moto), .up(_add_map_x_148_up), .right(_add_map_x_148_right), .down(_add_map_x_148_down), .left(_add_map_x_148_left), .start(_add_map_x_148_start), .goal(_add_map_x_148_goal), .now(_add_map_x_148_now));
add_map add_map_x_147 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_147_add_exe), .data_out(_add_map_x_147_data_out), .data_out_index(_add_map_x_147_data_out_index), .data_near(_add_map_x_147_data_near), .wall_t_out(_add_map_x_147_wall_t_out), .data_org(_add_map_x_147_data_org), .data_org_near(_add_map_x_147_data_org_near), .s_g(_add_map_x_147_s_g), .s_g_near(_add_map_x_147_s_g_near), .moto_org_near(_add_map_x_147_moto_org_near), .moto_org_near1(_add_map_x_147_moto_org_near1), .moto_org_near2(_add_map_x_147_moto_org_near2), .moto_org_near3(_add_map_x_147_moto_org_near3), .moto_org(_add_map_x_147_moto_org), .sg_up(_add_map_x_147_sg_up), .sg_down(_add_map_x_147_sg_down), .sg_left(_add_map_x_147_sg_left), .sg_right(_add_map_x_147_sg_right), .wall_t_in(_add_map_x_147_wall_t_in), .moto(_add_map_x_147_moto), .up(_add_map_x_147_up), .right(_add_map_x_147_right), .down(_add_map_x_147_down), .left(_add_map_x_147_left), .start(_add_map_x_147_start), .goal(_add_map_x_147_goal), .now(_add_map_x_147_now));
add_map add_map_x_146 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_146_add_exe), .data_out(_add_map_x_146_data_out), .data_out_index(_add_map_x_146_data_out_index), .data_near(_add_map_x_146_data_near), .wall_t_out(_add_map_x_146_wall_t_out), .data_org(_add_map_x_146_data_org), .data_org_near(_add_map_x_146_data_org_near), .s_g(_add_map_x_146_s_g), .s_g_near(_add_map_x_146_s_g_near), .moto_org_near(_add_map_x_146_moto_org_near), .moto_org_near1(_add_map_x_146_moto_org_near1), .moto_org_near2(_add_map_x_146_moto_org_near2), .moto_org_near3(_add_map_x_146_moto_org_near3), .moto_org(_add_map_x_146_moto_org), .sg_up(_add_map_x_146_sg_up), .sg_down(_add_map_x_146_sg_down), .sg_left(_add_map_x_146_sg_left), .sg_right(_add_map_x_146_sg_right), .wall_t_in(_add_map_x_146_wall_t_in), .moto(_add_map_x_146_moto), .up(_add_map_x_146_up), .right(_add_map_x_146_right), .down(_add_map_x_146_down), .left(_add_map_x_146_left), .start(_add_map_x_146_start), .goal(_add_map_x_146_goal), .now(_add_map_x_146_now));
add_map add_map_x_145 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_145_add_exe), .data_out(_add_map_x_145_data_out), .data_out_index(_add_map_x_145_data_out_index), .data_near(_add_map_x_145_data_near), .wall_t_out(_add_map_x_145_wall_t_out), .data_org(_add_map_x_145_data_org), .data_org_near(_add_map_x_145_data_org_near), .s_g(_add_map_x_145_s_g), .s_g_near(_add_map_x_145_s_g_near), .moto_org_near(_add_map_x_145_moto_org_near), .moto_org_near1(_add_map_x_145_moto_org_near1), .moto_org_near2(_add_map_x_145_moto_org_near2), .moto_org_near3(_add_map_x_145_moto_org_near3), .moto_org(_add_map_x_145_moto_org), .sg_up(_add_map_x_145_sg_up), .sg_down(_add_map_x_145_sg_down), .sg_left(_add_map_x_145_sg_left), .sg_right(_add_map_x_145_sg_right), .wall_t_in(_add_map_x_145_wall_t_in), .moto(_add_map_x_145_moto), .up(_add_map_x_145_up), .right(_add_map_x_145_right), .down(_add_map_x_145_down), .left(_add_map_x_145_left), .start(_add_map_x_145_start), .goal(_add_map_x_145_goal), .now(_add_map_x_145_now));
add_map add_map_x_144 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_144_add_exe), .data_out(_add_map_x_144_data_out), .data_out_index(_add_map_x_144_data_out_index), .data_near(_add_map_x_144_data_near), .wall_t_out(_add_map_x_144_wall_t_out), .data_org(_add_map_x_144_data_org), .data_org_near(_add_map_x_144_data_org_near), .s_g(_add_map_x_144_s_g), .s_g_near(_add_map_x_144_s_g_near), .moto_org_near(_add_map_x_144_moto_org_near), .moto_org_near1(_add_map_x_144_moto_org_near1), .moto_org_near2(_add_map_x_144_moto_org_near2), .moto_org_near3(_add_map_x_144_moto_org_near3), .moto_org(_add_map_x_144_moto_org), .sg_up(_add_map_x_144_sg_up), .sg_down(_add_map_x_144_sg_down), .sg_left(_add_map_x_144_sg_left), .sg_right(_add_map_x_144_sg_right), .wall_t_in(_add_map_x_144_wall_t_in), .moto(_add_map_x_144_moto), .up(_add_map_x_144_up), .right(_add_map_x_144_right), .down(_add_map_x_144_down), .left(_add_map_x_144_left), .start(_add_map_x_144_start), .goal(_add_map_x_144_goal), .now(_add_map_x_144_now));
add_map add_map_x_143 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_143_add_exe), .data_out(_add_map_x_143_data_out), .data_out_index(_add_map_x_143_data_out_index), .data_near(_add_map_x_143_data_near), .wall_t_out(_add_map_x_143_wall_t_out), .data_org(_add_map_x_143_data_org), .data_org_near(_add_map_x_143_data_org_near), .s_g(_add_map_x_143_s_g), .s_g_near(_add_map_x_143_s_g_near), .moto_org_near(_add_map_x_143_moto_org_near), .moto_org_near1(_add_map_x_143_moto_org_near1), .moto_org_near2(_add_map_x_143_moto_org_near2), .moto_org_near3(_add_map_x_143_moto_org_near3), .moto_org(_add_map_x_143_moto_org), .sg_up(_add_map_x_143_sg_up), .sg_down(_add_map_x_143_sg_down), .sg_left(_add_map_x_143_sg_left), .sg_right(_add_map_x_143_sg_right), .wall_t_in(_add_map_x_143_wall_t_in), .moto(_add_map_x_143_moto), .up(_add_map_x_143_up), .right(_add_map_x_143_right), .down(_add_map_x_143_down), .left(_add_map_x_143_left), .start(_add_map_x_143_start), .goal(_add_map_x_143_goal), .now(_add_map_x_143_now));
add_map add_map_x_142 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_142_add_exe), .data_out(_add_map_x_142_data_out), .data_out_index(_add_map_x_142_data_out_index), .data_near(_add_map_x_142_data_near), .wall_t_out(_add_map_x_142_wall_t_out), .data_org(_add_map_x_142_data_org), .data_org_near(_add_map_x_142_data_org_near), .s_g(_add_map_x_142_s_g), .s_g_near(_add_map_x_142_s_g_near), .moto_org_near(_add_map_x_142_moto_org_near), .moto_org_near1(_add_map_x_142_moto_org_near1), .moto_org_near2(_add_map_x_142_moto_org_near2), .moto_org_near3(_add_map_x_142_moto_org_near3), .moto_org(_add_map_x_142_moto_org), .sg_up(_add_map_x_142_sg_up), .sg_down(_add_map_x_142_sg_down), .sg_left(_add_map_x_142_sg_left), .sg_right(_add_map_x_142_sg_right), .wall_t_in(_add_map_x_142_wall_t_in), .moto(_add_map_x_142_moto), .up(_add_map_x_142_up), .right(_add_map_x_142_right), .down(_add_map_x_142_down), .left(_add_map_x_142_left), .start(_add_map_x_142_start), .goal(_add_map_x_142_goal), .now(_add_map_x_142_now));
add_map add_map_x_141 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_141_add_exe), .data_out(_add_map_x_141_data_out), .data_out_index(_add_map_x_141_data_out_index), .data_near(_add_map_x_141_data_near), .wall_t_out(_add_map_x_141_wall_t_out), .data_org(_add_map_x_141_data_org), .data_org_near(_add_map_x_141_data_org_near), .s_g(_add_map_x_141_s_g), .s_g_near(_add_map_x_141_s_g_near), .moto_org_near(_add_map_x_141_moto_org_near), .moto_org_near1(_add_map_x_141_moto_org_near1), .moto_org_near2(_add_map_x_141_moto_org_near2), .moto_org_near3(_add_map_x_141_moto_org_near3), .moto_org(_add_map_x_141_moto_org), .sg_up(_add_map_x_141_sg_up), .sg_down(_add_map_x_141_sg_down), .sg_left(_add_map_x_141_sg_left), .sg_right(_add_map_x_141_sg_right), .wall_t_in(_add_map_x_141_wall_t_in), .moto(_add_map_x_141_moto), .up(_add_map_x_141_up), .right(_add_map_x_141_right), .down(_add_map_x_141_down), .left(_add_map_x_141_left), .start(_add_map_x_141_start), .goal(_add_map_x_141_goal), .now(_add_map_x_141_now));
add_map add_map_x_140 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_140_add_exe), .data_out(_add_map_x_140_data_out), .data_out_index(_add_map_x_140_data_out_index), .data_near(_add_map_x_140_data_near), .wall_t_out(_add_map_x_140_wall_t_out), .data_org(_add_map_x_140_data_org), .data_org_near(_add_map_x_140_data_org_near), .s_g(_add_map_x_140_s_g), .s_g_near(_add_map_x_140_s_g_near), .moto_org_near(_add_map_x_140_moto_org_near), .moto_org_near1(_add_map_x_140_moto_org_near1), .moto_org_near2(_add_map_x_140_moto_org_near2), .moto_org_near3(_add_map_x_140_moto_org_near3), .moto_org(_add_map_x_140_moto_org), .sg_up(_add_map_x_140_sg_up), .sg_down(_add_map_x_140_sg_down), .sg_left(_add_map_x_140_sg_left), .sg_right(_add_map_x_140_sg_right), .wall_t_in(_add_map_x_140_wall_t_in), .moto(_add_map_x_140_moto), .up(_add_map_x_140_up), .right(_add_map_x_140_right), .down(_add_map_x_140_down), .left(_add_map_x_140_left), .start(_add_map_x_140_start), .goal(_add_map_x_140_goal), .now(_add_map_x_140_now));
add_map add_map_x_139 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_139_add_exe), .data_out(_add_map_x_139_data_out), .data_out_index(_add_map_x_139_data_out_index), .data_near(_add_map_x_139_data_near), .wall_t_out(_add_map_x_139_wall_t_out), .data_org(_add_map_x_139_data_org), .data_org_near(_add_map_x_139_data_org_near), .s_g(_add_map_x_139_s_g), .s_g_near(_add_map_x_139_s_g_near), .moto_org_near(_add_map_x_139_moto_org_near), .moto_org_near1(_add_map_x_139_moto_org_near1), .moto_org_near2(_add_map_x_139_moto_org_near2), .moto_org_near3(_add_map_x_139_moto_org_near3), .moto_org(_add_map_x_139_moto_org), .sg_up(_add_map_x_139_sg_up), .sg_down(_add_map_x_139_sg_down), .sg_left(_add_map_x_139_sg_left), .sg_right(_add_map_x_139_sg_right), .wall_t_in(_add_map_x_139_wall_t_in), .moto(_add_map_x_139_moto), .up(_add_map_x_139_up), .right(_add_map_x_139_right), .down(_add_map_x_139_down), .left(_add_map_x_139_left), .start(_add_map_x_139_start), .goal(_add_map_x_139_goal), .now(_add_map_x_139_now));
add_map add_map_x_138 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_138_add_exe), .data_out(_add_map_x_138_data_out), .data_out_index(_add_map_x_138_data_out_index), .data_near(_add_map_x_138_data_near), .wall_t_out(_add_map_x_138_wall_t_out), .data_org(_add_map_x_138_data_org), .data_org_near(_add_map_x_138_data_org_near), .s_g(_add_map_x_138_s_g), .s_g_near(_add_map_x_138_s_g_near), .moto_org_near(_add_map_x_138_moto_org_near), .moto_org_near1(_add_map_x_138_moto_org_near1), .moto_org_near2(_add_map_x_138_moto_org_near2), .moto_org_near3(_add_map_x_138_moto_org_near3), .moto_org(_add_map_x_138_moto_org), .sg_up(_add_map_x_138_sg_up), .sg_down(_add_map_x_138_sg_down), .sg_left(_add_map_x_138_sg_left), .sg_right(_add_map_x_138_sg_right), .wall_t_in(_add_map_x_138_wall_t_in), .moto(_add_map_x_138_moto), .up(_add_map_x_138_up), .right(_add_map_x_138_right), .down(_add_map_x_138_down), .left(_add_map_x_138_left), .start(_add_map_x_138_start), .goal(_add_map_x_138_goal), .now(_add_map_x_138_now));
add_map add_map_x_137 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_137_add_exe), .data_out(_add_map_x_137_data_out), .data_out_index(_add_map_x_137_data_out_index), .data_near(_add_map_x_137_data_near), .wall_t_out(_add_map_x_137_wall_t_out), .data_org(_add_map_x_137_data_org), .data_org_near(_add_map_x_137_data_org_near), .s_g(_add_map_x_137_s_g), .s_g_near(_add_map_x_137_s_g_near), .moto_org_near(_add_map_x_137_moto_org_near), .moto_org_near1(_add_map_x_137_moto_org_near1), .moto_org_near2(_add_map_x_137_moto_org_near2), .moto_org_near3(_add_map_x_137_moto_org_near3), .moto_org(_add_map_x_137_moto_org), .sg_up(_add_map_x_137_sg_up), .sg_down(_add_map_x_137_sg_down), .sg_left(_add_map_x_137_sg_left), .sg_right(_add_map_x_137_sg_right), .wall_t_in(_add_map_x_137_wall_t_in), .moto(_add_map_x_137_moto), .up(_add_map_x_137_up), .right(_add_map_x_137_right), .down(_add_map_x_137_down), .left(_add_map_x_137_left), .start(_add_map_x_137_start), .goal(_add_map_x_137_goal), .now(_add_map_x_137_now));
add_map add_map_x_136 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_136_add_exe), .data_out(_add_map_x_136_data_out), .data_out_index(_add_map_x_136_data_out_index), .data_near(_add_map_x_136_data_near), .wall_t_out(_add_map_x_136_wall_t_out), .data_org(_add_map_x_136_data_org), .data_org_near(_add_map_x_136_data_org_near), .s_g(_add_map_x_136_s_g), .s_g_near(_add_map_x_136_s_g_near), .moto_org_near(_add_map_x_136_moto_org_near), .moto_org_near1(_add_map_x_136_moto_org_near1), .moto_org_near2(_add_map_x_136_moto_org_near2), .moto_org_near3(_add_map_x_136_moto_org_near3), .moto_org(_add_map_x_136_moto_org), .sg_up(_add_map_x_136_sg_up), .sg_down(_add_map_x_136_sg_down), .sg_left(_add_map_x_136_sg_left), .sg_right(_add_map_x_136_sg_right), .wall_t_in(_add_map_x_136_wall_t_in), .moto(_add_map_x_136_moto), .up(_add_map_x_136_up), .right(_add_map_x_136_right), .down(_add_map_x_136_down), .left(_add_map_x_136_left), .start(_add_map_x_136_start), .goal(_add_map_x_136_goal), .now(_add_map_x_136_now));
add_map add_map_x_135 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_135_add_exe), .data_out(_add_map_x_135_data_out), .data_out_index(_add_map_x_135_data_out_index), .data_near(_add_map_x_135_data_near), .wall_t_out(_add_map_x_135_wall_t_out), .data_org(_add_map_x_135_data_org), .data_org_near(_add_map_x_135_data_org_near), .s_g(_add_map_x_135_s_g), .s_g_near(_add_map_x_135_s_g_near), .moto_org_near(_add_map_x_135_moto_org_near), .moto_org_near1(_add_map_x_135_moto_org_near1), .moto_org_near2(_add_map_x_135_moto_org_near2), .moto_org_near3(_add_map_x_135_moto_org_near3), .moto_org(_add_map_x_135_moto_org), .sg_up(_add_map_x_135_sg_up), .sg_down(_add_map_x_135_sg_down), .sg_left(_add_map_x_135_sg_left), .sg_right(_add_map_x_135_sg_right), .wall_t_in(_add_map_x_135_wall_t_in), .moto(_add_map_x_135_moto), .up(_add_map_x_135_up), .right(_add_map_x_135_right), .down(_add_map_x_135_down), .left(_add_map_x_135_left), .start(_add_map_x_135_start), .goal(_add_map_x_135_goal), .now(_add_map_x_135_now));
add_map add_map_x_134 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_134_add_exe), .data_out(_add_map_x_134_data_out), .data_out_index(_add_map_x_134_data_out_index), .data_near(_add_map_x_134_data_near), .wall_t_out(_add_map_x_134_wall_t_out), .data_org(_add_map_x_134_data_org), .data_org_near(_add_map_x_134_data_org_near), .s_g(_add_map_x_134_s_g), .s_g_near(_add_map_x_134_s_g_near), .moto_org_near(_add_map_x_134_moto_org_near), .moto_org_near1(_add_map_x_134_moto_org_near1), .moto_org_near2(_add_map_x_134_moto_org_near2), .moto_org_near3(_add_map_x_134_moto_org_near3), .moto_org(_add_map_x_134_moto_org), .sg_up(_add_map_x_134_sg_up), .sg_down(_add_map_x_134_sg_down), .sg_left(_add_map_x_134_sg_left), .sg_right(_add_map_x_134_sg_right), .wall_t_in(_add_map_x_134_wall_t_in), .moto(_add_map_x_134_moto), .up(_add_map_x_134_up), .right(_add_map_x_134_right), .down(_add_map_x_134_down), .left(_add_map_x_134_left), .start(_add_map_x_134_start), .goal(_add_map_x_134_goal), .now(_add_map_x_134_now));
add_map add_map_x_133 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_133_add_exe), .data_out(_add_map_x_133_data_out), .data_out_index(_add_map_x_133_data_out_index), .data_near(_add_map_x_133_data_near), .wall_t_out(_add_map_x_133_wall_t_out), .data_org(_add_map_x_133_data_org), .data_org_near(_add_map_x_133_data_org_near), .s_g(_add_map_x_133_s_g), .s_g_near(_add_map_x_133_s_g_near), .moto_org_near(_add_map_x_133_moto_org_near), .moto_org_near1(_add_map_x_133_moto_org_near1), .moto_org_near2(_add_map_x_133_moto_org_near2), .moto_org_near3(_add_map_x_133_moto_org_near3), .moto_org(_add_map_x_133_moto_org), .sg_up(_add_map_x_133_sg_up), .sg_down(_add_map_x_133_sg_down), .sg_left(_add_map_x_133_sg_left), .sg_right(_add_map_x_133_sg_right), .wall_t_in(_add_map_x_133_wall_t_in), .moto(_add_map_x_133_moto), .up(_add_map_x_133_up), .right(_add_map_x_133_right), .down(_add_map_x_133_down), .left(_add_map_x_133_left), .start(_add_map_x_133_start), .goal(_add_map_x_133_goal), .now(_add_map_x_133_now));
add_map add_map_x_132 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_132_add_exe), .data_out(_add_map_x_132_data_out), .data_out_index(_add_map_x_132_data_out_index), .data_near(_add_map_x_132_data_near), .wall_t_out(_add_map_x_132_wall_t_out), .data_org(_add_map_x_132_data_org), .data_org_near(_add_map_x_132_data_org_near), .s_g(_add_map_x_132_s_g), .s_g_near(_add_map_x_132_s_g_near), .moto_org_near(_add_map_x_132_moto_org_near), .moto_org_near1(_add_map_x_132_moto_org_near1), .moto_org_near2(_add_map_x_132_moto_org_near2), .moto_org_near3(_add_map_x_132_moto_org_near3), .moto_org(_add_map_x_132_moto_org), .sg_up(_add_map_x_132_sg_up), .sg_down(_add_map_x_132_sg_down), .sg_left(_add_map_x_132_sg_left), .sg_right(_add_map_x_132_sg_right), .wall_t_in(_add_map_x_132_wall_t_in), .moto(_add_map_x_132_moto), .up(_add_map_x_132_up), .right(_add_map_x_132_right), .down(_add_map_x_132_down), .left(_add_map_x_132_left), .start(_add_map_x_132_start), .goal(_add_map_x_132_goal), .now(_add_map_x_132_now));
add_map add_map_x_131 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_131_add_exe), .data_out(_add_map_x_131_data_out), .data_out_index(_add_map_x_131_data_out_index), .data_near(_add_map_x_131_data_near), .wall_t_out(_add_map_x_131_wall_t_out), .data_org(_add_map_x_131_data_org), .data_org_near(_add_map_x_131_data_org_near), .s_g(_add_map_x_131_s_g), .s_g_near(_add_map_x_131_s_g_near), .moto_org_near(_add_map_x_131_moto_org_near), .moto_org_near1(_add_map_x_131_moto_org_near1), .moto_org_near2(_add_map_x_131_moto_org_near2), .moto_org_near3(_add_map_x_131_moto_org_near3), .moto_org(_add_map_x_131_moto_org), .sg_up(_add_map_x_131_sg_up), .sg_down(_add_map_x_131_sg_down), .sg_left(_add_map_x_131_sg_left), .sg_right(_add_map_x_131_sg_right), .wall_t_in(_add_map_x_131_wall_t_in), .moto(_add_map_x_131_moto), .up(_add_map_x_131_up), .right(_add_map_x_131_right), .down(_add_map_x_131_down), .left(_add_map_x_131_left), .start(_add_map_x_131_start), .goal(_add_map_x_131_goal), .now(_add_map_x_131_now));
add_map add_map_x_130 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_130_add_exe), .data_out(_add_map_x_130_data_out), .data_out_index(_add_map_x_130_data_out_index), .data_near(_add_map_x_130_data_near), .wall_t_out(_add_map_x_130_wall_t_out), .data_org(_add_map_x_130_data_org), .data_org_near(_add_map_x_130_data_org_near), .s_g(_add_map_x_130_s_g), .s_g_near(_add_map_x_130_s_g_near), .moto_org_near(_add_map_x_130_moto_org_near), .moto_org_near1(_add_map_x_130_moto_org_near1), .moto_org_near2(_add_map_x_130_moto_org_near2), .moto_org_near3(_add_map_x_130_moto_org_near3), .moto_org(_add_map_x_130_moto_org), .sg_up(_add_map_x_130_sg_up), .sg_down(_add_map_x_130_sg_down), .sg_left(_add_map_x_130_sg_left), .sg_right(_add_map_x_130_sg_right), .wall_t_in(_add_map_x_130_wall_t_in), .moto(_add_map_x_130_moto), .up(_add_map_x_130_up), .right(_add_map_x_130_right), .down(_add_map_x_130_down), .left(_add_map_x_130_left), .start(_add_map_x_130_start), .goal(_add_map_x_130_goal), .now(_add_map_x_130_now));
add_map add_map_x_129 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_129_add_exe), .data_out(_add_map_x_129_data_out), .data_out_index(_add_map_x_129_data_out_index), .data_near(_add_map_x_129_data_near), .wall_t_out(_add_map_x_129_wall_t_out), .data_org(_add_map_x_129_data_org), .data_org_near(_add_map_x_129_data_org_near), .s_g(_add_map_x_129_s_g), .s_g_near(_add_map_x_129_s_g_near), .moto_org_near(_add_map_x_129_moto_org_near), .moto_org_near1(_add_map_x_129_moto_org_near1), .moto_org_near2(_add_map_x_129_moto_org_near2), .moto_org_near3(_add_map_x_129_moto_org_near3), .moto_org(_add_map_x_129_moto_org), .sg_up(_add_map_x_129_sg_up), .sg_down(_add_map_x_129_sg_down), .sg_left(_add_map_x_129_sg_left), .sg_right(_add_map_x_129_sg_right), .wall_t_in(_add_map_x_129_wall_t_in), .moto(_add_map_x_129_moto), .up(_add_map_x_129_up), .right(_add_map_x_129_right), .down(_add_map_x_129_down), .left(_add_map_x_129_left), .start(_add_map_x_129_start), .goal(_add_map_x_129_goal), .now(_add_map_x_129_now));
add_map add_map_x_128 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_128_add_exe), .data_out(_add_map_x_128_data_out), .data_out_index(_add_map_x_128_data_out_index), .data_near(_add_map_x_128_data_near), .wall_t_out(_add_map_x_128_wall_t_out), .data_org(_add_map_x_128_data_org), .data_org_near(_add_map_x_128_data_org_near), .s_g(_add_map_x_128_s_g), .s_g_near(_add_map_x_128_s_g_near), .moto_org_near(_add_map_x_128_moto_org_near), .moto_org_near1(_add_map_x_128_moto_org_near1), .moto_org_near2(_add_map_x_128_moto_org_near2), .moto_org_near3(_add_map_x_128_moto_org_near3), .moto_org(_add_map_x_128_moto_org), .sg_up(_add_map_x_128_sg_up), .sg_down(_add_map_x_128_sg_down), .sg_left(_add_map_x_128_sg_left), .sg_right(_add_map_x_128_sg_right), .wall_t_in(_add_map_x_128_wall_t_in), .moto(_add_map_x_128_moto), .up(_add_map_x_128_up), .right(_add_map_x_128_right), .down(_add_map_x_128_down), .left(_add_map_x_128_left), .start(_add_map_x_128_start), .goal(_add_map_x_128_goal), .now(_add_map_x_128_now));
add_map add_map_x_127 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_127_add_exe), .data_out(_add_map_x_127_data_out), .data_out_index(_add_map_x_127_data_out_index), .data_near(_add_map_x_127_data_near), .wall_t_out(_add_map_x_127_wall_t_out), .data_org(_add_map_x_127_data_org), .data_org_near(_add_map_x_127_data_org_near), .s_g(_add_map_x_127_s_g), .s_g_near(_add_map_x_127_s_g_near), .moto_org_near(_add_map_x_127_moto_org_near), .moto_org_near1(_add_map_x_127_moto_org_near1), .moto_org_near2(_add_map_x_127_moto_org_near2), .moto_org_near3(_add_map_x_127_moto_org_near3), .moto_org(_add_map_x_127_moto_org), .sg_up(_add_map_x_127_sg_up), .sg_down(_add_map_x_127_sg_down), .sg_left(_add_map_x_127_sg_left), .sg_right(_add_map_x_127_sg_right), .wall_t_in(_add_map_x_127_wall_t_in), .moto(_add_map_x_127_moto), .up(_add_map_x_127_up), .right(_add_map_x_127_right), .down(_add_map_x_127_down), .left(_add_map_x_127_left), .start(_add_map_x_127_start), .goal(_add_map_x_127_goal), .now(_add_map_x_127_now));
add_map add_map_x_126 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_126_add_exe), .data_out(_add_map_x_126_data_out), .data_out_index(_add_map_x_126_data_out_index), .data_near(_add_map_x_126_data_near), .wall_t_out(_add_map_x_126_wall_t_out), .data_org(_add_map_x_126_data_org), .data_org_near(_add_map_x_126_data_org_near), .s_g(_add_map_x_126_s_g), .s_g_near(_add_map_x_126_s_g_near), .moto_org_near(_add_map_x_126_moto_org_near), .moto_org_near1(_add_map_x_126_moto_org_near1), .moto_org_near2(_add_map_x_126_moto_org_near2), .moto_org_near3(_add_map_x_126_moto_org_near3), .moto_org(_add_map_x_126_moto_org), .sg_up(_add_map_x_126_sg_up), .sg_down(_add_map_x_126_sg_down), .sg_left(_add_map_x_126_sg_left), .sg_right(_add_map_x_126_sg_right), .wall_t_in(_add_map_x_126_wall_t_in), .moto(_add_map_x_126_moto), .up(_add_map_x_126_up), .right(_add_map_x_126_right), .down(_add_map_x_126_down), .left(_add_map_x_126_left), .start(_add_map_x_126_start), .goal(_add_map_x_126_goal), .now(_add_map_x_126_now));
add_map add_map_x_125 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_125_add_exe), .data_out(_add_map_x_125_data_out), .data_out_index(_add_map_x_125_data_out_index), .data_near(_add_map_x_125_data_near), .wall_t_out(_add_map_x_125_wall_t_out), .data_org(_add_map_x_125_data_org), .data_org_near(_add_map_x_125_data_org_near), .s_g(_add_map_x_125_s_g), .s_g_near(_add_map_x_125_s_g_near), .moto_org_near(_add_map_x_125_moto_org_near), .moto_org_near1(_add_map_x_125_moto_org_near1), .moto_org_near2(_add_map_x_125_moto_org_near2), .moto_org_near3(_add_map_x_125_moto_org_near3), .moto_org(_add_map_x_125_moto_org), .sg_up(_add_map_x_125_sg_up), .sg_down(_add_map_x_125_sg_down), .sg_left(_add_map_x_125_sg_left), .sg_right(_add_map_x_125_sg_right), .wall_t_in(_add_map_x_125_wall_t_in), .moto(_add_map_x_125_moto), .up(_add_map_x_125_up), .right(_add_map_x_125_right), .down(_add_map_x_125_down), .left(_add_map_x_125_left), .start(_add_map_x_125_start), .goal(_add_map_x_125_goal), .now(_add_map_x_125_now));
add_map add_map_x_124 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_124_add_exe), .data_out(_add_map_x_124_data_out), .data_out_index(_add_map_x_124_data_out_index), .data_near(_add_map_x_124_data_near), .wall_t_out(_add_map_x_124_wall_t_out), .data_org(_add_map_x_124_data_org), .data_org_near(_add_map_x_124_data_org_near), .s_g(_add_map_x_124_s_g), .s_g_near(_add_map_x_124_s_g_near), .moto_org_near(_add_map_x_124_moto_org_near), .moto_org_near1(_add_map_x_124_moto_org_near1), .moto_org_near2(_add_map_x_124_moto_org_near2), .moto_org_near3(_add_map_x_124_moto_org_near3), .moto_org(_add_map_x_124_moto_org), .sg_up(_add_map_x_124_sg_up), .sg_down(_add_map_x_124_sg_down), .sg_left(_add_map_x_124_sg_left), .sg_right(_add_map_x_124_sg_right), .wall_t_in(_add_map_x_124_wall_t_in), .moto(_add_map_x_124_moto), .up(_add_map_x_124_up), .right(_add_map_x_124_right), .down(_add_map_x_124_down), .left(_add_map_x_124_left), .start(_add_map_x_124_start), .goal(_add_map_x_124_goal), .now(_add_map_x_124_now));
add_map add_map_x_123 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_123_add_exe), .data_out(_add_map_x_123_data_out), .data_out_index(_add_map_x_123_data_out_index), .data_near(_add_map_x_123_data_near), .wall_t_out(_add_map_x_123_wall_t_out), .data_org(_add_map_x_123_data_org), .data_org_near(_add_map_x_123_data_org_near), .s_g(_add_map_x_123_s_g), .s_g_near(_add_map_x_123_s_g_near), .moto_org_near(_add_map_x_123_moto_org_near), .moto_org_near1(_add_map_x_123_moto_org_near1), .moto_org_near2(_add_map_x_123_moto_org_near2), .moto_org_near3(_add_map_x_123_moto_org_near3), .moto_org(_add_map_x_123_moto_org), .sg_up(_add_map_x_123_sg_up), .sg_down(_add_map_x_123_sg_down), .sg_left(_add_map_x_123_sg_left), .sg_right(_add_map_x_123_sg_right), .wall_t_in(_add_map_x_123_wall_t_in), .moto(_add_map_x_123_moto), .up(_add_map_x_123_up), .right(_add_map_x_123_right), .down(_add_map_x_123_down), .left(_add_map_x_123_left), .start(_add_map_x_123_start), .goal(_add_map_x_123_goal), .now(_add_map_x_123_now));
add_map add_map_x_122 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_122_add_exe), .data_out(_add_map_x_122_data_out), .data_out_index(_add_map_x_122_data_out_index), .data_near(_add_map_x_122_data_near), .wall_t_out(_add_map_x_122_wall_t_out), .data_org(_add_map_x_122_data_org), .data_org_near(_add_map_x_122_data_org_near), .s_g(_add_map_x_122_s_g), .s_g_near(_add_map_x_122_s_g_near), .moto_org_near(_add_map_x_122_moto_org_near), .moto_org_near1(_add_map_x_122_moto_org_near1), .moto_org_near2(_add_map_x_122_moto_org_near2), .moto_org_near3(_add_map_x_122_moto_org_near3), .moto_org(_add_map_x_122_moto_org), .sg_up(_add_map_x_122_sg_up), .sg_down(_add_map_x_122_sg_down), .sg_left(_add_map_x_122_sg_left), .sg_right(_add_map_x_122_sg_right), .wall_t_in(_add_map_x_122_wall_t_in), .moto(_add_map_x_122_moto), .up(_add_map_x_122_up), .right(_add_map_x_122_right), .down(_add_map_x_122_down), .left(_add_map_x_122_left), .start(_add_map_x_122_start), .goal(_add_map_x_122_goal), .now(_add_map_x_122_now));
add_map add_map_x_121 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_121_add_exe), .data_out(_add_map_x_121_data_out), .data_out_index(_add_map_x_121_data_out_index), .data_near(_add_map_x_121_data_near), .wall_t_out(_add_map_x_121_wall_t_out), .data_org(_add_map_x_121_data_org), .data_org_near(_add_map_x_121_data_org_near), .s_g(_add_map_x_121_s_g), .s_g_near(_add_map_x_121_s_g_near), .moto_org_near(_add_map_x_121_moto_org_near), .moto_org_near1(_add_map_x_121_moto_org_near1), .moto_org_near2(_add_map_x_121_moto_org_near2), .moto_org_near3(_add_map_x_121_moto_org_near3), .moto_org(_add_map_x_121_moto_org), .sg_up(_add_map_x_121_sg_up), .sg_down(_add_map_x_121_sg_down), .sg_left(_add_map_x_121_sg_left), .sg_right(_add_map_x_121_sg_right), .wall_t_in(_add_map_x_121_wall_t_in), .moto(_add_map_x_121_moto), .up(_add_map_x_121_up), .right(_add_map_x_121_right), .down(_add_map_x_121_down), .left(_add_map_x_121_left), .start(_add_map_x_121_start), .goal(_add_map_x_121_goal), .now(_add_map_x_121_now));
add_map add_map_x_120 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_120_add_exe), .data_out(_add_map_x_120_data_out), .data_out_index(_add_map_x_120_data_out_index), .data_near(_add_map_x_120_data_near), .wall_t_out(_add_map_x_120_wall_t_out), .data_org(_add_map_x_120_data_org), .data_org_near(_add_map_x_120_data_org_near), .s_g(_add_map_x_120_s_g), .s_g_near(_add_map_x_120_s_g_near), .moto_org_near(_add_map_x_120_moto_org_near), .moto_org_near1(_add_map_x_120_moto_org_near1), .moto_org_near2(_add_map_x_120_moto_org_near2), .moto_org_near3(_add_map_x_120_moto_org_near3), .moto_org(_add_map_x_120_moto_org), .sg_up(_add_map_x_120_sg_up), .sg_down(_add_map_x_120_sg_down), .sg_left(_add_map_x_120_sg_left), .sg_right(_add_map_x_120_sg_right), .wall_t_in(_add_map_x_120_wall_t_in), .moto(_add_map_x_120_moto), .up(_add_map_x_120_up), .right(_add_map_x_120_right), .down(_add_map_x_120_down), .left(_add_map_x_120_left), .start(_add_map_x_120_start), .goal(_add_map_x_120_goal), .now(_add_map_x_120_now));
add_map add_map_x_119 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_119_add_exe), .data_out(_add_map_x_119_data_out), .data_out_index(_add_map_x_119_data_out_index), .data_near(_add_map_x_119_data_near), .wall_t_out(_add_map_x_119_wall_t_out), .data_org(_add_map_x_119_data_org), .data_org_near(_add_map_x_119_data_org_near), .s_g(_add_map_x_119_s_g), .s_g_near(_add_map_x_119_s_g_near), .moto_org_near(_add_map_x_119_moto_org_near), .moto_org_near1(_add_map_x_119_moto_org_near1), .moto_org_near2(_add_map_x_119_moto_org_near2), .moto_org_near3(_add_map_x_119_moto_org_near3), .moto_org(_add_map_x_119_moto_org), .sg_up(_add_map_x_119_sg_up), .sg_down(_add_map_x_119_sg_down), .sg_left(_add_map_x_119_sg_left), .sg_right(_add_map_x_119_sg_right), .wall_t_in(_add_map_x_119_wall_t_in), .moto(_add_map_x_119_moto), .up(_add_map_x_119_up), .right(_add_map_x_119_right), .down(_add_map_x_119_down), .left(_add_map_x_119_left), .start(_add_map_x_119_start), .goal(_add_map_x_119_goal), .now(_add_map_x_119_now));
add_map add_map_x_118 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_118_add_exe), .data_out(_add_map_x_118_data_out), .data_out_index(_add_map_x_118_data_out_index), .data_near(_add_map_x_118_data_near), .wall_t_out(_add_map_x_118_wall_t_out), .data_org(_add_map_x_118_data_org), .data_org_near(_add_map_x_118_data_org_near), .s_g(_add_map_x_118_s_g), .s_g_near(_add_map_x_118_s_g_near), .moto_org_near(_add_map_x_118_moto_org_near), .moto_org_near1(_add_map_x_118_moto_org_near1), .moto_org_near2(_add_map_x_118_moto_org_near2), .moto_org_near3(_add_map_x_118_moto_org_near3), .moto_org(_add_map_x_118_moto_org), .sg_up(_add_map_x_118_sg_up), .sg_down(_add_map_x_118_sg_down), .sg_left(_add_map_x_118_sg_left), .sg_right(_add_map_x_118_sg_right), .wall_t_in(_add_map_x_118_wall_t_in), .moto(_add_map_x_118_moto), .up(_add_map_x_118_up), .right(_add_map_x_118_right), .down(_add_map_x_118_down), .left(_add_map_x_118_left), .start(_add_map_x_118_start), .goal(_add_map_x_118_goal), .now(_add_map_x_118_now));
add_map add_map_x_117 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_117_add_exe), .data_out(_add_map_x_117_data_out), .data_out_index(_add_map_x_117_data_out_index), .data_near(_add_map_x_117_data_near), .wall_t_out(_add_map_x_117_wall_t_out), .data_org(_add_map_x_117_data_org), .data_org_near(_add_map_x_117_data_org_near), .s_g(_add_map_x_117_s_g), .s_g_near(_add_map_x_117_s_g_near), .moto_org_near(_add_map_x_117_moto_org_near), .moto_org_near1(_add_map_x_117_moto_org_near1), .moto_org_near2(_add_map_x_117_moto_org_near2), .moto_org_near3(_add_map_x_117_moto_org_near3), .moto_org(_add_map_x_117_moto_org), .sg_up(_add_map_x_117_sg_up), .sg_down(_add_map_x_117_sg_down), .sg_left(_add_map_x_117_sg_left), .sg_right(_add_map_x_117_sg_right), .wall_t_in(_add_map_x_117_wall_t_in), .moto(_add_map_x_117_moto), .up(_add_map_x_117_up), .right(_add_map_x_117_right), .down(_add_map_x_117_down), .left(_add_map_x_117_left), .start(_add_map_x_117_start), .goal(_add_map_x_117_goal), .now(_add_map_x_117_now));
add_map add_map_x_116 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_116_add_exe), .data_out(_add_map_x_116_data_out), .data_out_index(_add_map_x_116_data_out_index), .data_near(_add_map_x_116_data_near), .wall_t_out(_add_map_x_116_wall_t_out), .data_org(_add_map_x_116_data_org), .data_org_near(_add_map_x_116_data_org_near), .s_g(_add_map_x_116_s_g), .s_g_near(_add_map_x_116_s_g_near), .moto_org_near(_add_map_x_116_moto_org_near), .moto_org_near1(_add_map_x_116_moto_org_near1), .moto_org_near2(_add_map_x_116_moto_org_near2), .moto_org_near3(_add_map_x_116_moto_org_near3), .moto_org(_add_map_x_116_moto_org), .sg_up(_add_map_x_116_sg_up), .sg_down(_add_map_x_116_sg_down), .sg_left(_add_map_x_116_sg_left), .sg_right(_add_map_x_116_sg_right), .wall_t_in(_add_map_x_116_wall_t_in), .moto(_add_map_x_116_moto), .up(_add_map_x_116_up), .right(_add_map_x_116_right), .down(_add_map_x_116_down), .left(_add_map_x_116_left), .start(_add_map_x_116_start), .goal(_add_map_x_116_goal), .now(_add_map_x_116_now));
add_map add_map_x_115 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_115_add_exe), .data_out(_add_map_x_115_data_out), .data_out_index(_add_map_x_115_data_out_index), .data_near(_add_map_x_115_data_near), .wall_t_out(_add_map_x_115_wall_t_out), .data_org(_add_map_x_115_data_org), .data_org_near(_add_map_x_115_data_org_near), .s_g(_add_map_x_115_s_g), .s_g_near(_add_map_x_115_s_g_near), .moto_org_near(_add_map_x_115_moto_org_near), .moto_org_near1(_add_map_x_115_moto_org_near1), .moto_org_near2(_add_map_x_115_moto_org_near2), .moto_org_near3(_add_map_x_115_moto_org_near3), .moto_org(_add_map_x_115_moto_org), .sg_up(_add_map_x_115_sg_up), .sg_down(_add_map_x_115_sg_down), .sg_left(_add_map_x_115_sg_left), .sg_right(_add_map_x_115_sg_right), .wall_t_in(_add_map_x_115_wall_t_in), .moto(_add_map_x_115_moto), .up(_add_map_x_115_up), .right(_add_map_x_115_right), .down(_add_map_x_115_down), .left(_add_map_x_115_left), .start(_add_map_x_115_start), .goal(_add_map_x_115_goal), .now(_add_map_x_115_now));
add_map add_map_x_114 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_114_add_exe), .data_out(_add_map_x_114_data_out), .data_out_index(_add_map_x_114_data_out_index), .data_near(_add_map_x_114_data_near), .wall_t_out(_add_map_x_114_wall_t_out), .data_org(_add_map_x_114_data_org), .data_org_near(_add_map_x_114_data_org_near), .s_g(_add_map_x_114_s_g), .s_g_near(_add_map_x_114_s_g_near), .moto_org_near(_add_map_x_114_moto_org_near), .moto_org_near1(_add_map_x_114_moto_org_near1), .moto_org_near2(_add_map_x_114_moto_org_near2), .moto_org_near3(_add_map_x_114_moto_org_near3), .moto_org(_add_map_x_114_moto_org), .sg_up(_add_map_x_114_sg_up), .sg_down(_add_map_x_114_sg_down), .sg_left(_add_map_x_114_sg_left), .sg_right(_add_map_x_114_sg_right), .wall_t_in(_add_map_x_114_wall_t_in), .moto(_add_map_x_114_moto), .up(_add_map_x_114_up), .right(_add_map_x_114_right), .down(_add_map_x_114_down), .left(_add_map_x_114_left), .start(_add_map_x_114_start), .goal(_add_map_x_114_goal), .now(_add_map_x_114_now));
add_map add_map_x_113 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_113_add_exe), .data_out(_add_map_x_113_data_out), .data_out_index(_add_map_x_113_data_out_index), .data_near(_add_map_x_113_data_near), .wall_t_out(_add_map_x_113_wall_t_out), .data_org(_add_map_x_113_data_org), .data_org_near(_add_map_x_113_data_org_near), .s_g(_add_map_x_113_s_g), .s_g_near(_add_map_x_113_s_g_near), .moto_org_near(_add_map_x_113_moto_org_near), .moto_org_near1(_add_map_x_113_moto_org_near1), .moto_org_near2(_add_map_x_113_moto_org_near2), .moto_org_near3(_add_map_x_113_moto_org_near3), .moto_org(_add_map_x_113_moto_org), .sg_up(_add_map_x_113_sg_up), .sg_down(_add_map_x_113_sg_down), .sg_left(_add_map_x_113_sg_left), .sg_right(_add_map_x_113_sg_right), .wall_t_in(_add_map_x_113_wall_t_in), .moto(_add_map_x_113_moto), .up(_add_map_x_113_up), .right(_add_map_x_113_right), .down(_add_map_x_113_down), .left(_add_map_x_113_left), .start(_add_map_x_113_start), .goal(_add_map_x_113_goal), .now(_add_map_x_113_now));
add_map add_map_x_112 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_112_add_exe), .data_out(_add_map_x_112_data_out), .data_out_index(_add_map_x_112_data_out_index), .data_near(_add_map_x_112_data_near), .wall_t_out(_add_map_x_112_wall_t_out), .data_org(_add_map_x_112_data_org), .data_org_near(_add_map_x_112_data_org_near), .s_g(_add_map_x_112_s_g), .s_g_near(_add_map_x_112_s_g_near), .moto_org_near(_add_map_x_112_moto_org_near), .moto_org_near1(_add_map_x_112_moto_org_near1), .moto_org_near2(_add_map_x_112_moto_org_near2), .moto_org_near3(_add_map_x_112_moto_org_near3), .moto_org(_add_map_x_112_moto_org), .sg_up(_add_map_x_112_sg_up), .sg_down(_add_map_x_112_sg_down), .sg_left(_add_map_x_112_sg_left), .sg_right(_add_map_x_112_sg_right), .wall_t_in(_add_map_x_112_wall_t_in), .moto(_add_map_x_112_moto), .up(_add_map_x_112_up), .right(_add_map_x_112_right), .down(_add_map_x_112_down), .left(_add_map_x_112_left), .start(_add_map_x_112_start), .goal(_add_map_x_112_goal), .now(_add_map_x_112_now));
add_map add_map_x_111 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_111_add_exe), .data_out(_add_map_x_111_data_out), .data_out_index(_add_map_x_111_data_out_index), .data_near(_add_map_x_111_data_near), .wall_t_out(_add_map_x_111_wall_t_out), .data_org(_add_map_x_111_data_org), .data_org_near(_add_map_x_111_data_org_near), .s_g(_add_map_x_111_s_g), .s_g_near(_add_map_x_111_s_g_near), .moto_org_near(_add_map_x_111_moto_org_near), .moto_org_near1(_add_map_x_111_moto_org_near1), .moto_org_near2(_add_map_x_111_moto_org_near2), .moto_org_near3(_add_map_x_111_moto_org_near3), .moto_org(_add_map_x_111_moto_org), .sg_up(_add_map_x_111_sg_up), .sg_down(_add_map_x_111_sg_down), .sg_left(_add_map_x_111_sg_left), .sg_right(_add_map_x_111_sg_right), .wall_t_in(_add_map_x_111_wall_t_in), .moto(_add_map_x_111_moto), .up(_add_map_x_111_up), .right(_add_map_x_111_right), .down(_add_map_x_111_down), .left(_add_map_x_111_left), .start(_add_map_x_111_start), .goal(_add_map_x_111_goal), .now(_add_map_x_111_now));
add_map add_map_x_110 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_110_add_exe), .data_out(_add_map_x_110_data_out), .data_out_index(_add_map_x_110_data_out_index), .data_near(_add_map_x_110_data_near), .wall_t_out(_add_map_x_110_wall_t_out), .data_org(_add_map_x_110_data_org), .data_org_near(_add_map_x_110_data_org_near), .s_g(_add_map_x_110_s_g), .s_g_near(_add_map_x_110_s_g_near), .moto_org_near(_add_map_x_110_moto_org_near), .moto_org_near1(_add_map_x_110_moto_org_near1), .moto_org_near2(_add_map_x_110_moto_org_near2), .moto_org_near3(_add_map_x_110_moto_org_near3), .moto_org(_add_map_x_110_moto_org), .sg_up(_add_map_x_110_sg_up), .sg_down(_add_map_x_110_sg_down), .sg_left(_add_map_x_110_sg_left), .sg_right(_add_map_x_110_sg_right), .wall_t_in(_add_map_x_110_wall_t_in), .moto(_add_map_x_110_moto), .up(_add_map_x_110_up), .right(_add_map_x_110_right), .down(_add_map_x_110_down), .left(_add_map_x_110_left), .start(_add_map_x_110_start), .goal(_add_map_x_110_goal), .now(_add_map_x_110_now));
add_map add_map_x_109 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_109_add_exe), .data_out(_add_map_x_109_data_out), .data_out_index(_add_map_x_109_data_out_index), .data_near(_add_map_x_109_data_near), .wall_t_out(_add_map_x_109_wall_t_out), .data_org(_add_map_x_109_data_org), .data_org_near(_add_map_x_109_data_org_near), .s_g(_add_map_x_109_s_g), .s_g_near(_add_map_x_109_s_g_near), .moto_org_near(_add_map_x_109_moto_org_near), .moto_org_near1(_add_map_x_109_moto_org_near1), .moto_org_near2(_add_map_x_109_moto_org_near2), .moto_org_near3(_add_map_x_109_moto_org_near3), .moto_org(_add_map_x_109_moto_org), .sg_up(_add_map_x_109_sg_up), .sg_down(_add_map_x_109_sg_down), .sg_left(_add_map_x_109_sg_left), .sg_right(_add_map_x_109_sg_right), .wall_t_in(_add_map_x_109_wall_t_in), .moto(_add_map_x_109_moto), .up(_add_map_x_109_up), .right(_add_map_x_109_right), .down(_add_map_x_109_down), .left(_add_map_x_109_left), .start(_add_map_x_109_start), .goal(_add_map_x_109_goal), .now(_add_map_x_109_now));
add_map add_map_x_108 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_108_add_exe), .data_out(_add_map_x_108_data_out), .data_out_index(_add_map_x_108_data_out_index), .data_near(_add_map_x_108_data_near), .wall_t_out(_add_map_x_108_wall_t_out), .data_org(_add_map_x_108_data_org), .data_org_near(_add_map_x_108_data_org_near), .s_g(_add_map_x_108_s_g), .s_g_near(_add_map_x_108_s_g_near), .moto_org_near(_add_map_x_108_moto_org_near), .moto_org_near1(_add_map_x_108_moto_org_near1), .moto_org_near2(_add_map_x_108_moto_org_near2), .moto_org_near3(_add_map_x_108_moto_org_near3), .moto_org(_add_map_x_108_moto_org), .sg_up(_add_map_x_108_sg_up), .sg_down(_add_map_x_108_sg_down), .sg_left(_add_map_x_108_sg_left), .sg_right(_add_map_x_108_sg_right), .wall_t_in(_add_map_x_108_wall_t_in), .moto(_add_map_x_108_moto), .up(_add_map_x_108_up), .right(_add_map_x_108_right), .down(_add_map_x_108_down), .left(_add_map_x_108_left), .start(_add_map_x_108_start), .goal(_add_map_x_108_goal), .now(_add_map_x_108_now));
add_map add_map_x_107 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_107_add_exe), .data_out(_add_map_x_107_data_out), .data_out_index(_add_map_x_107_data_out_index), .data_near(_add_map_x_107_data_near), .wall_t_out(_add_map_x_107_wall_t_out), .data_org(_add_map_x_107_data_org), .data_org_near(_add_map_x_107_data_org_near), .s_g(_add_map_x_107_s_g), .s_g_near(_add_map_x_107_s_g_near), .moto_org_near(_add_map_x_107_moto_org_near), .moto_org_near1(_add_map_x_107_moto_org_near1), .moto_org_near2(_add_map_x_107_moto_org_near2), .moto_org_near3(_add_map_x_107_moto_org_near3), .moto_org(_add_map_x_107_moto_org), .sg_up(_add_map_x_107_sg_up), .sg_down(_add_map_x_107_sg_down), .sg_left(_add_map_x_107_sg_left), .sg_right(_add_map_x_107_sg_right), .wall_t_in(_add_map_x_107_wall_t_in), .moto(_add_map_x_107_moto), .up(_add_map_x_107_up), .right(_add_map_x_107_right), .down(_add_map_x_107_down), .left(_add_map_x_107_left), .start(_add_map_x_107_start), .goal(_add_map_x_107_goal), .now(_add_map_x_107_now));
add_map add_map_x_106 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_106_add_exe), .data_out(_add_map_x_106_data_out), .data_out_index(_add_map_x_106_data_out_index), .data_near(_add_map_x_106_data_near), .wall_t_out(_add_map_x_106_wall_t_out), .data_org(_add_map_x_106_data_org), .data_org_near(_add_map_x_106_data_org_near), .s_g(_add_map_x_106_s_g), .s_g_near(_add_map_x_106_s_g_near), .moto_org_near(_add_map_x_106_moto_org_near), .moto_org_near1(_add_map_x_106_moto_org_near1), .moto_org_near2(_add_map_x_106_moto_org_near2), .moto_org_near3(_add_map_x_106_moto_org_near3), .moto_org(_add_map_x_106_moto_org), .sg_up(_add_map_x_106_sg_up), .sg_down(_add_map_x_106_sg_down), .sg_left(_add_map_x_106_sg_left), .sg_right(_add_map_x_106_sg_right), .wall_t_in(_add_map_x_106_wall_t_in), .moto(_add_map_x_106_moto), .up(_add_map_x_106_up), .right(_add_map_x_106_right), .down(_add_map_x_106_down), .left(_add_map_x_106_left), .start(_add_map_x_106_start), .goal(_add_map_x_106_goal), .now(_add_map_x_106_now));
add_map add_map_x_105 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_105_add_exe), .data_out(_add_map_x_105_data_out), .data_out_index(_add_map_x_105_data_out_index), .data_near(_add_map_x_105_data_near), .wall_t_out(_add_map_x_105_wall_t_out), .data_org(_add_map_x_105_data_org), .data_org_near(_add_map_x_105_data_org_near), .s_g(_add_map_x_105_s_g), .s_g_near(_add_map_x_105_s_g_near), .moto_org_near(_add_map_x_105_moto_org_near), .moto_org_near1(_add_map_x_105_moto_org_near1), .moto_org_near2(_add_map_x_105_moto_org_near2), .moto_org_near3(_add_map_x_105_moto_org_near3), .moto_org(_add_map_x_105_moto_org), .sg_up(_add_map_x_105_sg_up), .sg_down(_add_map_x_105_sg_down), .sg_left(_add_map_x_105_sg_left), .sg_right(_add_map_x_105_sg_right), .wall_t_in(_add_map_x_105_wall_t_in), .moto(_add_map_x_105_moto), .up(_add_map_x_105_up), .right(_add_map_x_105_right), .down(_add_map_x_105_down), .left(_add_map_x_105_left), .start(_add_map_x_105_start), .goal(_add_map_x_105_goal), .now(_add_map_x_105_now));
add_map add_map_x_104 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_104_add_exe), .data_out(_add_map_x_104_data_out), .data_out_index(_add_map_x_104_data_out_index), .data_near(_add_map_x_104_data_near), .wall_t_out(_add_map_x_104_wall_t_out), .data_org(_add_map_x_104_data_org), .data_org_near(_add_map_x_104_data_org_near), .s_g(_add_map_x_104_s_g), .s_g_near(_add_map_x_104_s_g_near), .moto_org_near(_add_map_x_104_moto_org_near), .moto_org_near1(_add_map_x_104_moto_org_near1), .moto_org_near2(_add_map_x_104_moto_org_near2), .moto_org_near3(_add_map_x_104_moto_org_near3), .moto_org(_add_map_x_104_moto_org), .sg_up(_add_map_x_104_sg_up), .sg_down(_add_map_x_104_sg_down), .sg_left(_add_map_x_104_sg_left), .sg_right(_add_map_x_104_sg_right), .wall_t_in(_add_map_x_104_wall_t_in), .moto(_add_map_x_104_moto), .up(_add_map_x_104_up), .right(_add_map_x_104_right), .down(_add_map_x_104_down), .left(_add_map_x_104_left), .start(_add_map_x_104_start), .goal(_add_map_x_104_goal), .now(_add_map_x_104_now));
add_map add_map_x_103 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_103_add_exe), .data_out(_add_map_x_103_data_out), .data_out_index(_add_map_x_103_data_out_index), .data_near(_add_map_x_103_data_near), .wall_t_out(_add_map_x_103_wall_t_out), .data_org(_add_map_x_103_data_org), .data_org_near(_add_map_x_103_data_org_near), .s_g(_add_map_x_103_s_g), .s_g_near(_add_map_x_103_s_g_near), .moto_org_near(_add_map_x_103_moto_org_near), .moto_org_near1(_add_map_x_103_moto_org_near1), .moto_org_near2(_add_map_x_103_moto_org_near2), .moto_org_near3(_add_map_x_103_moto_org_near3), .moto_org(_add_map_x_103_moto_org), .sg_up(_add_map_x_103_sg_up), .sg_down(_add_map_x_103_sg_down), .sg_left(_add_map_x_103_sg_left), .sg_right(_add_map_x_103_sg_right), .wall_t_in(_add_map_x_103_wall_t_in), .moto(_add_map_x_103_moto), .up(_add_map_x_103_up), .right(_add_map_x_103_right), .down(_add_map_x_103_down), .left(_add_map_x_103_left), .start(_add_map_x_103_start), .goal(_add_map_x_103_goal), .now(_add_map_x_103_now));
add_map add_map_x_102 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_102_add_exe), .data_out(_add_map_x_102_data_out), .data_out_index(_add_map_x_102_data_out_index), .data_near(_add_map_x_102_data_near), .wall_t_out(_add_map_x_102_wall_t_out), .data_org(_add_map_x_102_data_org), .data_org_near(_add_map_x_102_data_org_near), .s_g(_add_map_x_102_s_g), .s_g_near(_add_map_x_102_s_g_near), .moto_org_near(_add_map_x_102_moto_org_near), .moto_org_near1(_add_map_x_102_moto_org_near1), .moto_org_near2(_add_map_x_102_moto_org_near2), .moto_org_near3(_add_map_x_102_moto_org_near3), .moto_org(_add_map_x_102_moto_org), .sg_up(_add_map_x_102_sg_up), .sg_down(_add_map_x_102_sg_down), .sg_left(_add_map_x_102_sg_left), .sg_right(_add_map_x_102_sg_right), .wall_t_in(_add_map_x_102_wall_t_in), .moto(_add_map_x_102_moto), .up(_add_map_x_102_up), .right(_add_map_x_102_right), .down(_add_map_x_102_down), .left(_add_map_x_102_left), .start(_add_map_x_102_start), .goal(_add_map_x_102_goal), .now(_add_map_x_102_now));
add_map add_map_x_101 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_101_add_exe), .data_out(_add_map_x_101_data_out), .data_out_index(_add_map_x_101_data_out_index), .data_near(_add_map_x_101_data_near), .wall_t_out(_add_map_x_101_wall_t_out), .data_org(_add_map_x_101_data_org), .data_org_near(_add_map_x_101_data_org_near), .s_g(_add_map_x_101_s_g), .s_g_near(_add_map_x_101_s_g_near), .moto_org_near(_add_map_x_101_moto_org_near), .moto_org_near1(_add_map_x_101_moto_org_near1), .moto_org_near2(_add_map_x_101_moto_org_near2), .moto_org_near3(_add_map_x_101_moto_org_near3), .moto_org(_add_map_x_101_moto_org), .sg_up(_add_map_x_101_sg_up), .sg_down(_add_map_x_101_sg_down), .sg_left(_add_map_x_101_sg_left), .sg_right(_add_map_x_101_sg_right), .wall_t_in(_add_map_x_101_wall_t_in), .moto(_add_map_x_101_moto), .up(_add_map_x_101_up), .right(_add_map_x_101_right), .down(_add_map_x_101_down), .left(_add_map_x_101_left), .start(_add_map_x_101_start), .goal(_add_map_x_101_goal), .now(_add_map_x_101_now));
add_map add_map_x_100 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_100_add_exe), .data_out(_add_map_x_100_data_out), .data_out_index(_add_map_x_100_data_out_index), .data_near(_add_map_x_100_data_near), .wall_t_out(_add_map_x_100_wall_t_out), .data_org(_add_map_x_100_data_org), .data_org_near(_add_map_x_100_data_org_near), .s_g(_add_map_x_100_s_g), .s_g_near(_add_map_x_100_s_g_near), .moto_org_near(_add_map_x_100_moto_org_near), .moto_org_near1(_add_map_x_100_moto_org_near1), .moto_org_near2(_add_map_x_100_moto_org_near2), .moto_org_near3(_add_map_x_100_moto_org_near3), .moto_org(_add_map_x_100_moto_org), .sg_up(_add_map_x_100_sg_up), .sg_down(_add_map_x_100_sg_down), .sg_left(_add_map_x_100_sg_left), .sg_right(_add_map_x_100_sg_right), .wall_t_in(_add_map_x_100_wall_t_in), .moto(_add_map_x_100_moto), .up(_add_map_x_100_up), .right(_add_map_x_100_right), .down(_add_map_x_100_down), .left(_add_map_x_100_left), .start(_add_map_x_100_start), .goal(_add_map_x_100_goal), .now(_add_map_x_100_now));
add_map add_map_x_99 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_99_add_exe), .data_out(_add_map_x_99_data_out), .data_out_index(_add_map_x_99_data_out_index), .data_near(_add_map_x_99_data_near), .wall_t_out(_add_map_x_99_wall_t_out), .data_org(_add_map_x_99_data_org), .data_org_near(_add_map_x_99_data_org_near), .s_g(_add_map_x_99_s_g), .s_g_near(_add_map_x_99_s_g_near), .moto_org_near(_add_map_x_99_moto_org_near), .moto_org_near1(_add_map_x_99_moto_org_near1), .moto_org_near2(_add_map_x_99_moto_org_near2), .moto_org_near3(_add_map_x_99_moto_org_near3), .moto_org(_add_map_x_99_moto_org), .sg_up(_add_map_x_99_sg_up), .sg_down(_add_map_x_99_sg_down), .sg_left(_add_map_x_99_sg_left), .sg_right(_add_map_x_99_sg_right), .wall_t_in(_add_map_x_99_wall_t_in), .moto(_add_map_x_99_moto), .up(_add_map_x_99_up), .right(_add_map_x_99_right), .down(_add_map_x_99_down), .left(_add_map_x_99_left), .start(_add_map_x_99_start), .goal(_add_map_x_99_goal), .now(_add_map_x_99_now));
add_map add_map_x_98 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_98_add_exe), .data_out(_add_map_x_98_data_out), .data_out_index(_add_map_x_98_data_out_index), .data_near(_add_map_x_98_data_near), .wall_t_out(_add_map_x_98_wall_t_out), .data_org(_add_map_x_98_data_org), .data_org_near(_add_map_x_98_data_org_near), .s_g(_add_map_x_98_s_g), .s_g_near(_add_map_x_98_s_g_near), .moto_org_near(_add_map_x_98_moto_org_near), .moto_org_near1(_add_map_x_98_moto_org_near1), .moto_org_near2(_add_map_x_98_moto_org_near2), .moto_org_near3(_add_map_x_98_moto_org_near3), .moto_org(_add_map_x_98_moto_org), .sg_up(_add_map_x_98_sg_up), .sg_down(_add_map_x_98_sg_down), .sg_left(_add_map_x_98_sg_left), .sg_right(_add_map_x_98_sg_right), .wall_t_in(_add_map_x_98_wall_t_in), .moto(_add_map_x_98_moto), .up(_add_map_x_98_up), .right(_add_map_x_98_right), .down(_add_map_x_98_down), .left(_add_map_x_98_left), .start(_add_map_x_98_start), .goal(_add_map_x_98_goal), .now(_add_map_x_98_now));
add_map add_map_x_97 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_97_add_exe), .data_out(_add_map_x_97_data_out), .data_out_index(_add_map_x_97_data_out_index), .data_near(_add_map_x_97_data_near), .wall_t_out(_add_map_x_97_wall_t_out), .data_org(_add_map_x_97_data_org), .data_org_near(_add_map_x_97_data_org_near), .s_g(_add_map_x_97_s_g), .s_g_near(_add_map_x_97_s_g_near), .moto_org_near(_add_map_x_97_moto_org_near), .moto_org_near1(_add_map_x_97_moto_org_near1), .moto_org_near2(_add_map_x_97_moto_org_near2), .moto_org_near3(_add_map_x_97_moto_org_near3), .moto_org(_add_map_x_97_moto_org), .sg_up(_add_map_x_97_sg_up), .sg_down(_add_map_x_97_sg_down), .sg_left(_add_map_x_97_sg_left), .sg_right(_add_map_x_97_sg_right), .wall_t_in(_add_map_x_97_wall_t_in), .moto(_add_map_x_97_moto), .up(_add_map_x_97_up), .right(_add_map_x_97_right), .down(_add_map_x_97_down), .left(_add_map_x_97_left), .start(_add_map_x_97_start), .goal(_add_map_x_97_goal), .now(_add_map_x_97_now));
add_map add_map_x_96 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_96_add_exe), .data_out(_add_map_x_96_data_out), .data_out_index(_add_map_x_96_data_out_index), .data_near(_add_map_x_96_data_near), .wall_t_out(_add_map_x_96_wall_t_out), .data_org(_add_map_x_96_data_org), .data_org_near(_add_map_x_96_data_org_near), .s_g(_add_map_x_96_s_g), .s_g_near(_add_map_x_96_s_g_near), .moto_org_near(_add_map_x_96_moto_org_near), .moto_org_near1(_add_map_x_96_moto_org_near1), .moto_org_near2(_add_map_x_96_moto_org_near2), .moto_org_near3(_add_map_x_96_moto_org_near3), .moto_org(_add_map_x_96_moto_org), .sg_up(_add_map_x_96_sg_up), .sg_down(_add_map_x_96_sg_down), .sg_left(_add_map_x_96_sg_left), .sg_right(_add_map_x_96_sg_right), .wall_t_in(_add_map_x_96_wall_t_in), .moto(_add_map_x_96_moto), .up(_add_map_x_96_up), .right(_add_map_x_96_right), .down(_add_map_x_96_down), .left(_add_map_x_96_left), .start(_add_map_x_96_start), .goal(_add_map_x_96_goal), .now(_add_map_x_96_now));
add_map add_map_x_95 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_95_add_exe), .data_out(_add_map_x_95_data_out), .data_out_index(_add_map_x_95_data_out_index), .data_near(_add_map_x_95_data_near), .wall_t_out(_add_map_x_95_wall_t_out), .data_org(_add_map_x_95_data_org), .data_org_near(_add_map_x_95_data_org_near), .s_g(_add_map_x_95_s_g), .s_g_near(_add_map_x_95_s_g_near), .moto_org_near(_add_map_x_95_moto_org_near), .moto_org_near1(_add_map_x_95_moto_org_near1), .moto_org_near2(_add_map_x_95_moto_org_near2), .moto_org_near3(_add_map_x_95_moto_org_near3), .moto_org(_add_map_x_95_moto_org), .sg_up(_add_map_x_95_sg_up), .sg_down(_add_map_x_95_sg_down), .sg_left(_add_map_x_95_sg_left), .sg_right(_add_map_x_95_sg_right), .wall_t_in(_add_map_x_95_wall_t_in), .moto(_add_map_x_95_moto), .up(_add_map_x_95_up), .right(_add_map_x_95_right), .down(_add_map_x_95_down), .left(_add_map_x_95_left), .start(_add_map_x_95_start), .goal(_add_map_x_95_goal), .now(_add_map_x_95_now));
add_map add_map_x_94 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_94_add_exe), .data_out(_add_map_x_94_data_out), .data_out_index(_add_map_x_94_data_out_index), .data_near(_add_map_x_94_data_near), .wall_t_out(_add_map_x_94_wall_t_out), .data_org(_add_map_x_94_data_org), .data_org_near(_add_map_x_94_data_org_near), .s_g(_add_map_x_94_s_g), .s_g_near(_add_map_x_94_s_g_near), .moto_org_near(_add_map_x_94_moto_org_near), .moto_org_near1(_add_map_x_94_moto_org_near1), .moto_org_near2(_add_map_x_94_moto_org_near2), .moto_org_near3(_add_map_x_94_moto_org_near3), .moto_org(_add_map_x_94_moto_org), .sg_up(_add_map_x_94_sg_up), .sg_down(_add_map_x_94_sg_down), .sg_left(_add_map_x_94_sg_left), .sg_right(_add_map_x_94_sg_right), .wall_t_in(_add_map_x_94_wall_t_in), .moto(_add_map_x_94_moto), .up(_add_map_x_94_up), .right(_add_map_x_94_right), .down(_add_map_x_94_down), .left(_add_map_x_94_left), .start(_add_map_x_94_start), .goal(_add_map_x_94_goal), .now(_add_map_x_94_now));
add_map add_map_x_93 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_93_add_exe), .data_out(_add_map_x_93_data_out), .data_out_index(_add_map_x_93_data_out_index), .data_near(_add_map_x_93_data_near), .wall_t_out(_add_map_x_93_wall_t_out), .data_org(_add_map_x_93_data_org), .data_org_near(_add_map_x_93_data_org_near), .s_g(_add_map_x_93_s_g), .s_g_near(_add_map_x_93_s_g_near), .moto_org_near(_add_map_x_93_moto_org_near), .moto_org_near1(_add_map_x_93_moto_org_near1), .moto_org_near2(_add_map_x_93_moto_org_near2), .moto_org_near3(_add_map_x_93_moto_org_near3), .moto_org(_add_map_x_93_moto_org), .sg_up(_add_map_x_93_sg_up), .sg_down(_add_map_x_93_sg_down), .sg_left(_add_map_x_93_sg_left), .sg_right(_add_map_x_93_sg_right), .wall_t_in(_add_map_x_93_wall_t_in), .moto(_add_map_x_93_moto), .up(_add_map_x_93_up), .right(_add_map_x_93_right), .down(_add_map_x_93_down), .left(_add_map_x_93_left), .start(_add_map_x_93_start), .goal(_add_map_x_93_goal), .now(_add_map_x_93_now));
add_map add_map_x_92 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_92_add_exe), .data_out(_add_map_x_92_data_out), .data_out_index(_add_map_x_92_data_out_index), .data_near(_add_map_x_92_data_near), .wall_t_out(_add_map_x_92_wall_t_out), .data_org(_add_map_x_92_data_org), .data_org_near(_add_map_x_92_data_org_near), .s_g(_add_map_x_92_s_g), .s_g_near(_add_map_x_92_s_g_near), .moto_org_near(_add_map_x_92_moto_org_near), .moto_org_near1(_add_map_x_92_moto_org_near1), .moto_org_near2(_add_map_x_92_moto_org_near2), .moto_org_near3(_add_map_x_92_moto_org_near3), .moto_org(_add_map_x_92_moto_org), .sg_up(_add_map_x_92_sg_up), .sg_down(_add_map_x_92_sg_down), .sg_left(_add_map_x_92_sg_left), .sg_right(_add_map_x_92_sg_right), .wall_t_in(_add_map_x_92_wall_t_in), .moto(_add_map_x_92_moto), .up(_add_map_x_92_up), .right(_add_map_x_92_right), .down(_add_map_x_92_down), .left(_add_map_x_92_left), .start(_add_map_x_92_start), .goal(_add_map_x_92_goal), .now(_add_map_x_92_now));
add_map add_map_x_91 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_91_add_exe), .data_out(_add_map_x_91_data_out), .data_out_index(_add_map_x_91_data_out_index), .data_near(_add_map_x_91_data_near), .wall_t_out(_add_map_x_91_wall_t_out), .data_org(_add_map_x_91_data_org), .data_org_near(_add_map_x_91_data_org_near), .s_g(_add_map_x_91_s_g), .s_g_near(_add_map_x_91_s_g_near), .moto_org_near(_add_map_x_91_moto_org_near), .moto_org_near1(_add_map_x_91_moto_org_near1), .moto_org_near2(_add_map_x_91_moto_org_near2), .moto_org_near3(_add_map_x_91_moto_org_near3), .moto_org(_add_map_x_91_moto_org), .sg_up(_add_map_x_91_sg_up), .sg_down(_add_map_x_91_sg_down), .sg_left(_add_map_x_91_sg_left), .sg_right(_add_map_x_91_sg_right), .wall_t_in(_add_map_x_91_wall_t_in), .moto(_add_map_x_91_moto), .up(_add_map_x_91_up), .right(_add_map_x_91_right), .down(_add_map_x_91_down), .left(_add_map_x_91_left), .start(_add_map_x_91_start), .goal(_add_map_x_91_goal), .now(_add_map_x_91_now));
add_map add_map_x_90 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_90_add_exe), .data_out(_add_map_x_90_data_out), .data_out_index(_add_map_x_90_data_out_index), .data_near(_add_map_x_90_data_near), .wall_t_out(_add_map_x_90_wall_t_out), .data_org(_add_map_x_90_data_org), .data_org_near(_add_map_x_90_data_org_near), .s_g(_add_map_x_90_s_g), .s_g_near(_add_map_x_90_s_g_near), .moto_org_near(_add_map_x_90_moto_org_near), .moto_org_near1(_add_map_x_90_moto_org_near1), .moto_org_near2(_add_map_x_90_moto_org_near2), .moto_org_near3(_add_map_x_90_moto_org_near3), .moto_org(_add_map_x_90_moto_org), .sg_up(_add_map_x_90_sg_up), .sg_down(_add_map_x_90_sg_down), .sg_left(_add_map_x_90_sg_left), .sg_right(_add_map_x_90_sg_right), .wall_t_in(_add_map_x_90_wall_t_in), .moto(_add_map_x_90_moto), .up(_add_map_x_90_up), .right(_add_map_x_90_right), .down(_add_map_x_90_down), .left(_add_map_x_90_left), .start(_add_map_x_90_start), .goal(_add_map_x_90_goal), .now(_add_map_x_90_now));
add_map add_map_x_89 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_89_add_exe), .data_out(_add_map_x_89_data_out), .data_out_index(_add_map_x_89_data_out_index), .data_near(_add_map_x_89_data_near), .wall_t_out(_add_map_x_89_wall_t_out), .data_org(_add_map_x_89_data_org), .data_org_near(_add_map_x_89_data_org_near), .s_g(_add_map_x_89_s_g), .s_g_near(_add_map_x_89_s_g_near), .moto_org_near(_add_map_x_89_moto_org_near), .moto_org_near1(_add_map_x_89_moto_org_near1), .moto_org_near2(_add_map_x_89_moto_org_near2), .moto_org_near3(_add_map_x_89_moto_org_near3), .moto_org(_add_map_x_89_moto_org), .sg_up(_add_map_x_89_sg_up), .sg_down(_add_map_x_89_sg_down), .sg_left(_add_map_x_89_sg_left), .sg_right(_add_map_x_89_sg_right), .wall_t_in(_add_map_x_89_wall_t_in), .moto(_add_map_x_89_moto), .up(_add_map_x_89_up), .right(_add_map_x_89_right), .down(_add_map_x_89_down), .left(_add_map_x_89_left), .start(_add_map_x_89_start), .goal(_add_map_x_89_goal), .now(_add_map_x_89_now));
add_map add_map_x_88 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_88_add_exe), .data_out(_add_map_x_88_data_out), .data_out_index(_add_map_x_88_data_out_index), .data_near(_add_map_x_88_data_near), .wall_t_out(_add_map_x_88_wall_t_out), .data_org(_add_map_x_88_data_org), .data_org_near(_add_map_x_88_data_org_near), .s_g(_add_map_x_88_s_g), .s_g_near(_add_map_x_88_s_g_near), .moto_org_near(_add_map_x_88_moto_org_near), .moto_org_near1(_add_map_x_88_moto_org_near1), .moto_org_near2(_add_map_x_88_moto_org_near2), .moto_org_near3(_add_map_x_88_moto_org_near3), .moto_org(_add_map_x_88_moto_org), .sg_up(_add_map_x_88_sg_up), .sg_down(_add_map_x_88_sg_down), .sg_left(_add_map_x_88_sg_left), .sg_right(_add_map_x_88_sg_right), .wall_t_in(_add_map_x_88_wall_t_in), .moto(_add_map_x_88_moto), .up(_add_map_x_88_up), .right(_add_map_x_88_right), .down(_add_map_x_88_down), .left(_add_map_x_88_left), .start(_add_map_x_88_start), .goal(_add_map_x_88_goal), .now(_add_map_x_88_now));
add_map add_map_x_87 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_87_add_exe), .data_out(_add_map_x_87_data_out), .data_out_index(_add_map_x_87_data_out_index), .data_near(_add_map_x_87_data_near), .wall_t_out(_add_map_x_87_wall_t_out), .data_org(_add_map_x_87_data_org), .data_org_near(_add_map_x_87_data_org_near), .s_g(_add_map_x_87_s_g), .s_g_near(_add_map_x_87_s_g_near), .moto_org_near(_add_map_x_87_moto_org_near), .moto_org_near1(_add_map_x_87_moto_org_near1), .moto_org_near2(_add_map_x_87_moto_org_near2), .moto_org_near3(_add_map_x_87_moto_org_near3), .moto_org(_add_map_x_87_moto_org), .sg_up(_add_map_x_87_sg_up), .sg_down(_add_map_x_87_sg_down), .sg_left(_add_map_x_87_sg_left), .sg_right(_add_map_x_87_sg_right), .wall_t_in(_add_map_x_87_wall_t_in), .moto(_add_map_x_87_moto), .up(_add_map_x_87_up), .right(_add_map_x_87_right), .down(_add_map_x_87_down), .left(_add_map_x_87_left), .start(_add_map_x_87_start), .goal(_add_map_x_87_goal), .now(_add_map_x_87_now));
add_map add_map_x_86 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_86_add_exe), .data_out(_add_map_x_86_data_out), .data_out_index(_add_map_x_86_data_out_index), .data_near(_add_map_x_86_data_near), .wall_t_out(_add_map_x_86_wall_t_out), .data_org(_add_map_x_86_data_org), .data_org_near(_add_map_x_86_data_org_near), .s_g(_add_map_x_86_s_g), .s_g_near(_add_map_x_86_s_g_near), .moto_org_near(_add_map_x_86_moto_org_near), .moto_org_near1(_add_map_x_86_moto_org_near1), .moto_org_near2(_add_map_x_86_moto_org_near2), .moto_org_near3(_add_map_x_86_moto_org_near3), .moto_org(_add_map_x_86_moto_org), .sg_up(_add_map_x_86_sg_up), .sg_down(_add_map_x_86_sg_down), .sg_left(_add_map_x_86_sg_left), .sg_right(_add_map_x_86_sg_right), .wall_t_in(_add_map_x_86_wall_t_in), .moto(_add_map_x_86_moto), .up(_add_map_x_86_up), .right(_add_map_x_86_right), .down(_add_map_x_86_down), .left(_add_map_x_86_left), .start(_add_map_x_86_start), .goal(_add_map_x_86_goal), .now(_add_map_x_86_now));
add_map add_map_x_85 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_85_add_exe), .data_out(_add_map_x_85_data_out), .data_out_index(_add_map_x_85_data_out_index), .data_near(_add_map_x_85_data_near), .wall_t_out(_add_map_x_85_wall_t_out), .data_org(_add_map_x_85_data_org), .data_org_near(_add_map_x_85_data_org_near), .s_g(_add_map_x_85_s_g), .s_g_near(_add_map_x_85_s_g_near), .moto_org_near(_add_map_x_85_moto_org_near), .moto_org_near1(_add_map_x_85_moto_org_near1), .moto_org_near2(_add_map_x_85_moto_org_near2), .moto_org_near3(_add_map_x_85_moto_org_near3), .moto_org(_add_map_x_85_moto_org), .sg_up(_add_map_x_85_sg_up), .sg_down(_add_map_x_85_sg_down), .sg_left(_add_map_x_85_sg_left), .sg_right(_add_map_x_85_sg_right), .wall_t_in(_add_map_x_85_wall_t_in), .moto(_add_map_x_85_moto), .up(_add_map_x_85_up), .right(_add_map_x_85_right), .down(_add_map_x_85_down), .left(_add_map_x_85_left), .start(_add_map_x_85_start), .goal(_add_map_x_85_goal), .now(_add_map_x_85_now));
add_map add_map_x_84 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_84_add_exe), .data_out(_add_map_x_84_data_out), .data_out_index(_add_map_x_84_data_out_index), .data_near(_add_map_x_84_data_near), .wall_t_out(_add_map_x_84_wall_t_out), .data_org(_add_map_x_84_data_org), .data_org_near(_add_map_x_84_data_org_near), .s_g(_add_map_x_84_s_g), .s_g_near(_add_map_x_84_s_g_near), .moto_org_near(_add_map_x_84_moto_org_near), .moto_org_near1(_add_map_x_84_moto_org_near1), .moto_org_near2(_add_map_x_84_moto_org_near2), .moto_org_near3(_add_map_x_84_moto_org_near3), .moto_org(_add_map_x_84_moto_org), .sg_up(_add_map_x_84_sg_up), .sg_down(_add_map_x_84_sg_down), .sg_left(_add_map_x_84_sg_left), .sg_right(_add_map_x_84_sg_right), .wall_t_in(_add_map_x_84_wall_t_in), .moto(_add_map_x_84_moto), .up(_add_map_x_84_up), .right(_add_map_x_84_right), .down(_add_map_x_84_down), .left(_add_map_x_84_left), .start(_add_map_x_84_start), .goal(_add_map_x_84_goal), .now(_add_map_x_84_now));
add_map add_map_x_83 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_83_add_exe), .data_out(_add_map_x_83_data_out), .data_out_index(_add_map_x_83_data_out_index), .data_near(_add_map_x_83_data_near), .wall_t_out(_add_map_x_83_wall_t_out), .data_org(_add_map_x_83_data_org), .data_org_near(_add_map_x_83_data_org_near), .s_g(_add_map_x_83_s_g), .s_g_near(_add_map_x_83_s_g_near), .moto_org_near(_add_map_x_83_moto_org_near), .moto_org_near1(_add_map_x_83_moto_org_near1), .moto_org_near2(_add_map_x_83_moto_org_near2), .moto_org_near3(_add_map_x_83_moto_org_near3), .moto_org(_add_map_x_83_moto_org), .sg_up(_add_map_x_83_sg_up), .sg_down(_add_map_x_83_sg_down), .sg_left(_add_map_x_83_sg_left), .sg_right(_add_map_x_83_sg_right), .wall_t_in(_add_map_x_83_wall_t_in), .moto(_add_map_x_83_moto), .up(_add_map_x_83_up), .right(_add_map_x_83_right), .down(_add_map_x_83_down), .left(_add_map_x_83_left), .start(_add_map_x_83_start), .goal(_add_map_x_83_goal), .now(_add_map_x_83_now));
add_map add_map_x_82 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_82_add_exe), .data_out(_add_map_x_82_data_out), .data_out_index(_add_map_x_82_data_out_index), .data_near(_add_map_x_82_data_near), .wall_t_out(_add_map_x_82_wall_t_out), .data_org(_add_map_x_82_data_org), .data_org_near(_add_map_x_82_data_org_near), .s_g(_add_map_x_82_s_g), .s_g_near(_add_map_x_82_s_g_near), .moto_org_near(_add_map_x_82_moto_org_near), .moto_org_near1(_add_map_x_82_moto_org_near1), .moto_org_near2(_add_map_x_82_moto_org_near2), .moto_org_near3(_add_map_x_82_moto_org_near3), .moto_org(_add_map_x_82_moto_org), .sg_up(_add_map_x_82_sg_up), .sg_down(_add_map_x_82_sg_down), .sg_left(_add_map_x_82_sg_left), .sg_right(_add_map_x_82_sg_right), .wall_t_in(_add_map_x_82_wall_t_in), .moto(_add_map_x_82_moto), .up(_add_map_x_82_up), .right(_add_map_x_82_right), .down(_add_map_x_82_down), .left(_add_map_x_82_left), .start(_add_map_x_82_start), .goal(_add_map_x_82_goal), .now(_add_map_x_82_now));
add_map add_map_x_81 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_81_add_exe), .data_out(_add_map_x_81_data_out), .data_out_index(_add_map_x_81_data_out_index), .data_near(_add_map_x_81_data_near), .wall_t_out(_add_map_x_81_wall_t_out), .data_org(_add_map_x_81_data_org), .data_org_near(_add_map_x_81_data_org_near), .s_g(_add_map_x_81_s_g), .s_g_near(_add_map_x_81_s_g_near), .moto_org_near(_add_map_x_81_moto_org_near), .moto_org_near1(_add_map_x_81_moto_org_near1), .moto_org_near2(_add_map_x_81_moto_org_near2), .moto_org_near3(_add_map_x_81_moto_org_near3), .moto_org(_add_map_x_81_moto_org), .sg_up(_add_map_x_81_sg_up), .sg_down(_add_map_x_81_sg_down), .sg_left(_add_map_x_81_sg_left), .sg_right(_add_map_x_81_sg_right), .wall_t_in(_add_map_x_81_wall_t_in), .moto(_add_map_x_81_moto), .up(_add_map_x_81_up), .right(_add_map_x_81_right), .down(_add_map_x_81_down), .left(_add_map_x_81_left), .start(_add_map_x_81_start), .goal(_add_map_x_81_goal), .now(_add_map_x_81_now));
add_map add_map_x_80 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_80_add_exe), .data_out(_add_map_x_80_data_out), .data_out_index(_add_map_x_80_data_out_index), .data_near(_add_map_x_80_data_near), .wall_t_out(_add_map_x_80_wall_t_out), .data_org(_add_map_x_80_data_org), .data_org_near(_add_map_x_80_data_org_near), .s_g(_add_map_x_80_s_g), .s_g_near(_add_map_x_80_s_g_near), .moto_org_near(_add_map_x_80_moto_org_near), .moto_org_near1(_add_map_x_80_moto_org_near1), .moto_org_near2(_add_map_x_80_moto_org_near2), .moto_org_near3(_add_map_x_80_moto_org_near3), .moto_org(_add_map_x_80_moto_org), .sg_up(_add_map_x_80_sg_up), .sg_down(_add_map_x_80_sg_down), .sg_left(_add_map_x_80_sg_left), .sg_right(_add_map_x_80_sg_right), .wall_t_in(_add_map_x_80_wall_t_in), .moto(_add_map_x_80_moto), .up(_add_map_x_80_up), .right(_add_map_x_80_right), .down(_add_map_x_80_down), .left(_add_map_x_80_left), .start(_add_map_x_80_start), .goal(_add_map_x_80_goal), .now(_add_map_x_80_now));
add_map add_map_x_79 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_79_add_exe), .data_out(_add_map_x_79_data_out), .data_out_index(_add_map_x_79_data_out_index), .data_near(_add_map_x_79_data_near), .wall_t_out(_add_map_x_79_wall_t_out), .data_org(_add_map_x_79_data_org), .data_org_near(_add_map_x_79_data_org_near), .s_g(_add_map_x_79_s_g), .s_g_near(_add_map_x_79_s_g_near), .moto_org_near(_add_map_x_79_moto_org_near), .moto_org_near1(_add_map_x_79_moto_org_near1), .moto_org_near2(_add_map_x_79_moto_org_near2), .moto_org_near3(_add_map_x_79_moto_org_near3), .moto_org(_add_map_x_79_moto_org), .sg_up(_add_map_x_79_sg_up), .sg_down(_add_map_x_79_sg_down), .sg_left(_add_map_x_79_sg_left), .sg_right(_add_map_x_79_sg_right), .wall_t_in(_add_map_x_79_wall_t_in), .moto(_add_map_x_79_moto), .up(_add_map_x_79_up), .right(_add_map_x_79_right), .down(_add_map_x_79_down), .left(_add_map_x_79_left), .start(_add_map_x_79_start), .goal(_add_map_x_79_goal), .now(_add_map_x_79_now));
add_map add_map_x_78 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_78_add_exe), .data_out(_add_map_x_78_data_out), .data_out_index(_add_map_x_78_data_out_index), .data_near(_add_map_x_78_data_near), .wall_t_out(_add_map_x_78_wall_t_out), .data_org(_add_map_x_78_data_org), .data_org_near(_add_map_x_78_data_org_near), .s_g(_add_map_x_78_s_g), .s_g_near(_add_map_x_78_s_g_near), .moto_org_near(_add_map_x_78_moto_org_near), .moto_org_near1(_add_map_x_78_moto_org_near1), .moto_org_near2(_add_map_x_78_moto_org_near2), .moto_org_near3(_add_map_x_78_moto_org_near3), .moto_org(_add_map_x_78_moto_org), .sg_up(_add_map_x_78_sg_up), .sg_down(_add_map_x_78_sg_down), .sg_left(_add_map_x_78_sg_left), .sg_right(_add_map_x_78_sg_right), .wall_t_in(_add_map_x_78_wall_t_in), .moto(_add_map_x_78_moto), .up(_add_map_x_78_up), .right(_add_map_x_78_right), .down(_add_map_x_78_down), .left(_add_map_x_78_left), .start(_add_map_x_78_start), .goal(_add_map_x_78_goal), .now(_add_map_x_78_now));
add_map add_map_x_77 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_77_add_exe), .data_out(_add_map_x_77_data_out), .data_out_index(_add_map_x_77_data_out_index), .data_near(_add_map_x_77_data_near), .wall_t_out(_add_map_x_77_wall_t_out), .data_org(_add_map_x_77_data_org), .data_org_near(_add_map_x_77_data_org_near), .s_g(_add_map_x_77_s_g), .s_g_near(_add_map_x_77_s_g_near), .moto_org_near(_add_map_x_77_moto_org_near), .moto_org_near1(_add_map_x_77_moto_org_near1), .moto_org_near2(_add_map_x_77_moto_org_near2), .moto_org_near3(_add_map_x_77_moto_org_near3), .moto_org(_add_map_x_77_moto_org), .sg_up(_add_map_x_77_sg_up), .sg_down(_add_map_x_77_sg_down), .sg_left(_add_map_x_77_sg_left), .sg_right(_add_map_x_77_sg_right), .wall_t_in(_add_map_x_77_wall_t_in), .moto(_add_map_x_77_moto), .up(_add_map_x_77_up), .right(_add_map_x_77_right), .down(_add_map_x_77_down), .left(_add_map_x_77_left), .start(_add_map_x_77_start), .goal(_add_map_x_77_goal), .now(_add_map_x_77_now));
add_map add_map_x_76 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_76_add_exe), .data_out(_add_map_x_76_data_out), .data_out_index(_add_map_x_76_data_out_index), .data_near(_add_map_x_76_data_near), .wall_t_out(_add_map_x_76_wall_t_out), .data_org(_add_map_x_76_data_org), .data_org_near(_add_map_x_76_data_org_near), .s_g(_add_map_x_76_s_g), .s_g_near(_add_map_x_76_s_g_near), .moto_org_near(_add_map_x_76_moto_org_near), .moto_org_near1(_add_map_x_76_moto_org_near1), .moto_org_near2(_add_map_x_76_moto_org_near2), .moto_org_near3(_add_map_x_76_moto_org_near3), .moto_org(_add_map_x_76_moto_org), .sg_up(_add_map_x_76_sg_up), .sg_down(_add_map_x_76_sg_down), .sg_left(_add_map_x_76_sg_left), .sg_right(_add_map_x_76_sg_right), .wall_t_in(_add_map_x_76_wall_t_in), .moto(_add_map_x_76_moto), .up(_add_map_x_76_up), .right(_add_map_x_76_right), .down(_add_map_x_76_down), .left(_add_map_x_76_left), .start(_add_map_x_76_start), .goal(_add_map_x_76_goal), .now(_add_map_x_76_now));
add_map add_map_x_75 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_75_add_exe), .data_out(_add_map_x_75_data_out), .data_out_index(_add_map_x_75_data_out_index), .data_near(_add_map_x_75_data_near), .wall_t_out(_add_map_x_75_wall_t_out), .data_org(_add_map_x_75_data_org), .data_org_near(_add_map_x_75_data_org_near), .s_g(_add_map_x_75_s_g), .s_g_near(_add_map_x_75_s_g_near), .moto_org_near(_add_map_x_75_moto_org_near), .moto_org_near1(_add_map_x_75_moto_org_near1), .moto_org_near2(_add_map_x_75_moto_org_near2), .moto_org_near3(_add_map_x_75_moto_org_near3), .moto_org(_add_map_x_75_moto_org), .sg_up(_add_map_x_75_sg_up), .sg_down(_add_map_x_75_sg_down), .sg_left(_add_map_x_75_sg_left), .sg_right(_add_map_x_75_sg_right), .wall_t_in(_add_map_x_75_wall_t_in), .moto(_add_map_x_75_moto), .up(_add_map_x_75_up), .right(_add_map_x_75_right), .down(_add_map_x_75_down), .left(_add_map_x_75_left), .start(_add_map_x_75_start), .goal(_add_map_x_75_goal), .now(_add_map_x_75_now));
add_map add_map_x_74 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_74_add_exe), .data_out(_add_map_x_74_data_out), .data_out_index(_add_map_x_74_data_out_index), .data_near(_add_map_x_74_data_near), .wall_t_out(_add_map_x_74_wall_t_out), .data_org(_add_map_x_74_data_org), .data_org_near(_add_map_x_74_data_org_near), .s_g(_add_map_x_74_s_g), .s_g_near(_add_map_x_74_s_g_near), .moto_org_near(_add_map_x_74_moto_org_near), .moto_org_near1(_add_map_x_74_moto_org_near1), .moto_org_near2(_add_map_x_74_moto_org_near2), .moto_org_near3(_add_map_x_74_moto_org_near3), .moto_org(_add_map_x_74_moto_org), .sg_up(_add_map_x_74_sg_up), .sg_down(_add_map_x_74_sg_down), .sg_left(_add_map_x_74_sg_left), .sg_right(_add_map_x_74_sg_right), .wall_t_in(_add_map_x_74_wall_t_in), .moto(_add_map_x_74_moto), .up(_add_map_x_74_up), .right(_add_map_x_74_right), .down(_add_map_x_74_down), .left(_add_map_x_74_left), .start(_add_map_x_74_start), .goal(_add_map_x_74_goal), .now(_add_map_x_74_now));
add_map add_map_x_73 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_73_add_exe), .data_out(_add_map_x_73_data_out), .data_out_index(_add_map_x_73_data_out_index), .data_near(_add_map_x_73_data_near), .wall_t_out(_add_map_x_73_wall_t_out), .data_org(_add_map_x_73_data_org), .data_org_near(_add_map_x_73_data_org_near), .s_g(_add_map_x_73_s_g), .s_g_near(_add_map_x_73_s_g_near), .moto_org_near(_add_map_x_73_moto_org_near), .moto_org_near1(_add_map_x_73_moto_org_near1), .moto_org_near2(_add_map_x_73_moto_org_near2), .moto_org_near3(_add_map_x_73_moto_org_near3), .moto_org(_add_map_x_73_moto_org), .sg_up(_add_map_x_73_sg_up), .sg_down(_add_map_x_73_sg_down), .sg_left(_add_map_x_73_sg_left), .sg_right(_add_map_x_73_sg_right), .wall_t_in(_add_map_x_73_wall_t_in), .moto(_add_map_x_73_moto), .up(_add_map_x_73_up), .right(_add_map_x_73_right), .down(_add_map_x_73_down), .left(_add_map_x_73_left), .start(_add_map_x_73_start), .goal(_add_map_x_73_goal), .now(_add_map_x_73_now));
add_map add_map_x_72 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_72_add_exe), .data_out(_add_map_x_72_data_out), .data_out_index(_add_map_x_72_data_out_index), .data_near(_add_map_x_72_data_near), .wall_t_out(_add_map_x_72_wall_t_out), .data_org(_add_map_x_72_data_org), .data_org_near(_add_map_x_72_data_org_near), .s_g(_add_map_x_72_s_g), .s_g_near(_add_map_x_72_s_g_near), .moto_org_near(_add_map_x_72_moto_org_near), .moto_org_near1(_add_map_x_72_moto_org_near1), .moto_org_near2(_add_map_x_72_moto_org_near2), .moto_org_near3(_add_map_x_72_moto_org_near3), .moto_org(_add_map_x_72_moto_org), .sg_up(_add_map_x_72_sg_up), .sg_down(_add_map_x_72_sg_down), .sg_left(_add_map_x_72_sg_left), .sg_right(_add_map_x_72_sg_right), .wall_t_in(_add_map_x_72_wall_t_in), .moto(_add_map_x_72_moto), .up(_add_map_x_72_up), .right(_add_map_x_72_right), .down(_add_map_x_72_down), .left(_add_map_x_72_left), .start(_add_map_x_72_start), .goal(_add_map_x_72_goal), .now(_add_map_x_72_now));
add_map add_map_x_71 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_71_add_exe), .data_out(_add_map_x_71_data_out), .data_out_index(_add_map_x_71_data_out_index), .data_near(_add_map_x_71_data_near), .wall_t_out(_add_map_x_71_wall_t_out), .data_org(_add_map_x_71_data_org), .data_org_near(_add_map_x_71_data_org_near), .s_g(_add_map_x_71_s_g), .s_g_near(_add_map_x_71_s_g_near), .moto_org_near(_add_map_x_71_moto_org_near), .moto_org_near1(_add_map_x_71_moto_org_near1), .moto_org_near2(_add_map_x_71_moto_org_near2), .moto_org_near3(_add_map_x_71_moto_org_near3), .moto_org(_add_map_x_71_moto_org), .sg_up(_add_map_x_71_sg_up), .sg_down(_add_map_x_71_sg_down), .sg_left(_add_map_x_71_sg_left), .sg_right(_add_map_x_71_sg_right), .wall_t_in(_add_map_x_71_wall_t_in), .moto(_add_map_x_71_moto), .up(_add_map_x_71_up), .right(_add_map_x_71_right), .down(_add_map_x_71_down), .left(_add_map_x_71_left), .start(_add_map_x_71_start), .goal(_add_map_x_71_goal), .now(_add_map_x_71_now));
add_map add_map_x_70 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_70_add_exe), .data_out(_add_map_x_70_data_out), .data_out_index(_add_map_x_70_data_out_index), .data_near(_add_map_x_70_data_near), .wall_t_out(_add_map_x_70_wall_t_out), .data_org(_add_map_x_70_data_org), .data_org_near(_add_map_x_70_data_org_near), .s_g(_add_map_x_70_s_g), .s_g_near(_add_map_x_70_s_g_near), .moto_org_near(_add_map_x_70_moto_org_near), .moto_org_near1(_add_map_x_70_moto_org_near1), .moto_org_near2(_add_map_x_70_moto_org_near2), .moto_org_near3(_add_map_x_70_moto_org_near3), .moto_org(_add_map_x_70_moto_org), .sg_up(_add_map_x_70_sg_up), .sg_down(_add_map_x_70_sg_down), .sg_left(_add_map_x_70_sg_left), .sg_right(_add_map_x_70_sg_right), .wall_t_in(_add_map_x_70_wall_t_in), .moto(_add_map_x_70_moto), .up(_add_map_x_70_up), .right(_add_map_x_70_right), .down(_add_map_x_70_down), .left(_add_map_x_70_left), .start(_add_map_x_70_start), .goal(_add_map_x_70_goal), .now(_add_map_x_70_now));
add_map add_map_x_69 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_69_add_exe), .data_out(_add_map_x_69_data_out), .data_out_index(_add_map_x_69_data_out_index), .data_near(_add_map_x_69_data_near), .wall_t_out(_add_map_x_69_wall_t_out), .data_org(_add_map_x_69_data_org), .data_org_near(_add_map_x_69_data_org_near), .s_g(_add_map_x_69_s_g), .s_g_near(_add_map_x_69_s_g_near), .moto_org_near(_add_map_x_69_moto_org_near), .moto_org_near1(_add_map_x_69_moto_org_near1), .moto_org_near2(_add_map_x_69_moto_org_near2), .moto_org_near3(_add_map_x_69_moto_org_near3), .moto_org(_add_map_x_69_moto_org), .sg_up(_add_map_x_69_sg_up), .sg_down(_add_map_x_69_sg_down), .sg_left(_add_map_x_69_sg_left), .sg_right(_add_map_x_69_sg_right), .wall_t_in(_add_map_x_69_wall_t_in), .moto(_add_map_x_69_moto), .up(_add_map_x_69_up), .right(_add_map_x_69_right), .down(_add_map_x_69_down), .left(_add_map_x_69_left), .start(_add_map_x_69_start), .goal(_add_map_x_69_goal), .now(_add_map_x_69_now));
add_map add_map_x_68 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_68_add_exe), .data_out(_add_map_x_68_data_out), .data_out_index(_add_map_x_68_data_out_index), .data_near(_add_map_x_68_data_near), .wall_t_out(_add_map_x_68_wall_t_out), .data_org(_add_map_x_68_data_org), .data_org_near(_add_map_x_68_data_org_near), .s_g(_add_map_x_68_s_g), .s_g_near(_add_map_x_68_s_g_near), .moto_org_near(_add_map_x_68_moto_org_near), .moto_org_near1(_add_map_x_68_moto_org_near1), .moto_org_near2(_add_map_x_68_moto_org_near2), .moto_org_near3(_add_map_x_68_moto_org_near3), .moto_org(_add_map_x_68_moto_org), .sg_up(_add_map_x_68_sg_up), .sg_down(_add_map_x_68_sg_down), .sg_left(_add_map_x_68_sg_left), .sg_right(_add_map_x_68_sg_right), .wall_t_in(_add_map_x_68_wall_t_in), .moto(_add_map_x_68_moto), .up(_add_map_x_68_up), .right(_add_map_x_68_right), .down(_add_map_x_68_down), .left(_add_map_x_68_left), .start(_add_map_x_68_start), .goal(_add_map_x_68_goal), .now(_add_map_x_68_now));
add_map add_map_x_67 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_67_add_exe), .data_out(_add_map_x_67_data_out), .data_out_index(_add_map_x_67_data_out_index), .data_near(_add_map_x_67_data_near), .wall_t_out(_add_map_x_67_wall_t_out), .data_org(_add_map_x_67_data_org), .data_org_near(_add_map_x_67_data_org_near), .s_g(_add_map_x_67_s_g), .s_g_near(_add_map_x_67_s_g_near), .moto_org_near(_add_map_x_67_moto_org_near), .moto_org_near1(_add_map_x_67_moto_org_near1), .moto_org_near2(_add_map_x_67_moto_org_near2), .moto_org_near3(_add_map_x_67_moto_org_near3), .moto_org(_add_map_x_67_moto_org), .sg_up(_add_map_x_67_sg_up), .sg_down(_add_map_x_67_sg_down), .sg_left(_add_map_x_67_sg_left), .sg_right(_add_map_x_67_sg_right), .wall_t_in(_add_map_x_67_wall_t_in), .moto(_add_map_x_67_moto), .up(_add_map_x_67_up), .right(_add_map_x_67_right), .down(_add_map_x_67_down), .left(_add_map_x_67_left), .start(_add_map_x_67_start), .goal(_add_map_x_67_goal), .now(_add_map_x_67_now));
add_map add_map_x_66 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_66_add_exe), .data_out(_add_map_x_66_data_out), .data_out_index(_add_map_x_66_data_out_index), .data_near(_add_map_x_66_data_near), .wall_t_out(_add_map_x_66_wall_t_out), .data_org(_add_map_x_66_data_org), .data_org_near(_add_map_x_66_data_org_near), .s_g(_add_map_x_66_s_g), .s_g_near(_add_map_x_66_s_g_near), .moto_org_near(_add_map_x_66_moto_org_near), .moto_org_near1(_add_map_x_66_moto_org_near1), .moto_org_near2(_add_map_x_66_moto_org_near2), .moto_org_near3(_add_map_x_66_moto_org_near3), .moto_org(_add_map_x_66_moto_org), .sg_up(_add_map_x_66_sg_up), .sg_down(_add_map_x_66_sg_down), .sg_left(_add_map_x_66_sg_left), .sg_right(_add_map_x_66_sg_right), .wall_t_in(_add_map_x_66_wall_t_in), .moto(_add_map_x_66_moto), .up(_add_map_x_66_up), .right(_add_map_x_66_right), .down(_add_map_x_66_down), .left(_add_map_x_66_left), .start(_add_map_x_66_start), .goal(_add_map_x_66_goal), .now(_add_map_x_66_now));
add_map add_map_x_65 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_65_add_exe), .data_out(_add_map_x_65_data_out), .data_out_index(_add_map_x_65_data_out_index), .data_near(_add_map_x_65_data_near), .wall_t_out(_add_map_x_65_wall_t_out), .data_org(_add_map_x_65_data_org), .data_org_near(_add_map_x_65_data_org_near), .s_g(_add_map_x_65_s_g), .s_g_near(_add_map_x_65_s_g_near), .moto_org_near(_add_map_x_65_moto_org_near), .moto_org_near1(_add_map_x_65_moto_org_near1), .moto_org_near2(_add_map_x_65_moto_org_near2), .moto_org_near3(_add_map_x_65_moto_org_near3), .moto_org(_add_map_x_65_moto_org), .sg_up(_add_map_x_65_sg_up), .sg_down(_add_map_x_65_sg_down), .sg_left(_add_map_x_65_sg_left), .sg_right(_add_map_x_65_sg_right), .wall_t_in(_add_map_x_65_wall_t_in), .moto(_add_map_x_65_moto), .up(_add_map_x_65_up), .right(_add_map_x_65_right), .down(_add_map_x_65_down), .left(_add_map_x_65_left), .start(_add_map_x_65_start), .goal(_add_map_x_65_goal), .now(_add_map_x_65_now));
add_map add_map_x_64 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_64_add_exe), .data_out(_add_map_x_64_data_out), .data_out_index(_add_map_x_64_data_out_index), .data_near(_add_map_x_64_data_near), .wall_t_out(_add_map_x_64_wall_t_out), .data_org(_add_map_x_64_data_org), .data_org_near(_add_map_x_64_data_org_near), .s_g(_add_map_x_64_s_g), .s_g_near(_add_map_x_64_s_g_near), .moto_org_near(_add_map_x_64_moto_org_near), .moto_org_near1(_add_map_x_64_moto_org_near1), .moto_org_near2(_add_map_x_64_moto_org_near2), .moto_org_near3(_add_map_x_64_moto_org_near3), .moto_org(_add_map_x_64_moto_org), .sg_up(_add_map_x_64_sg_up), .sg_down(_add_map_x_64_sg_down), .sg_left(_add_map_x_64_sg_left), .sg_right(_add_map_x_64_sg_right), .wall_t_in(_add_map_x_64_wall_t_in), .moto(_add_map_x_64_moto), .up(_add_map_x_64_up), .right(_add_map_x_64_right), .down(_add_map_x_64_down), .left(_add_map_x_64_left), .start(_add_map_x_64_start), .goal(_add_map_x_64_goal), .now(_add_map_x_64_now));
add_map add_map_x_63 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_63_add_exe), .data_out(_add_map_x_63_data_out), .data_out_index(_add_map_x_63_data_out_index), .data_near(_add_map_x_63_data_near), .wall_t_out(_add_map_x_63_wall_t_out), .data_org(_add_map_x_63_data_org), .data_org_near(_add_map_x_63_data_org_near), .s_g(_add_map_x_63_s_g), .s_g_near(_add_map_x_63_s_g_near), .moto_org_near(_add_map_x_63_moto_org_near), .moto_org_near1(_add_map_x_63_moto_org_near1), .moto_org_near2(_add_map_x_63_moto_org_near2), .moto_org_near3(_add_map_x_63_moto_org_near3), .moto_org(_add_map_x_63_moto_org), .sg_up(_add_map_x_63_sg_up), .sg_down(_add_map_x_63_sg_down), .sg_left(_add_map_x_63_sg_left), .sg_right(_add_map_x_63_sg_right), .wall_t_in(_add_map_x_63_wall_t_in), .moto(_add_map_x_63_moto), .up(_add_map_x_63_up), .right(_add_map_x_63_right), .down(_add_map_x_63_down), .left(_add_map_x_63_left), .start(_add_map_x_63_start), .goal(_add_map_x_63_goal), .now(_add_map_x_63_now));
add_map add_map_x_62 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_62_add_exe), .data_out(_add_map_x_62_data_out), .data_out_index(_add_map_x_62_data_out_index), .data_near(_add_map_x_62_data_near), .wall_t_out(_add_map_x_62_wall_t_out), .data_org(_add_map_x_62_data_org), .data_org_near(_add_map_x_62_data_org_near), .s_g(_add_map_x_62_s_g), .s_g_near(_add_map_x_62_s_g_near), .moto_org_near(_add_map_x_62_moto_org_near), .moto_org_near1(_add_map_x_62_moto_org_near1), .moto_org_near2(_add_map_x_62_moto_org_near2), .moto_org_near3(_add_map_x_62_moto_org_near3), .moto_org(_add_map_x_62_moto_org), .sg_up(_add_map_x_62_sg_up), .sg_down(_add_map_x_62_sg_down), .sg_left(_add_map_x_62_sg_left), .sg_right(_add_map_x_62_sg_right), .wall_t_in(_add_map_x_62_wall_t_in), .moto(_add_map_x_62_moto), .up(_add_map_x_62_up), .right(_add_map_x_62_right), .down(_add_map_x_62_down), .left(_add_map_x_62_left), .start(_add_map_x_62_start), .goal(_add_map_x_62_goal), .now(_add_map_x_62_now));
add_map add_map_x_61 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_61_add_exe), .data_out(_add_map_x_61_data_out), .data_out_index(_add_map_x_61_data_out_index), .data_near(_add_map_x_61_data_near), .wall_t_out(_add_map_x_61_wall_t_out), .data_org(_add_map_x_61_data_org), .data_org_near(_add_map_x_61_data_org_near), .s_g(_add_map_x_61_s_g), .s_g_near(_add_map_x_61_s_g_near), .moto_org_near(_add_map_x_61_moto_org_near), .moto_org_near1(_add_map_x_61_moto_org_near1), .moto_org_near2(_add_map_x_61_moto_org_near2), .moto_org_near3(_add_map_x_61_moto_org_near3), .moto_org(_add_map_x_61_moto_org), .sg_up(_add_map_x_61_sg_up), .sg_down(_add_map_x_61_sg_down), .sg_left(_add_map_x_61_sg_left), .sg_right(_add_map_x_61_sg_right), .wall_t_in(_add_map_x_61_wall_t_in), .moto(_add_map_x_61_moto), .up(_add_map_x_61_up), .right(_add_map_x_61_right), .down(_add_map_x_61_down), .left(_add_map_x_61_left), .start(_add_map_x_61_start), .goal(_add_map_x_61_goal), .now(_add_map_x_61_now));
add_map add_map_x_60 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_60_add_exe), .data_out(_add_map_x_60_data_out), .data_out_index(_add_map_x_60_data_out_index), .data_near(_add_map_x_60_data_near), .wall_t_out(_add_map_x_60_wall_t_out), .data_org(_add_map_x_60_data_org), .data_org_near(_add_map_x_60_data_org_near), .s_g(_add_map_x_60_s_g), .s_g_near(_add_map_x_60_s_g_near), .moto_org_near(_add_map_x_60_moto_org_near), .moto_org_near1(_add_map_x_60_moto_org_near1), .moto_org_near2(_add_map_x_60_moto_org_near2), .moto_org_near3(_add_map_x_60_moto_org_near3), .moto_org(_add_map_x_60_moto_org), .sg_up(_add_map_x_60_sg_up), .sg_down(_add_map_x_60_sg_down), .sg_left(_add_map_x_60_sg_left), .sg_right(_add_map_x_60_sg_right), .wall_t_in(_add_map_x_60_wall_t_in), .moto(_add_map_x_60_moto), .up(_add_map_x_60_up), .right(_add_map_x_60_right), .down(_add_map_x_60_down), .left(_add_map_x_60_left), .start(_add_map_x_60_start), .goal(_add_map_x_60_goal), .now(_add_map_x_60_now));
add_map add_map_x_59 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_59_add_exe), .data_out(_add_map_x_59_data_out), .data_out_index(_add_map_x_59_data_out_index), .data_near(_add_map_x_59_data_near), .wall_t_out(_add_map_x_59_wall_t_out), .data_org(_add_map_x_59_data_org), .data_org_near(_add_map_x_59_data_org_near), .s_g(_add_map_x_59_s_g), .s_g_near(_add_map_x_59_s_g_near), .moto_org_near(_add_map_x_59_moto_org_near), .moto_org_near1(_add_map_x_59_moto_org_near1), .moto_org_near2(_add_map_x_59_moto_org_near2), .moto_org_near3(_add_map_x_59_moto_org_near3), .moto_org(_add_map_x_59_moto_org), .sg_up(_add_map_x_59_sg_up), .sg_down(_add_map_x_59_sg_down), .sg_left(_add_map_x_59_sg_left), .sg_right(_add_map_x_59_sg_right), .wall_t_in(_add_map_x_59_wall_t_in), .moto(_add_map_x_59_moto), .up(_add_map_x_59_up), .right(_add_map_x_59_right), .down(_add_map_x_59_down), .left(_add_map_x_59_left), .start(_add_map_x_59_start), .goal(_add_map_x_59_goal), .now(_add_map_x_59_now));
add_map add_map_x_58 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_58_add_exe), .data_out(_add_map_x_58_data_out), .data_out_index(_add_map_x_58_data_out_index), .data_near(_add_map_x_58_data_near), .wall_t_out(_add_map_x_58_wall_t_out), .data_org(_add_map_x_58_data_org), .data_org_near(_add_map_x_58_data_org_near), .s_g(_add_map_x_58_s_g), .s_g_near(_add_map_x_58_s_g_near), .moto_org_near(_add_map_x_58_moto_org_near), .moto_org_near1(_add_map_x_58_moto_org_near1), .moto_org_near2(_add_map_x_58_moto_org_near2), .moto_org_near3(_add_map_x_58_moto_org_near3), .moto_org(_add_map_x_58_moto_org), .sg_up(_add_map_x_58_sg_up), .sg_down(_add_map_x_58_sg_down), .sg_left(_add_map_x_58_sg_left), .sg_right(_add_map_x_58_sg_right), .wall_t_in(_add_map_x_58_wall_t_in), .moto(_add_map_x_58_moto), .up(_add_map_x_58_up), .right(_add_map_x_58_right), .down(_add_map_x_58_down), .left(_add_map_x_58_left), .start(_add_map_x_58_start), .goal(_add_map_x_58_goal), .now(_add_map_x_58_now));
add_map add_map_x_57 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_57_add_exe), .data_out(_add_map_x_57_data_out), .data_out_index(_add_map_x_57_data_out_index), .data_near(_add_map_x_57_data_near), .wall_t_out(_add_map_x_57_wall_t_out), .data_org(_add_map_x_57_data_org), .data_org_near(_add_map_x_57_data_org_near), .s_g(_add_map_x_57_s_g), .s_g_near(_add_map_x_57_s_g_near), .moto_org_near(_add_map_x_57_moto_org_near), .moto_org_near1(_add_map_x_57_moto_org_near1), .moto_org_near2(_add_map_x_57_moto_org_near2), .moto_org_near3(_add_map_x_57_moto_org_near3), .moto_org(_add_map_x_57_moto_org), .sg_up(_add_map_x_57_sg_up), .sg_down(_add_map_x_57_sg_down), .sg_left(_add_map_x_57_sg_left), .sg_right(_add_map_x_57_sg_right), .wall_t_in(_add_map_x_57_wall_t_in), .moto(_add_map_x_57_moto), .up(_add_map_x_57_up), .right(_add_map_x_57_right), .down(_add_map_x_57_down), .left(_add_map_x_57_left), .start(_add_map_x_57_start), .goal(_add_map_x_57_goal), .now(_add_map_x_57_now));
add_map add_map_x_56 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_56_add_exe), .data_out(_add_map_x_56_data_out), .data_out_index(_add_map_x_56_data_out_index), .data_near(_add_map_x_56_data_near), .wall_t_out(_add_map_x_56_wall_t_out), .data_org(_add_map_x_56_data_org), .data_org_near(_add_map_x_56_data_org_near), .s_g(_add_map_x_56_s_g), .s_g_near(_add_map_x_56_s_g_near), .moto_org_near(_add_map_x_56_moto_org_near), .moto_org_near1(_add_map_x_56_moto_org_near1), .moto_org_near2(_add_map_x_56_moto_org_near2), .moto_org_near3(_add_map_x_56_moto_org_near3), .moto_org(_add_map_x_56_moto_org), .sg_up(_add_map_x_56_sg_up), .sg_down(_add_map_x_56_sg_down), .sg_left(_add_map_x_56_sg_left), .sg_right(_add_map_x_56_sg_right), .wall_t_in(_add_map_x_56_wall_t_in), .moto(_add_map_x_56_moto), .up(_add_map_x_56_up), .right(_add_map_x_56_right), .down(_add_map_x_56_down), .left(_add_map_x_56_left), .start(_add_map_x_56_start), .goal(_add_map_x_56_goal), .now(_add_map_x_56_now));
add_map add_map_x_55 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_55_add_exe), .data_out(_add_map_x_55_data_out), .data_out_index(_add_map_x_55_data_out_index), .data_near(_add_map_x_55_data_near), .wall_t_out(_add_map_x_55_wall_t_out), .data_org(_add_map_x_55_data_org), .data_org_near(_add_map_x_55_data_org_near), .s_g(_add_map_x_55_s_g), .s_g_near(_add_map_x_55_s_g_near), .moto_org_near(_add_map_x_55_moto_org_near), .moto_org_near1(_add_map_x_55_moto_org_near1), .moto_org_near2(_add_map_x_55_moto_org_near2), .moto_org_near3(_add_map_x_55_moto_org_near3), .moto_org(_add_map_x_55_moto_org), .sg_up(_add_map_x_55_sg_up), .sg_down(_add_map_x_55_sg_down), .sg_left(_add_map_x_55_sg_left), .sg_right(_add_map_x_55_sg_right), .wall_t_in(_add_map_x_55_wall_t_in), .moto(_add_map_x_55_moto), .up(_add_map_x_55_up), .right(_add_map_x_55_right), .down(_add_map_x_55_down), .left(_add_map_x_55_left), .start(_add_map_x_55_start), .goal(_add_map_x_55_goal), .now(_add_map_x_55_now));
add_map add_map_x_54 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_54_add_exe), .data_out(_add_map_x_54_data_out), .data_out_index(_add_map_x_54_data_out_index), .data_near(_add_map_x_54_data_near), .wall_t_out(_add_map_x_54_wall_t_out), .data_org(_add_map_x_54_data_org), .data_org_near(_add_map_x_54_data_org_near), .s_g(_add_map_x_54_s_g), .s_g_near(_add_map_x_54_s_g_near), .moto_org_near(_add_map_x_54_moto_org_near), .moto_org_near1(_add_map_x_54_moto_org_near1), .moto_org_near2(_add_map_x_54_moto_org_near2), .moto_org_near3(_add_map_x_54_moto_org_near3), .moto_org(_add_map_x_54_moto_org), .sg_up(_add_map_x_54_sg_up), .sg_down(_add_map_x_54_sg_down), .sg_left(_add_map_x_54_sg_left), .sg_right(_add_map_x_54_sg_right), .wall_t_in(_add_map_x_54_wall_t_in), .moto(_add_map_x_54_moto), .up(_add_map_x_54_up), .right(_add_map_x_54_right), .down(_add_map_x_54_down), .left(_add_map_x_54_left), .start(_add_map_x_54_start), .goal(_add_map_x_54_goal), .now(_add_map_x_54_now));
add_map add_map_x_53 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_53_add_exe), .data_out(_add_map_x_53_data_out), .data_out_index(_add_map_x_53_data_out_index), .data_near(_add_map_x_53_data_near), .wall_t_out(_add_map_x_53_wall_t_out), .data_org(_add_map_x_53_data_org), .data_org_near(_add_map_x_53_data_org_near), .s_g(_add_map_x_53_s_g), .s_g_near(_add_map_x_53_s_g_near), .moto_org_near(_add_map_x_53_moto_org_near), .moto_org_near1(_add_map_x_53_moto_org_near1), .moto_org_near2(_add_map_x_53_moto_org_near2), .moto_org_near3(_add_map_x_53_moto_org_near3), .moto_org(_add_map_x_53_moto_org), .sg_up(_add_map_x_53_sg_up), .sg_down(_add_map_x_53_sg_down), .sg_left(_add_map_x_53_sg_left), .sg_right(_add_map_x_53_sg_right), .wall_t_in(_add_map_x_53_wall_t_in), .moto(_add_map_x_53_moto), .up(_add_map_x_53_up), .right(_add_map_x_53_right), .down(_add_map_x_53_down), .left(_add_map_x_53_left), .start(_add_map_x_53_start), .goal(_add_map_x_53_goal), .now(_add_map_x_53_now));
add_map add_map_x_52 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_52_add_exe), .data_out(_add_map_x_52_data_out), .data_out_index(_add_map_x_52_data_out_index), .data_near(_add_map_x_52_data_near), .wall_t_out(_add_map_x_52_wall_t_out), .data_org(_add_map_x_52_data_org), .data_org_near(_add_map_x_52_data_org_near), .s_g(_add_map_x_52_s_g), .s_g_near(_add_map_x_52_s_g_near), .moto_org_near(_add_map_x_52_moto_org_near), .moto_org_near1(_add_map_x_52_moto_org_near1), .moto_org_near2(_add_map_x_52_moto_org_near2), .moto_org_near3(_add_map_x_52_moto_org_near3), .moto_org(_add_map_x_52_moto_org), .sg_up(_add_map_x_52_sg_up), .sg_down(_add_map_x_52_sg_down), .sg_left(_add_map_x_52_sg_left), .sg_right(_add_map_x_52_sg_right), .wall_t_in(_add_map_x_52_wall_t_in), .moto(_add_map_x_52_moto), .up(_add_map_x_52_up), .right(_add_map_x_52_right), .down(_add_map_x_52_down), .left(_add_map_x_52_left), .start(_add_map_x_52_start), .goal(_add_map_x_52_goal), .now(_add_map_x_52_now));
add_map add_map_x_51 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_51_add_exe), .data_out(_add_map_x_51_data_out), .data_out_index(_add_map_x_51_data_out_index), .data_near(_add_map_x_51_data_near), .wall_t_out(_add_map_x_51_wall_t_out), .data_org(_add_map_x_51_data_org), .data_org_near(_add_map_x_51_data_org_near), .s_g(_add_map_x_51_s_g), .s_g_near(_add_map_x_51_s_g_near), .moto_org_near(_add_map_x_51_moto_org_near), .moto_org_near1(_add_map_x_51_moto_org_near1), .moto_org_near2(_add_map_x_51_moto_org_near2), .moto_org_near3(_add_map_x_51_moto_org_near3), .moto_org(_add_map_x_51_moto_org), .sg_up(_add_map_x_51_sg_up), .sg_down(_add_map_x_51_sg_down), .sg_left(_add_map_x_51_sg_left), .sg_right(_add_map_x_51_sg_right), .wall_t_in(_add_map_x_51_wall_t_in), .moto(_add_map_x_51_moto), .up(_add_map_x_51_up), .right(_add_map_x_51_right), .down(_add_map_x_51_down), .left(_add_map_x_51_left), .start(_add_map_x_51_start), .goal(_add_map_x_51_goal), .now(_add_map_x_51_now));
add_map add_map_x_50 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_50_add_exe), .data_out(_add_map_x_50_data_out), .data_out_index(_add_map_x_50_data_out_index), .data_near(_add_map_x_50_data_near), .wall_t_out(_add_map_x_50_wall_t_out), .data_org(_add_map_x_50_data_org), .data_org_near(_add_map_x_50_data_org_near), .s_g(_add_map_x_50_s_g), .s_g_near(_add_map_x_50_s_g_near), .moto_org_near(_add_map_x_50_moto_org_near), .moto_org_near1(_add_map_x_50_moto_org_near1), .moto_org_near2(_add_map_x_50_moto_org_near2), .moto_org_near3(_add_map_x_50_moto_org_near3), .moto_org(_add_map_x_50_moto_org), .sg_up(_add_map_x_50_sg_up), .sg_down(_add_map_x_50_sg_down), .sg_left(_add_map_x_50_sg_left), .sg_right(_add_map_x_50_sg_right), .wall_t_in(_add_map_x_50_wall_t_in), .moto(_add_map_x_50_moto), .up(_add_map_x_50_up), .right(_add_map_x_50_right), .down(_add_map_x_50_down), .left(_add_map_x_50_left), .start(_add_map_x_50_start), .goal(_add_map_x_50_goal), .now(_add_map_x_50_now));
add_map add_map_x_49 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_49_add_exe), .data_out(_add_map_x_49_data_out), .data_out_index(_add_map_x_49_data_out_index), .data_near(_add_map_x_49_data_near), .wall_t_out(_add_map_x_49_wall_t_out), .data_org(_add_map_x_49_data_org), .data_org_near(_add_map_x_49_data_org_near), .s_g(_add_map_x_49_s_g), .s_g_near(_add_map_x_49_s_g_near), .moto_org_near(_add_map_x_49_moto_org_near), .moto_org_near1(_add_map_x_49_moto_org_near1), .moto_org_near2(_add_map_x_49_moto_org_near2), .moto_org_near3(_add_map_x_49_moto_org_near3), .moto_org(_add_map_x_49_moto_org), .sg_up(_add_map_x_49_sg_up), .sg_down(_add_map_x_49_sg_down), .sg_left(_add_map_x_49_sg_left), .sg_right(_add_map_x_49_sg_right), .wall_t_in(_add_map_x_49_wall_t_in), .moto(_add_map_x_49_moto), .up(_add_map_x_49_up), .right(_add_map_x_49_right), .down(_add_map_x_49_down), .left(_add_map_x_49_left), .start(_add_map_x_49_start), .goal(_add_map_x_49_goal), .now(_add_map_x_49_now));
add_map add_map_x_48 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_48_add_exe), .data_out(_add_map_x_48_data_out), .data_out_index(_add_map_x_48_data_out_index), .data_near(_add_map_x_48_data_near), .wall_t_out(_add_map_x_48_wall_t_out), .data_org(_add_map_x_48_data_org), .data_org_near(_add_map_x_48_data_org_near), .s_g(_add_map_x_48_s_g), .s_g_near(_add_map_x_48_s_g_near), .moto_org_near(_add_map_x_48_moto_org_near), .moto_org_near1(_add_map_x_48_moto_org_near1), .moto_org_near2(_add_map_x_48_moto_org_near2), .moto_org_near3(_add_map_x_48_moto_org_near3), .moto_org(_add_map_x_48_moto_org), .sg_up(_add_map_x_48_sg_up), .sg_down(_add_map_x_48_sg_down), .sg_left(_add_map_x_48_sg_left), .sg_right(_add_map_x_48_sg_right), .wall_t_in(_add_map_x_48_wall_t_in), .moto(_add_map_x_48_moto), .up(_add_map_x_48_up), .right(_add_map_x_48_right), .down(_add_map_x_48_down), .left(_add_map_x_48_left), .start(_add_map_x_48_start), .goal(_add_map_x_48_goal), .now(_add_map_x_48_now));
add_map add_map_x_47 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_47_add_exe), .data_out(_add_map_x_47_data_out), .data_out_index(_add_map_x_47_data_out_index), .data_near(_add_map_x_47_data_near), .wall_t_out(_add_map_x_47_wall_t_out), .data_org(_add_map_x_47_data_org), .data_org_near(_add_map_x_47_data_org_near), .s_g(_add_map_x_47_s_g), .s_g_near(_add_map_x_47_s_g_near), .moto_org_near(_add_map_x_47_moto_org_near), .moto_org_near1(_add_map_x_47_moto_org_near1), .moto_org_near2(_add_map_x_47_moto_org_near2), .moto_org_near3(_add_map_x_47_moto_org_near3), .moto_org(_add_map_x_47_moto_org), .sg_up(_add_map_x_47_sg_up), .sg_down(_add_map_x_47_sg_down), .sg_left(_add_map_x_47_sg_left), .sg_right(_add_map_x_47_sg_right), .wall_t_in(_add_map_x_47_wall_t_in), .moto(_add_map_x_47_moto), .up(_add_map_x_47_up), .right(_add_map_x_47_right), .down(_add_map_x_47_down), .left(_add_map_x_47_left), .start(_add_map_x_47_start), .goal(_add_map_x_47_goal), .now(_add_map_x_47_now));
add_map add_map_x_46 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_46_add_exe), .data_out(_add_map_x_46_data_out), .data_out_index(_add_map_x_46_data_out_index), .data_near(_add_map_x_46_data_near), .wall_t_out(_add_map_x_46_wall_t_out), .data_org(_add_map_x_46_data_org), .data_org_near(_add_map_x_46_data_org_near), .s_g(_add_map_x_46_s_g), .s_g_near(_add_map_x_46_s_g_near), .moto_org_near(_add_map_x_46_moto_org_near), .moto_org_near1(_add_map_x_46_moto_org_near1), .moto_org_near2(_add_map_x_46_moto_org_near2), .moto_org_near3(_add_map_x_46_moto_org_near3), .moto_org(_add_map_x_46_moto_org), .sg_up(_add_map_x_46_sg_up), .sg_down(_add_map_x_46_sg_down), .sg_left(_add_map_x_46_sg_left), .sg_right(_add_map_x_46_sg_right), .wall_t_in(_add_map_x_46_wall_t_in), .moto(_add_map_x_46_moto), .up(_add_map_x_46_up), .right(_add_map_x_46_right), .down(_add_map_x_46_down), .left(_add_map_x_46_left), .start(_add_map_x_46_start), .goal(_add_map_x_46_goal), .now(_add_map_x_46_now));
add_map add_map_x_45 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_45_add_exe), .data_out(_add_map_x_45_data_out), .data_out_index(_add_map_x_45_data_out_index), .data_near(_add_map_x_45_data_near), .wall_t_out(_add_map_x_45_wall_t_out), .data_org(_add_map_x_45_data_org), .data_org_near(_add_map_x_45_data_org_near), .s_g(_add_map_x_45_s_g), .s_g_near(_add_map_x_45_s_g_near), .moto_org_near(_add_map_x_45_moto_org_near), .moto_org_near1(_add_map_x_45_moto_org_near1), .moto_org_near2(_add_map_x_45_moto_org_near2), .moto_org_near3(_add_map_x_45_moto_org_near3), .moto_org(_add_map_x_45_moto_org), .sg_up(_add_map_x_45_sg_up), .sg_down(_add_map_x_45_sg_down), .sg_left(_add_map_x_45_sg_left), .sg_right(_add_map_x_45_sg_right), .wall_t_in(_add_map_x_45_wall_t_in), .moto(_add_map_x_45_moto), .up(_add_map_x_45_up), .right(_add_map_x_45_right), .down(_add_map_x_45_down), .left(_add_map_x_45_left), .start(_add_map_x_45_start), .goal(_add_map_x_45_goal), .now(_add_map_x_45_now));
add_map add_map_x_44 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_44_add_exe), .data_out(_add_map_x_44_data_out), .data_out_index(_add_map_x_44_data_out_index), .data_near(_add_map_x_44_data_near), .wall_t_out(_add_map_x_44_wall_t_out), .data_org(_add_map_x_44_data_org), .data_org_near(_add_map_x_44_data_org_near), .s_g(_add_map_x_44_s_g), .s_g_near(_add_map_x_44_s_g_near), .moto_org_near(_add_map_x_44_moto_org_near), .moto_org_near1(_add_map_x_44_moto_org_near1), .moto_org_near2(_add_map_x_44_moto_org_near2), .moto_org_near3(_add_map_x_44_moto_org_near3), .moto_org(_add_map_x_44_moto_org), .sg_up(_add_map_x_44_sg_up), .sg_down(_add_map_x_44_sg_down), .sg_left(_add_map_x_44_sg_left), .sg_right(_add_map_x_44_sg_right), .wall_t_in(_add_map_x_44_wall_t_in), .moto(_add_map_x_44_moto), .up(_add_map_x_44_up), .right(_add_map_x_44_right), .down(_add_map_x_44_down), .left(_add_map_x_44_left), .start(_add_map_x_44_start), .goal(_add_map_x_44_goal), .now(_add_map_x_44_now));
add_map add_map_x_43 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_43_add_exe), .data_out(_add_map_x_43_data_out), .data_out_index(_add_map_x_43_data_out_index), .data_near(_add_map_x_43_data_near), .wall_t_out(_add_map_x_43_wall_t_out), .data_org(_add_map_x_43_data_org), .data_org_near(_add_map_x_43_data_org_near), .s_g(_add_map_x_43_s_g), .s_g_near(_add_map_x_43_s_g_near), .moto_org_near(_add_map_x_43_moto_org_near), .moto_org_near1(_add_map_x_43_moto_org_near1), .moto_org_near2(_add_map_x_43_moto_org_near2), .moto_org_near3(_add_map_x_43_moto_org_near3), .moto_org(_add_map_x_43_moto_org), .sg_up(_add_map_x_43_sg_up), .sg_down(_add_map_x_43_sg_down), .sg_left(_add_map_x_43_sg_left), .sg_right(_add_map_x_43_sg_right), .wall_t_in(_add_map_x_43_wall_t_in), .moto(_add_map_x_43_moto), .up(_add_map_x_43_up), .right(_add_map_x_43_right), .down(_add_map_x_43_down), .left(_add_map_x_43_left), .start(_add_map_x_43_start), .goal(_add_map_x_43_goal), .now(_add_map_x_43_now));
add_map add_map_x_42 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_42_add_exe), .data_out(_add_map_x_42_data_out), .data_out_index(_add_map_x_42_data_out_index), .data_near(_add_map_x_42_data_near), .wall_t_out(_add_map_x_42_wall_t_out), .data_org(_add_map_x_42_data_org), .data_org_near(_add_map_x_42_data_org_near), .s_g(_add_map_x_42_s_g), .s_g_near(_add_map_x_42_s_g_near), .moto_org_near(_add_map_x_42_moto_org_near), .moto_org_near1(_add_map_x_42_moto_org_near1), .moto_org_near2(_add_map_x_42_moto_org_near2), .moto_org_near3(_add_map_x_42_moto_org_near3), .moto_org(_add_map_x_42_moto_org), .sg_up(_add_map_x_42_sg_up), .sg_down(_add_map_x_42_sg_down), .sg_left(_add_map_x_42_sg_left), .sg_right(_add_map_x_42_sg_right), .wall_t_in(_add_map_x_42_wall_t_in), .moto(_add_map_x_42_moto), .up(_add_map_x_42_up), .right(_add_map_x_42_right), .down(_add_map_x_42_down), .left(_add_map_x_42_left), .start(_add_map_x_42_start), .goal(_add_map_x_42_goal), .now(_add_map_x_42_now));
add_map add_map_x_41 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_41_add_exe), .data_out(_add_map_x_41_data_out), .data_out_index(_add_map_x_41_data_out_index), .data_near(_add_map_x_41_data_near), .wall_t_out(_add_map_x_41_wall_t_out), .data_org(_add_map_x_41_data_org), .data_org_near(_add_map_x_41_data_org_near), .s_g(_add_map_x_41_s_g), .s_g_near(_add_map_x_41_s_g_near), .moto_org_near(_add_map_x_41_moto_org_near), .moto_org_near1(_add_map_x_41_moto_org_near1), .moto_org_near2(_add_map_x_41_moto_org_near2), .moto_org_near3(_add_map_x_41_moto_org_near3), .moto_org(_add_map_x_41_moto_org), .sg_up(_add_map_x_41_sg_up), .sg_down(_add_map_x_41_sg_down), .sg_left(_add_map_x_41_sg_left), .sg_right(_add_map_x_41_sg_right), .wall_t_in(_add_map_x_41_wall_t_in), .moto(_add_map_x_41_moto), .up(_add_map_x_41_up), .right(_add_map_x_41_right), .down(_add_map_x_41_down), .left(_add_map_x_41_left), .start(_add_map_x_41_start), .goal(_add_map_x_41_goal), .now(_add_map_x_41_now));
add_map add_map_x_40 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_40_add_exe), .data_out(_add_map_x_40_data_out), .data_out_index(_add_map_x_40_data_out_index), .data_near(_add_map_x_40_data_near), .wall_t_out(_add_map_x_40_wall_t_out), .data_org(_add_map_x_40_data_org), .data_org_near(_add_map_x_40_data_org_near), .s_g(_add_map_x_40_s_g), .s_g_near(_add_map_x_40_s_g_near), .moto_org_near(_add_map_x_40_moto_org_near), .moto_org_near1(_add_map_x_40_moto_org_near1), .moto_org_near2(_add_map_x_40_moto_org_near2), .moto_org_near3(_add_map_x_40_moto_org_near3), .moto_org(_add_map_x_40_moto_org), .sg_up(_add_map_x_40_sg_up), .sg_down(_add_map_x_40_sg_down), .sg_left(_add_map_x_40_sg_left), .sg_right(_add_map_x_40_sg_right), .wall_t_in(_add_map_x_40_wall_t_in), .moto(_add_map_x_40_moto), .up(_add_map_x_40_up), .right(_add_map_x_40_right), .down(_add_map_x_40_down), .left(_add_map_x_40_left), .start(_add_map_x_40_start), .goal(_add_map_x_40_goal), .now(_add_map_x_40_now));
add_map add_map_x_39 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_39_add_exe), .data_out(_add_map_x_39_data_out), .data_out_index(_add_map_x_39_data_out_index), .data_near(_add_map_x_39_data_near), .wall_t_out(_add_map_x_39_wall_t_out), .data_org(_add_map_x_39_data_org), .data_org_near(_add_map_x_39_data_org_near), .s_g(_add_map_x_39_s_g), .s_g_near(_add_map_x_39_s_g_near), .moto_org_near(_add_map_x_39_moto_org_near), .moto_org_near1(_add_map_x_39_moto_org_near1), .moto_org_near2(_add_map_x_39_moto_org_near2), .moto_org_near3(_add_map_x_39_moto_org_near3), .moto_org(_add_map_x_39_moto_org), .sg_up(_add_map_x_39_sg_up), .sg_down(_add_map_x_39_sg_down), .sg_left(_add_map_x_39_sg_left), .sg_right(_add_map_x_39_sg_right), .wall_t_in(_add_map_x_39_wall_t_in), .moto(_add_map_x_39_moto), .up(_add_map_x_39_up), .right(_add_map_x_39_right), .down(_add_map_x_39_down), .left(_add_map_x_39_left), .start(_add_map_x_39_start), .goal(_add_map_x_39_goal), .now(_add_map_x_39_now));
add_map add_map_x_38 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_38_add_exe), .data_out(_add_map_x_38_data_out), .data_out_index(_add_map_x_38_data_out_index), .data_near(_add_map_x_38_data_near), .wall_t_out(_add_map_x_38_wall_t_out), .data_org(_add_map_x_38_data_org), .data_org_near(_add_map_x_38_data_org_near), .s_g(_add_map_x_38_s_g), .s_g_near(_add_map_x_38_s_g_near), .moto_org_near(_add_map_x_38_moto_org_near), .moto_org_near1(_add_map_x_38_moto_org_near1), .moto_org_near2(_add_map_x_38_moto_org_near2), .moto_org_near3(_add_map_x_38_moto_org_near3), .moto_org(_add_map_x_38_moto_org), .sg_up(_add_map_x_38_sg_up), .sg_down(_add_map_x_38_sg_down), .sg_left(_add_map_x_38_sg_left), .sg_right(_add_map_x_38_sg_right), .wall_t_in(_add_map_x_38_wall_t_in), .moto(_add_map_x_38_moto), .up(_add_map_x_38_up), .right(_add_map_x_38_right), .down(_add_map_x_38_down), .left(_add_map_x_38_left), .start(_add_map_x_38_start), .goal(_add_map_x_38_goal), .now(_add_map_x_38_now));
add_map add_map_x_37 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_37_add_exe), .data_out(_add_map_x_37_data_out), .data_out_index(_add_map_x_37_data_out_index), .data_near(_add_map_x_37_data_near), .wall_t_out(_add_map_x_37_wall_t_out), .data_org(_add_map_x_37_data_org), .data_org_near(_add_map_x_37_data_org_near), .s_g(_add_map_x_37_s_g), .s_g_near(_add_map_x_37_s_g_near), .moto_org_near(_add_map_x_37_moto_org_near), .moto_org_near1(_add_map_x_37_moto_org_near1), .moto_org_near2(_add_map_x_37_moto_org_near2), .moto_org_near3(_add_map_x_37_moto_org_near3), .moto_org(_add_map_x_37_moto_org), .sg_up(_add_map_x_37_sg_up), .sg_down(_add_map_x_37_sg_down), .sg_left(_add_map_x_37_sg_left), .sg_right(_add_map_x_37_sg_right), .wall_t_in(_add_map_x_37_wall_t_in), .moto(_add_map_x_37_moto), .up(_add_map_x_37_up), .right(_add_map_x_37_right), .down(_add_map_x_37_down), .left(_add_map_x_37_left), .start(_add_map_x_37_start), .goal(_add_map_x_37_goal), .now(_add_map_x_37_now));
add_map add_map_x_36 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_36_add_exe), .data_out(_add_map_x_36_data_out), .data_out_index(_add_map_x_36_data_out_index), .data_near(_add_map_x_36_data_near), .wall_t_out(_add_map_x_36_wall_t_out), .data_org(_add_map_x_36_data_org), .data_org_near(_add_map_x_36_data_org_near), .s_g(_add_map_x_36_s_g), .s_g_near(_add_map_x_36_s_g_near), .moto_org_near(_add_map_x_36_moto_org_near), .moto_org_near1(_add_map_x_36_moto_org_near1), .moto_org_near2(_add_map_x_36_moto_org_near2), .moto_org_near3(_add_map_x_36_moto_org_near3), .moto_org(_add_map_x_36_moto_org), .sg_up(_add_map_x_36_sg_up), .sg_down(_add_map_x_36_sg_down), .sg_left(_add_map_x_36_sg_left), .sg_right(_add_map_x_36_sg_right), .wall_t_in(_add_map_x_36_wall_t_in), .moto(_add_map_x_36_moto), .up(_add_map_x_36_up), .right(_add_map_x_36_right), .down(_add_map_x_36_down), .left(_add_map_x_36_left), .start(_add_map_x_36_start), .goal(_add_map_x_36_goal), .now(_add_map_x_36_now));
add_map add_map_x_35 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_35_add_exe), .data_out(_add_map_x_35_data_out), .data_out_index(_add_map_x_35_data_out_index), .data_near(_add_map_x_35_data_near), .wall_t_out(_add_map_x_35_wall_t_out), .data_org(_add_map_x_35_data_org), .data_org_near(_add_map_x_35_data_org_near), .s_g(_add_map_x_35_s_g), .s_g_near(_add_map_x_35_s_g_near), .moto_org_near(_add_map_x_35_moto_org_near), .moto_org_near1(_add_map_x_35_moto_org_near1), .moto_org_near2(_add_map_x_35_moto_org_near2), .moto_org_near3(_add_map_x_35_moto_org_near3), .moto_org(_add_map_x_35_moto_org), .sg_up(_add_map_x_35_sg_up), .sg_down(_add_map_x_35_sg_down), .sg_left(_add_map_x_35_sg_left), .sg_right(_add_map_x_35_sg_right), .wall_t_in(_add_map_x_35_wall_t_in), .moto(_add_map_x_35_moto), .up(_add_map_x_35_up), .right(_add_map_x_35_right), .down(_add_map_x_35_down), .left(_add_map_x_35_left), .start(_add_map_x_35_start), .goal(_add_map_x_35_goal), .now(_add_map_x_35_now));
add_map add_map_x_34 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_34_add_exe), .data_out(_add_map_x_34_data_out), .data_out_index(_add_map_x_34_data_out_index), .data_near(_add_map_x_34_data_near), .wall_t_out(_add_map_x_34_wall_t_out), .data_org(_add_map_x_34_data_org), .data_org_near(_add_map_x_34_data_org_near), .s_g(_add_map_x_34_s_g), .s_g_near(_add_map_x_34_s_g_near), .moto_org_near(_add_map_x_34_moto_org_near), .moto_org_near1(_add_map_x_34_moto_org_near1), .moto_org_near2(_add_map_x_34_moto_org_near2), .moto_org_near3(_add_map_x_34_moto_org_near3), .moto_org(_add_map_x_34_moto_org), .sg_up(_add_map_x_34_sg_up), .sg_down(_add_map_x_34_sg_down), .sg_left(_add_map_x_34_sg_left), .sg_right(_add_map_x_34_sg_right), .wall_t_in(_add_map_x_34_wall_t_in), .moto(_add_map_x_34_moto), .up(_add_map_x_34_up), .right(_add_map_x_34_right), .down(_add_map_x_34_down), .left(_add_map_x_34_left), .start(_add_map_x_34_start), .goal(_add_map_x_34_goal), .now(_add_map_x_34_now));
add_map add_map_x_33 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_33_add_exe), .data_out(_add_map_x_33_data_out), .data_out_index(_add_map_x_33_data_out_index), .data_near(_add_map_x_33_data_near), .wall_t_out(_add_map_x_33_wall_t_out), .data_org(_add_map_x_33_data_org), .data_org_near(_add_map_x_33_data_org_near), .s_g(_add_map_x_33_s_g), .s_g_near(_add_map_x_33_s_g_near), .moto_org_near(_add_map_x_33_moto_org_near), .moto_org_near1(_add_map_x_33_moto_org_near1), .moto_org_near2(_add_map_x_33_moto_org_near2), .moto_org_near3(_add_map_x_33_moto_org_near3), .moto_org(_add_map_x_33_moto_org), .sg_up(_add_map_x_33_sg_up), .sg_down(_add_map_x_33_sg_down), .sg_left(_add_map_x_33_sg_left), .sg_right(_add_map_x_33_sg_right), .wall_t_in(_add_map_x_33_wall_t_in), .moto(_add_map_x_33_moto), .up(_add_map_x_33_up), .right(_add_map_x_33_right), .down(_add_map_x_33_down), .left(_add_map_x_33_left), .start(_add_map_x_33_start), .goal(_add_map_x_33_goal), .now(_add_map_x_33_now));
add_map add_map_x_32 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_32_add_exe), .data_out(_add_map_x_32_data_out), .data_out_index(_add_map_x_32_data_out_index), .data_near(_add_map_x_32_data_near), .wall_t_out(_add_map_x_32_wall_t_out), .data_org(_add_map_x_32_data_org), .data_org_near(_add_map_x_32_data_org_near), .s_g(_add_map_x_32_s_g), .s_g_near(_add_map_x_32_s_g_near), .moto_org_near(_add_map_x_32_moto_org_near), .moto_org_near1(_add_map_x_32_moto_org_near1), .moto_org_near2(_add_map_x_32_moto_org_near2), .moto_org_near3(_add_map_x_32_moto_org_near3), .moto_org(_add_map_x_32_moto_org), .sg_up(_add_map_x_32_sg_up), .sg_down(_add_map_x_32_sg_down), .sg_left(_add_map_x_32_sg_left), .sg_right(_add_map_x_32_sg_right), .wall_t_in(_add_map_x_32_wall_t_in), .moto(_add_map_x_32_moto), .up(_add_map_x_32_up), .right(_add_map_x_32_right), .down(_add_map_x_32_down), .left(_add_map_x_32_left), .start(_add_map_x_32_start), .goal(_add_map_x_32_goal), .now(_add_map_x_32_now));
add_map add_map_x_31 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_31_add_exe), .data_out(_add_map_x_31_data_out), .data_out_index(_add_map_x_31_data_out_index), .data_near(_add_map_x_31_data_near), .wall_t_out(_add_map_x_31_wall_t_out), .data_org(_add_map_x_31_data_org), .data_org_near(_add_map_x_31_data_org_near), .s_g(_add_map_x_31_s_g), .s_g_near(_add_map_x_31_s_g_near), .moto_org_near(_add_map_x_31_moto_org_near), .moto_org_near1(_add_map_x_31_moto_org_near1), .moto_org_near2(_add_map_x_31_moto_org_near2), .moto_org_near3(_add_map_x_31_moto_org_near3), .moto_org(_add_map_x_31_moto_org), .sg_up(_add_map_x_31_sg_up), .sg_down(_add_map_x_31_sg_down), .sg_left(_add_map_x_31_sg_left), .sg_right(_add_map_x_31_sg_right), .wall_t_in(_add_map_x_31_wall_t_in), .moto(_add_map_x_31_moto), .up(_add_map_x_31_up), .right(_add_map_x_31_right), .down(_add_map_x_31_down), .left(_add_map_x_31_left), .start(_add_map_x_31_start), .goal(_add_map_x_31_goal), .now(_add_map_x_31_now));
add_map add_map_x_30 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_30_add_exe), .data_out(_add_map_x_30_data_out), .data_out_index(_add_map_x_30_data_out_index), .data_near(_add_map_x_30_data_near), .wall_t_out(_add_map_x_30_wall_t_out), .data_org(_add_map_x_30_data_org), .data_org_near(_add_map_x_30_data_org_near), .s_g(_add_map_x_30_s_g), .s_g_near(_add_map_x_30_s_g_near), .moto_org_near(_add_map_x_30_moto_org_near), .moto_org_near1(_add_map_x_30_moto_org_near1), .moto_org_near2(_add_map_x_30_moto_org_near2), .moto_org_near3(_add_map_x_30_moto_org_near3), .moto_org(_add_map_x_30_moto_org), .sg_up(_add_map_x_30_sg_up), .sg_down(_add_map_x_30_sg_down), .sg_left(_add_map_x_30_sg_left), .sg_right(_add_map_x_30_sg_right), .wall_t_in(_add_map_x_30_wall_t_in), .moto(_add_map_x_30_moto), .up(_add_map_x_30_up), .right(_add_map_x_30_right), .down(_add_map_x_30_down), .left(_add_map_x_30_left), .start(_add_map_x_30_start), .goal(_add_map_x_30_goal), .now(_add_map_x_30_now));
add_map add_map_x_29 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_29_add_exe), .data_out(_add_map_x_29_data_out), .data_out_index(_add_map_x_29_data_out_index), .data_near(_add_map_x_29_data_near), .wall_t_out(_add_map_x_29_wall_t_out), .data_org(_add_map_x_29_data_org), .data_org_near(_add_map_x_29_data_org_near), .s_g(_add_map_x_29_s_g), .s_g_near(_add_map_x_29_s_g_near), .moto_org_near(_add_map_x_29_moto_org_near), .moto_org_near1(_add_map_x_29_moto_org_near1), .moto_org_near2(_add_map_x_29_moto_org_near2), .moto_org_near3(_add_map_x_29_moto_org_near3), .moto_org(_add_map_x_29_moto_org), .sg_up(_add_map_x_29_sg_up), .sg_down(_add_map_x_29_sg_down), .sg_left(_add_map_x_29_sg_left), .sg_right(_add_map_x_29_sg_right), .wall_t_in(_add_map_x_29_wall_t_in), .moto(_add_map_x_29_moto), .up(_add_map_x_29_up), .right(_add_map_x_29_right), .down(_add_map_x_29_down), .left(_add_map_x_29_left), .start(_add_map_x_29_start), .goal(_add_map_x_29_goal), .now(_add_map_x_29_now));
add_map add_map_x_28 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_28_add_exe), .data_out(_add_map_x_28_data_out), .data_out_index(_add_map_x_28_data_out_index), .data_near(_add_map_x_28_data_near), .wall_t_out(_add_map_x_28_wall_t_out), .data_org(_add_map_x_28_data_org), .data_org_near(_add_map_x_28_data_org_near), .s_g(_add_map_x_28_s_g), .s_g_near(_add_map_x_28_s_g_near), .moto_org_near(_add_map_x_28_moto_org_near), .moto_org_near1(_add_map_x_28_moto_org_near1), .moto_org_near2(_add_map_x_28_moto_org_near2), .moto_org_near3(_add_map_x_28_moto_org_near3), .moto_org(_add_map_x_28_moto_org), .sg_up(_add_map_x_28_sg_up), .sg_down(_add_map_x_28_sg_down), .sg_left(_add_map_x_28_sg_left), .sg_right(_add_map_x_28_sg_right), .wall_t_in(_add_map_x_28_wall_t_in), .moto(_add_map_x_28_moto), .up(_add_map_x_28_up), .right(_add_map_x_28_right), .down(_add_map_x_28_down), .left(_add_map_x_28_left), .start(_add_map_x_28_start), .goal(_add_map_x_28_goal), .now(_add_map_x_28_now));
add_map add_map_x_27 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_27_add_exe), .data_out(_add_map_x_27_data_out), .data_out_index(_add_map_x_27_data_out_index), .data_near(_add_map_x_27_data_near), .wall_t_out(_add_map_x_27_wall_t_out), .data_org(_add_map_x_27_data_org), .data_org_near(_add_map_x_27_data_org_near), .s_g(_add_map_x_27_s_g), .s_g_near(_add_map_x_27_s_g_near), .moto_org_near(_add_map_x_27_moto_org_near), .moto_org_near1(_add_map_x_27_moto_org_near1), .moto_org_near2(_add_map_x_27_moto_org_near2), .moto_org_near3(_add_map_x_27_moto_org_near3), .moto_org(_add_map_x_27_moto_org), .sg_up(_add_map_x_27_sg_up), .sg_down(_add_map_x_27_sg_down), .sg_left(_add_map_x_27_sg_left), .sg_right(_add_map_x_27_sg_right), .wall_t_in(_add_map_x_27_wall_t_in), .moto(_add_map_x_27_moto), .up(_add_map_x_27_up), .right(_add_map_x_27_right), .down(_add_map_x_27_down), .left(_add_map_x_27_left), .start(_add_map_x_27_start), .goal(_add_map_x_27_goal), .now(_add_map_x_27_now));
add_map add_map_x_26 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_26_add_exe), .data_out(_add_map_x_26_data_out), .data_out_index(_add_map_x_26_data_out_index), .data_near(_add_map_x_26_data_near), .wall_t_out(_add_map_x_26_wall_t_out), .data_org(_add_map_x_26_data_org), .data_org_near(_add_map_x_26_data_org_near), .s_g(_add_map_x_26_s_g), .s_g_near(_add_map_x_26_s_g_near), .moto_org_near(_add_map_x_26_moto_org_near), .moto_org_near1(_add_map_x_26_moto_org_near1), .moto_org_near2(_add_map_x_26_moto_org_near2), .moto_org_near3(_add_map_x_26_moto_org_near3), .moto_org(_add_map_x_26_moto_org), .sg_up(_add_map_x_26_sg_up), .sg_down(_add_map_x_26_sg_down), .sg_left(_add_map_x_26_sg_left), .sg_right(_add_map_x_26_sg_right), .wall_t_in(_add_map_x_26_wall_t_in), .moto(_add_map_x_26_moto), .up(_add_map_x_26_up), .right(_add_map_x_26_right), .down(_add_map_x_26_down), .left(_add_map_x_26_left), .start(_add_map_x_26_start), .goal(_add_map_x_26_goal), .now(_add_map_x_26_now));
add_map add_map_x_25 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_25_add_exe), .data_out(_add_map_x_25_data_out), .data_out_index(_add_map_x_25_data_out_index), .data_near(_add_map_x_25_data_near), .wall_t_out(_add_map_x_25_wall_t_out), .data_org(_add_map_x_25_data_org), .data_org_near(_add_map_x_25_data_org_near), .s_g(_add_map_x_25_s_g), .s_g_near(_add_map_x_25_s_g_near), .moto_org_near(_add_map_x_25_moto_org_near), .moto_org_near1(_add_map_x_25_moto_org_near1), .moto_org_near2(_add_map_x_25_moto_org_near2), .moto_org_near3(_add_map_x_25_moto_org_near3), .moto_org(_add_map_x_25_moto_org), .sg_up(_add_map_x_25_sg_up), .sg_down(_add_map_x_25_sg_down), .sg_left(_add_map_x_25_sg_left), .sg_right(_add_map_x_25_sg_right), .wall_t_in(_add_map_x_25_wall_t_in), .moto(_add_map_x_25_moto), .up(_add_map_x_25_up), .right(_add_map_x_25_right), .down(_add_map_x_25_down), .left(_add_map_x_25_left), .start(_add_map_x_25_start), .goal(_add_map_x_25_goal), .now(_add_map_x_25_now));
add_map add_map_x_24 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_24_add_exe), .data_out(_add_map_x_24_data_out), .data_out_index(_add_map_x_24_data_out_index), .data_near(_add_map_x_24_data_near), .wall_t_out(_add_map_x_24_wall_t_out), .data_org(_add_map_x_24_data_org), .data_org_near(_add_map_x_24_data_org_near), .s_g(_add_map_x_24_s_g), .s_g_near(_add_map_x_24_s_g_near), .moto_org_near(_add_map_x_24_moto_org_near), .moto_org_near1(_add_map_x_24_moto_org_near1), .moto_org_near2(_add_map_x_24_moto_org_near2), .moto_org_near3(_add_map_x_24_moto_org_near3), .moto_org(_add_map_x_24_moto_org), .sg_up(_add_map_x_24_sg_up), .sg_down(_add_map_x_24_sg_down), .sg_left(_add_map_x_24_sg_left), .sg_right(_add_map_x_24_sg_right), .wall_t_in(_add_map_x_24_wall_t_in), .moto(_add_map_x_24_moto), .up(_add_map_x_24_up), .right(_add_map_x_24_right), .down(_add_map_x_24_down), .left(_add_map_x_24_left), .start(_add_map_x_24_start), .goal(_add_map_x_24_goal), .now(_add_map_x_24_now));
add_map add_map_x_23 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_23_add_exe), .data_out(_add_map_x_23_data_out), .data_out_index(_add_map_x_23_data_out_index), .data_near(_add_map_x_23_data_near), .wall_t_out(_add_map_x_23_wall_t_out), .data_org(_add_map_x_23_data_org), .data_org_near(_add_map_x_23_data_org_near), .s_g(_add_map_x_23_s_g), .s_g_near(_add_map_x_23_s_g_near), .moto_org_near(_add_map_x_23_moto_org_near), .moto_org_near1(_add_map_x_23_moto_org_near1), .moto_org_near2(_add_map_x_23_moto_org_near2), .moto_org_near3(_add_map_x_23_moto_org_near3), .moto_org(_add_map_x_23_moto_org), .sg_up(_add_map_x_23_sg_up), .sg_down(_add_map_x_23_sg_down), .sg_left(_add_map_x_23_sg_left), .sg_right(_add_map_x_23_sg_right), .wall_t_in(_add_map_x_23_wall_t_in), .moto(_add_map_x_23_moto), .up(_add_map_x_23_up), .right(_add_map_x_23_right), .down(_add_map_x_23_down), .left(_add_map_x_23_left), .start(_add_map_x_23_start), .goal(_add_map_x_23_goal), .now(_add_map_x_23_now));
add_map add_map_x_22 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_22_add_exe), .data_out(_add_map_x_22_data_out), .data_out_index(_add_map_x_22_data_out_index), .data_near(_add_map_x_22_data_near), .wall_t_out(_add_map_x_22_wall_t_out), .data_org(_add_map_x_22_data_org), .data_org_near(_add_map_x_22_data_org_near), .s_g(_add_map_x_22_s_g), .s_g_near(_add_map_x_22_s_g_near), .moto_org_near(_add_map_x_22_moto_org_near), .moto_org_near1(_add_map_x_22_moto_org_near1), .moto_org_near2(_add_map_x_22_moto_org_near2), .moto_org_near3(_add_map_x_22_moto_org_near3), .moto_org(_add_map_x_22_moto_org), .sg_up(_add_map_x_22_sg_up), .sg_down(_add_map_x_22_sg_down), .sg_left(_add_map_x_22_sg_left), .sg_right(_add_map_x_22_sg_right), .wall_t_in(_add_map_x_22_wall_t_in), .moto(_add_map_x_22_moto), .up(_add_map_x_22_up), .right(_add_map_x_22_right), .down(_add_map_x_22_down), .left(_add_map_x_22_left), .start(_add_map_x_22_start), .goal(_add_map_x_22_goal), .now(_add_map_x_22_now));
add_map add_map_x_21 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_21_add_exe), .data_out(_add_map_x_21_data_out), .data_out_index(_add_map_x_21_data_out_index), .data_near(_add_map_x_21_data_near), .wall_t_out(_add_map_x_21_wall_t_out), .data_org(_add_map_x_21_data_org), .data_org_near(_add_map_x_21_data_org_near), .s_g(_add_map_x_21_s_g), .s_g_near(_add_map_x_21_s_g_near), .moto_org_near(_add_map_x_21_moto_org_near), .moto_org_near1(_add_map_x_21_moto_org_near1), .moto_org_near2(_add_map_x_21_moto_org_near2), .moto_org_near3(_add_map_x_21_moto_org_near3), .moto_org(_add_map_x_21_moto_org), .sg_up(_add_map_x_21_sg_up), .sg_down(_add_map_x_21_sg_down), .sg_left(_add_map_x_21_sg_left), .sg_right(_add_map_x_21_sg_right), .wall_t_in(_add_map_x_21_wall_t_in), .moto(_add_map_x_21_moto), .up(_add_map_x_21_up), .right(_add_map_x_21_right), .down(_add_map_x_21_down), .left(_add_map_x_21_left), .start(_add_map_x_21_start), .goal(_add_map_x_21_goal), .now(_add_map_x_21_now));
add_map add_map_x_20 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_20_add_exe), .data_out(_add_map_x_20_data_out), .data_out_index(_add_map_x_20_data_out_index), .data_near(_add_map_x_20_data_near), .wall_t_out(_add_map_x_20_wall_t_out), .data_org(_add_map_x_20_data_org), .data_org_near(_add_map_x_20_data_org_near), .s_g(_add_map_x_20_s_g), .s_g_near(_add_map_x_20_s_g_near), .moto_org_near(_add_map_x_20_moto_org_near), .moto_org_near1(_add_map_x_20_moto_org_near1), .moto_org_near2(_add_map_x_20_moto_org_near2), .moto_org_near3(_add_map_x_20_moto_org_near3), .moto_org(_add_map_x_20_moto_org), .sg_up(_add_map_x_20_sg_up), .sg_down(_add_map_x_20_sg_down), .sg_left(_add_map_x_20_sg_left), .sg_right(_add_map_x_20_sg_right), .wall_t_in(_add_map_x_20_wall_t_in), .moto(_add_map_x_20_moto), .up(_add_map_x_20_up), .right(_add_map_x_20_right), .down(_add_map_x_20_down), .left(_add_map_x_20_left), .start(_add_map_x_20_start), .goal(_add_map_x_20_goal), .now(_add_map_x_20_now));
add_map add_map_x_19 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_19_add_exe), .data_out(_add_map_x_19_data_out), .data_out_index(_add_map_x_19_data_out_index), .data_near(_add_map_x_19_data_near), .wall_t_out(_add_map_x_19_wall_t_out), .data_org(_add_map_x_19_data_org), .data_org_near(_add_map_x_19_data_org_near), .s_g(_add_map_x_19_s_g), .s_g_near(_add_map_x_19_s_g_near), .moto_org_near(_add_map_x_19_moto_org_near), .moto_org_near1(_add_map_x_19_moto_org_near1), .moto_org_near2(_add_map_x_19_moto_org_near2), .moto_org_near3(_add_map_x_19_moto_org_near3), .moto_org(_add_map_x_19_moto_org), .sg_up(_add_map_x_19_sg_up), .sg_down(_add_map_x_19_sg_down), .sg_left(_add_map_x_19_sg_left), .sg_right(_add_map_x_19_sg_right), .wall_t_in(_add_map_x_19_wall_t_in), .moto(_add_map_x_19_moto), .up(_add_map_x_19_up), .right(_add_map_x_19_right), .down(_add_map_x_19_down), .left(_add_map_x_19_left), .start(_add_map_x_19_start), .goal(_add_map_x_19_goal), .now(_add_map_x_19_now));
add_map add_map_x_18 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_18_add_exe), .data_out(_add_map_x_18_data_out), .data_out_index(_add_map_x_18_data_out_index), .data_near(_add_map_x_18_data_near), .wall_t_out(_add_map_x_18_wall_t_out), .data_org(_add_map_x_18_data_org), .data_org_near(_add_map_x_18_data_org_near), .s_g(_add_map_x_18_s_g), .s_g_near(_add_map_x_18_s_g_near), .moto_org_near(_add_map_x_18_moto_org_near), .moto_org_near1(_add_map_x_18_moto_org_near1), .moto_org_near2(_add_map_x_18_moto_org_near2), .moto_org_near3(_add_map_x_18_moto_org_near3), .moto_org(_add_map_x_18_moto_org), .sg_up(_add_map_x_18_sg_up), .sg_down(_add_map_x_18_sg_down), .sg_left(_add_map_x_18_sg_left), .sg_right(_add_map_x_18_sg_right), .wall_t_in(_add_map_x_18_wall_t_in), .moto(_add_map_x_18_moto), .up(_add_map_x_18_up), .right(_add_map_x_18_right), .down(_add_map_x_18_down), .left(_add_map_x_18_left), .start(_add_map_x_18_start), .goal(_add_map_x_18_goal), .now(_add_map_x_18_now));
add_map add_map_x_17 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_17_add_exe), .data_out(_add_map_x_17_data_out), .data_out_index(_add_map_x_17_data_out_index), .data_near(_add_map_x_17_data_near), .wall_t_out(_add_map_x_17_wall_t_out), .data_org(_add_map_x_17_data_org), .data_org_near(_add_map_x_17_data_org_near), .s_g(_add_map_x_17_s_g), .s_g_near(_add_map_x_17_s_g_near), .moto_org_near(_add_map_x_17_moto_org_near), .moto_org_near1(_add_map_x_17_moto_org_near1), .moto_org_near2(_add_map_x_17_moto_org_near2), .moto_org_near3(_add_map_x_17_moto_org_near3), .moto_org(_add_map_x_17_moto_org), .sg_up(_add_map_x_17_sg_up), .sg_down(_add_map_x_17_sg_down), .sg_left(_add_map_x_17_sg_left), .sg_right(_add_map_x_17_sg_right), .wall_t_in(_add_map_x_17_wall_t_in), .moto(_add_map_x_17_moto), .up(_add_map_x_17_up), .right(_add_map_x_17_right), .down(_add_map_x_17_down), .left(_add_map_x_17_left), .start(_add_map_x_17_start), .goal(_add_map_x_17_goal), .now(_add_map_x_17_now));
add_map add_map_x_16 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_16_add_exe), .data_out(_add_map_x_16_data_out), .data_out_index(_add_map_x_16_data_out_index), .data_near(_add_map_x_16_data_near), .wall_t_out(_add_map_x_16_wall_t_out), .data_org(_add_map_x_16_data_org), .data_org_near(_add_map_x_16_data_org_near), .s_g(_add_map_x_16_s_g), .s_g_near(_add_map_x_16_s_g_near), .moto_org_near(_add_map_x_16_moto_org_near), .moto_org_near1(_add_map_x_16_moto_org_near1), .moto_org_near2(_add_map_x_16_moto_org_near2), .moto_org_near3(_add_map_x_16_moto_org_near3), .moto_org(_add_map_x_16_moto_org), .sg_up(_add_map_x_16_sg_up), .sg_down(_add_map_x_16_sg_down), .sg_left(_add_map_x_16_sg_left), .sg_right(_add_map_x_16_sg_right), .wall_t_in(_add_map_x_16_wall_t_in), .moto(_add_map_x_16_moto), .up(_add_map_x_16_up), .right(_add_map_x_16_right), .down(_add_map_x_16_down), .left(_add_map_x_16_left), .start(_add_map_x_16_start), .goal(_add_map_x_16_goal), .now(_add_map_x_16_now));
add_map add_map_x_15 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_15_add_exe), .data_out(_add_map_x_15_data_out), .data_out_index(_add_map_x_15_data_out_index), .data_near(_add_map_x_15_data_near), .wall_t_out(_add_map_x_15_wall_t_out), .data_org(_add_map_x_15_data_org), .data_org_near(_add_map_x_15_data_org_near), .s_g(_add_map_x_15_s_g), .s_g_near(_add_map_x_15_s_g_near), .moto_org_near(_add_map_x_15_moto_org_near), .moto_org_near1(_add_map_x_15_moto_org_near1), .moto_org_near2(_add_map_x_15_moto_org_near2), .moto_org_near3(_add_map_x_15_moto_org_near3), .moto_org(_add_map_x_15_moto_org), .sg_up(_add_map_x_15_sg_up), .sg_down(_add_map_x_15_sg_down), .sg_left(_add_map_x_15_sg_left), .sg_right(_add_map_x_15_sg_right), .wall_t_in(_add_map_x_15_wall_t_in), .moto(_add_map_x_15_moto), .up(_add_map_x_15_up), .right(_add_map_x_15_right), .down(_add_map_x_15_down), .left(_add_map_x_15_left), .start(_add_map_x_15_start), .goal(_add_map_x_15_goal), .now(_add_map_x_15_now));
add_map add_map_x_14 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_14_add_exe), .data_out(_add_map_x_14_data_out), .data_out_index(_add_map_x_14_data_out_index), .data_near(_add_map_x_14_data_near), .wall_t_out(_add_map_x_14_wall_t_out), .data_org(_add_map_x_14_data_org), .data_org_near(_add_map_x_14_data_org_near), .s_g(_add_map_x_14_s_g), .s_g_near(_add_map_x_14_s_g_near), .moto_org_near(_add_map_x_14_moto_org_near), .moto_org_near1(_add_map_x_14_moto_org_near1), .moto_org_near2(_add_map_x_14_moto_org_near2), .moto_org_near3(_add_map_x_14_moto_org_near3), .moto_org(_add_map_x_14_moto_org), .sg_up(_add_map_x_14_sg_up), .sg_down(_add_map_x_14_sg_down), .sg_left(_add_map_x_14_sg_left), .sg_right(_add_map_x_14_sg_right), .wall_t_in(_add_map_x_14_wall_t_in), .moto(_add_map_x_14_moto), .up(_add_map_x_14_up), .right(_add_map_x_14_right), .down(_add_map_x_14_down), .left(_add_map_x_14_left), .start(_add_map_x_14_start), .goal(_add_map_x_14_goal), .now(_add_map_x_14_now));
add_map add_map_x_13 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_13_add_exe), .data_out(_add_map_x_13_data_out), .data_out_index(_add_map_x_13_data_out_index), .data_near(_add_map_x_13_data_near), .wall_t_out(_add_map_x_13_wall_t_out), .data_org(_add_map_x_13_data_org), .data_org_near(_add_map_x_13_data_org_near), .s_g(_add_map_x_13_s_g), .s_g_near(_add_map_x_13_s_g_near), .moto_org_near(_add_map_x_13_moto_org_near), .moto_org_near1(_add_map_x_13_moto_org_near1), .moto_org_near2(_add_map_x_13_moto_org_near2), .moto_org_near3(_add_map_x_13_moto_org_near3), .moto_org(_add_map_x_13_moto_org), .sg_up(_add_map_x_13_sg_up), .sg_down(_add_map_x_13_sg_down), .sg_left(_add_map_x_13_sg_left), .sg_right(_add_map_x_13_sg_right), .wall_t_in(_add_map_x_13_wall_t_in), .moto(_add_map_x_13_moto), .up(_add_map_x_13_up), .right(_add_map_x_13_right), .down(_add_map_x_13_down), .left(_add_map_x_13_left), .start(_add_map_x_13_start), .goal(_add_map_x_13_goal), .now(_add_map_x_13_now));
add_map add_map_x_12 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_12_add_exe), .data_out(_add_map_x_12_data_out), .data_out_index(_add_map_x_12_data_out_index), .data_near(_add_map_x_12_data_near), .wall_t_out(_add_map_x_12_wall_t_out), .data_org(_add_map_x_12_data_org), .data_org_near(_add_map_x_12_data_org_near), .s_g(_add_map_x_12_s_g), .s_g_near(_add_map_x_12_s_g_near), .moto_org_near(_add_map_x_12_moto_org_near), .moto_org_near1(_add_map_x_12_moto_org_near1), .moto_org_near2(_add_map_x_12_moto_org_near2), .moto_org_near3(_add_map_x_12_moto_org_near3), .moto_org(_add_map_x_12_moto_org), .sg_up(_add_map_x_12_sg_up), .sg_down(_add_map_x_12_sg_down), .sg_left(_add_map_x_12_sg_left), .sg_right(_add_map_x_12_sg_right), .wall_t_in(_add_map_x_12_wall_t_in), .moto(_add_map_x_12_moto), .up(_add_map_x_12_up), .right(_add_map_x_12_right), .down(_add_map_x_12_down), .left(_add_map_x_12_left), .start(_add_map_x_12_start), .goal(_add_map_x_12_goal), .now(_add_map_x_12_now));
add_map add_map_x_11 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_11_add_exe), .data_out(_add_map_x_11_data_out), .data_out_index(_add_map_x_11_data_out_index), .data_near(_add_map_x_11_data_near), .wall_t_out(_add_map_x_11_wall_t_out), .data_org(_add_map_x_11_data_org), .data_org_near(_add_map_x_11_data_org_near), .s_g(_add_map_x_11_s_g), .s_g_near(_add_map_x_11_s_g_near), .moto_org_near(_add_map_x_11_moto_org_near), .moto_org_near1(_add_map_x_11_moto_org_near1), .moto_org_near2(_add_map_x_11_moto_org_near2), .moto_org_near3(_add_map_x_11_moto_org_near3), .moto_org(_add_map_x_11_moto_org), .sg_up(_add_map_x_11_sg_up), .sg_down(_add_map_x_11_sg_down), .sg_left(_add_map_x_11_sg_left), .sg_right(_add_map_x_11_sg_right), .wall_t_in(_add_map_x_11_wall_t_in), .moto(_add_map_x_11_moto), .up(_add_map_x_11_up), .right(_add_map_x_11_right), .down(_add_map_x_11_down), .left(_add_map_x_11_left), .start(_add_map_x_11_start), .goal(_add_map_x_11_goal), .now(_add_map_x_11_now));
add_map add_map_x_10 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_10_add_exe), .data_out(_add_map_x_10_data_out), .data_out_index(_add_map_x_10_data_out_index), .data_near(_add_map_x_10_data_near), .wall_t_out(_add_map_x_10_wall_t_out), .data_org(_add_map_x_10_data_org), .data_org_near(_add_map_x_10_data_org_near), .s_g(_add_map_x_10_s_g), .s_g_near(_add_map_x_10_s_g_near), .moto_org_near(_add_map_x_10_moto_org_near), .moto_org_near1(_add_map_x_10_moto_org_near1), .moto_org_near2(_add_map_x_10_moto_org_near2), .moto_org_near3(_add_map_x_10_moto_org_near3), .moto_org(_add_map_x_10_moto_org), .sg_up(_add_map_x_10_sg_up), .sg_down(_add_map_x_10_sg_down), .sg_left(_add_map_x_10_sg_left), .sg_right(_add_map_x_10_sg_right), .wall_t_in(_add_map_x_10_wall_t_in), .moto(_add_map_x_10_moto), .up(_add_map_x_10_up), .right(_add_map_x_10_right), .down(_add_map_x_10_down), .left(_add_map_x_10_left), .start(_add_map_x_10_start), .goal(_add_map_x_10_goal), .now(_add_map_x_10_now));
add_map add_map_x_9 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_9_add_exe), .data_out(_add_map_x_9_data_out), .data_out_index(_add_map_x_9_data_out_index), .data_near(_add_map_x_9_data_near), .wall_t_out(_add_map_x_9_wall_t_out), .data_org(_add_map_x_9_data_org), .data_org_near(_add_map_x_9_data_org_near), .s_g(_add_map_x_9_s_g), .s_g_near(_add_map_x_9_s_g_near), .moto_org_near(_add_map_x_9_moto_org_near), .moto_org_near1(_add_map_x_9_moto_org_near1), .moto_org_near2(_add_map_x_9_moto_org_near2), .moto_org_near3(_add_map_x_9_moto_org_near3), .moto_org(_add_map_x_9_moto_org), .sg_up(_add_map_x_9_sg_up), .sg_down(_add_map_x_9_sg_down), .sg_left(_add_map_x_9_sg_left), .sg_right(_add_map_x_9_sg_right), .wall_t_in(_add_map_x_9_wall_t_in), .moto(_add_map_x_9_moto), .up(_add_map_x_9_up), .right(_add_map_x_9_right), .down(_add_map_x_9_down), .left(_add_map_x_9_left), .start(_add_map_x_9_start), .goal(_add_map_x_9_goal), .now(_add_map_x_9_now));
add_map add_map_x_8 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_8_add_exe), .data_out(_add_map_x_8_data_out), .data_out_index(_add_map_x_8_data_out_index), .data_near(_add_map_x_8_data_near), .wall_t_out(_add_map_x_8_wall_t_out), .data_org(_add_map_x_8_data_org), .data_org_near(_add_map_x_8_data_org_near), .s_g(_add_map_x_8_s_g), .s_g_near(_add_map_x_8_s_g_near), .moto_org_near(_add_map_x_8_moto_org_near), .moto_org_near1(_add_map_x_8_moto_org_near1), .moto_org_near2(_add_map_x_8_moto_org_near2), .moto_org_near3(_add_map_x_8_moto_org_near3), .moto_org(_add_map_x_8_moto_org), .sg_up(_add_map_x_8_sg_up), .sg_down(_add_map_x_8_sg_down), .sg_left(_add_map_x_8_sg_left), .sg_right(_add_map_x_8_sg_right), .wall_t_in(_add_map_x_8_wall_t_in), .moto(_add_map_x_8_moto), .up(_add_map_x_8_up), .right(_add_map_x_8_right), .down(_add_map_x_8_down), .left(_add_map_x_8_left), .start(_add_map_x_8_start), .goal(_add_map_x_8_goal), .now(_add_map_x_8_now));
add_map add_map_x_7 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_7_add_exe), .data_out(_add_map_x_7_data_out), .data_out_index(_add_map_x_7_data_out_index), .data_near(_add_map_x_7_data_near), .wall_t_out(_add_map_x_7_wall_t_out), .data_org(_add_map_x_7_data_org), .data_org_near(_add_map_x_7_data_org_near), .s_g(_add_map_x_7_s_g), .s_g_near(_add_map_x_7_s_g_near), .moto_org_near(_add_map_x_7_moto_org_near), .moto_org_near1(_add_map_x_7_moto_org_near1), .moto_org_near2(_add_map_x_7_moto_org_near2), .moto_org_near3(_add_map_x_7_moto_org_near3), .moto_org(_add_map_x_7_moto_org), .sg_up(_add_map_x_7_sg_up), .sg_down(_add_map_x_7_sg_down), .sg_left(_add_map_x_7_sg_left), .sg_right(_add_map_x_7_sg_right), .wall_t_in(_add_map_x_7_wall_t_in), .moto(_add_map_x_7_moto), .up(_add_map_x_7_up), .right(_add_map_x_7_right), .down(_add_map_x_7_down), .left(_add_map_x_7_left), .start(_add_map_x_7_start), .goal(_add_map_x_7_goal), .now(_add_map_x_7_now));
add_map add_map_x_6 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_6_add_exe), .data_out(_add_map_x_6_data_out), .data_out_index(_add_map_x_6_data_out_index), .data_near(_add_map_x_6_data_near), .wall_t_out(_add_map_x_6_wall_t_out), .data_org(_add_map_x_6_data_org), .data_org_near(_add_map_x_6_data_org_near), .s_g(_add_map_x_6_s_g), .s_g_near(_add_map_x_6_s_g_near), .moto_org_near(_add_map_x_6_moto_org_near), .moto_org_near1(_add_map_x_6_moto_org_near1), .moto_org_near2(_add_map_x_6_moto_org_near2), .moto_org_near3(_add_map_x_6_moto_org_near3), .moto_org(_add_map_x_6_moto_org), .sg_up(_add_map_x_6_sg_up), .sg_down(_add_map_x_6_sg_down), .sg_left(_add_map_x_6_sg_left), .sg_right(_add_map_x_6_sg_right), .wall_t_in(_add_map_x_6_wall_t_in), .moto(_add_map_x_6_moto), .up(_add_map_x_6_up), .right(_add_map_x_6_right), .down(_add_map_x_6_down), .left(_add_map_x_6_left), .start(_add_map_x_6_start), .goal(_add_map_x_6_goal), .now(_add_map_x_6_now));
add_map add_map_x_5 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_5_add_exe), .data_out(_add_map_x_5_data_out), .data_out_index(_add_map_x_5_data_out_index), .data_near(_add_map_x_5_data_near), .wall_t_out(_add_map_x_5_wall_t_out), .data_org(_add_map_x_5_data_org), .data_org_near(_add_map_x_5_data_org_near), .s_g(_add_map_x_5_s_g), .s_g_near(_add_map_x_5_s_g_near), .moto_org_near(_add_map_x_5_moto_org_near), .moto_org_near1(_add_map_x_5_moto_org_near1), .moto_org_near2(_add_map_x_5_moto_org_near2), .moto_org_near3(_add_map_x_5_moto_org_near3), .moto_org(_add_map_x_5_moto_org), .sg_up(_add_map_x_5_sg_up), .sg_down(_add_map_x_5_sg_down), .sg_left(_add_map_x_5_sg_left), .sg_right(_add_map_x_5_sg_right), .wall_t_in(_add_map_x_5_wall_t_in), .moto(_add_map_x_5_moto), .up(_add_map_x_5_up), .right(_add_map_x_5_right), .down(_add_map_x_5_down), .left(_add_map_x_5_left), .start(_add_map_x_5_start), .goal(_add_map_x_5_goal), .now(_add_map_x_5_now));
add_map add_map_x_4 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_4_add_exe), .data_out(_add_map_x_4_data_out), .data_out_index(_add_map_x_4_data_out_index), .data_near(_add_map_x_4_data_near), .wall_t_out(_add_map_x_4_wall_t_out), .data_org(_add_map_x_4_data_org), .data_org_near(_add_map_x_4_data_org_near), .s_g(_add_map_x_4_s_g), .s_g_near(_add_map_x_4_s_g_near), .moto_org_near(_add_map_x_4_moto_org_near), .moto_org_near1(_add_map_x_4_moto_org_near1), .moto_org_near2(_add_map_x_4_moto_org_near2), .moto_org_near3(_add_map_x_4_moto_org_near3), .moto_org(_add_map_x_4_moto_org), .sg_up(_add_map_x_4_sg_up), .sg_down(_add_map_x_4_sg_down), .sg_left(_add_map_x_4_sg_left), .sg_right(_add_map_x_4_sg_right), .wall_t_in(_add_map_x_4_wall_t_in), .moto(_add_map_x_4_moto), .up(_add_map_x_4_up), .right(_add_map_x_4_right), .down(_add_map_x_4_down), .left(_add_map_x_4_left), .start(_add_map_x_4_start), .goal(_add_map_x_4_goal), .now(_add_map_x_4_now));
add_map add_map_x_3 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_3_add_exe), .data_out(_add_map_x_3_data_out), .data_out_index(_add_map_x_3_data_out_index), .data_near(_add_map_x_3_data_near), .wall_t_out(_add_map_x_3_wall_t_out), .data_org(_add_map_x_3_data_org), .data_org_near(_add_map_x_3_data_org_near), .s_g(_add_map_x_3_s_g), .s_g_near(_add_map_x_3_s_g_near), .moto_org_near(_add_map_x_3_moto_org_near), .moto_org_near1(_add_map_x_3_moto_org_near1), .moto_org_near2(_add_map_x_3_moto_org_near2), .moto_org_near3(_add_map_x_3_moto_org_near3), .moto_org(_add_map_x_3_moto_org), .sg_up(_add_map_x_3_sg_up), .sg_down(_add_map_x_3_sg_down), .sg_left(_add_map_x_3_sg_left), .sg_right(_add_map_x_3_sg_right), .wall_t_in(_add_map_x_3_wall_t_in), .moto(_add_map_x_3_moto), .up(_add_map_x_3_up), .right(_add_map_x_3_right), .down(_add_map_x_3_down), .left(_add_map_x_3_left), .start(_add_map_x_3_start), .goal(_add_map_x_3_goal), .now(_add_map_x_3_now));
add_map add_map_x_2 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_2_add_exe), .data_out(_add_map_x_2_data_out), .data_out_index(_add_map_x_2_data_out_index), .data_near(_add_map_x_2_data_near), .wall_t_out(_add_map_x_2_wall_t_out), .data_org(_add_map_x_2_data_org), .data_org_near(_add_map_x_2_data_org_near), .s_g(_add_map_x_2_s_g), .s_g_near(_add_map_x_2_s_g_near), .moto_org_near(_add_map_x_2_moto_org_near), .moto_org_near1(_add_map_x_2_moto_org_near1), .moto_org_near2(_add_map_x_2_moto_org_near2), .moto_org_near3(_add_map_x_2_moto_org_near3), .moto_org(_add_map_x_2_moto_org), .sg_up(_add_map_x_2_sg_up), .sg_down(_add_map_x_2_sg_down), .sg_left(_add_map_x_2_sg_left), .sg_right(_add_map_x_2_sg_right), .wall_t_in(_add_map_x_2_wall_t_in), .moto(_add_map_x_2_moto), .up(_add_map_x_2_up), .right(_add_map_x_2_right), .down(_add_map_x_2_down), .left(_add_map_x_2_left), .start(_add_map_x_2_start), .goal(_add_map_x_2_goal), .now(_add_map_x_2_now));
add_map add_map_x_1 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_1_add_exe), .data_out(_add_map_x_1_data_out), .data_out_index(_add_map_x_1_data_out_index), .data_near(_add_map_x_1_data_near), .wall_t_out(_add_map_x_1_wall_t_out), .data_org(_add_map_x_1_data_org), .data_org_near(_add_map_x_1_data_org_near), .s_g(_add_map_x_1_s_g), .s_g_near(_add_map_x_1_s_g_near), .moto_org_near(_add_map_x_1_moto_org_near), .moto_org_near1(_add_map_x_1_moto_org_near1), .moto_org_near2(_add_map_x_1_moto_org_near2), .moto_org_near3(_add_map_x_1_moto_org_near3), .moto_org(_add_map_x_1_moto_org), .sg_up(_add_map_x_1_sg_up), .sg_down(_add_map_x_1_sg_down), .sg_left(_add_map_x_1_sg_left), .sg_right(_add_map_x_1_sg_right), .wall_t_in(_add_map_x_1_wall_t_in), .moto(_add_map_x_1_moto), .up(_add_map_x_1_up), .right(_add_map_x_1_right), .down(_add_map_x_1_down), .left(_add_map_x_1_left), .start(_add_map_x_1_start), .goal(_add_map_x_1_goal), .now(_add_map_x_1_now));

   assign  _add_map_x_moto_org_near = ((_net_4013)?data_in_org34:10'b0)|
    ((_net_21)?data_in_org33:10'b0);
   assign  _add_map_x_moto_org_near1 = ((_net_4012)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_20)?data_in_org35:10'b0);
   assign  _add_map_x_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_moto_org_near3 = ((_net_4010)?data_in_org65:10'b0)|
    ((_net_18)?data_in_org66:10'b0);
   assign  _add_map_x_moto_org = ((_net_4009)?data_in_org33:10'b0)|
    ((_net_17)?data_in_org34:10'b0);
   assign  _add_map_x_sg_up = ((_net_4008)?sg_in34:2'b0)|
    ((_net_16)?sg_in33:2'b0);
   assign  _add_map_x_sg_down = ((_net_4007)?3'b000:2'b0)|
    ((_net_15)?sg_in35:2'b0);
   assign  _add_map_x_sg_left = ((_net_4005)?sg_in65:2'b0)|
    ((_net_13)?sg_in66:2'b0);
   assign  _add_map_x_sg_right = 3'b000;
   assign  _add_map_x_wall_t_in = dig_w;
   assign  _add_map_x_moto = ((_net_4003)?data_in33:10'b0)|
    ((_net_11)?data_in34:10'b0);
   assign  _add_map_x_up = ((_net_4002)?data_in34:10'b0)|
    ((_net_10)?data_in33:10'b0);
   assign  _add_map_x_right = ((_net_4001)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_9)?data_in35:10'b0);
   assign  _add_map_x_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_left = ((_net_3999)?data_in65:10'b0)|
    ((_net_7)?data_in66:10'b0);
   assign  _add_map_x_start = start;
   assign  _add_map_x_goal = goal;
   assign  _add_map_x_now = ((_net_3996)?10'b0000100001:10'b0)|
    ((_net_4)?10'b0000100010:10'b0);
   assign  _add_map_x_add_exe = (_net_3995|_net_3);
   assign  _add_map_x_p_reset = p_reset;
   assign  _add_map_x_m_clock = m_clock;
   assign  _add_map_x_209_moto_org_near = ((_net_7984)?data_in_org477:10'b0)|
    ((_net_3992)?data_in_org478:10'b0);
   assign  _add_map_x_209_moto_org_near1 = ((_net_7983)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_3991)?data_in_org476:10'b0);
   assign  _add_map_x_209_moto_org_near2 = ((_net_7982)?data_in_org446:10'b0)|
    ((_net_3990)?data_in_org445:10'b0);
   assign  _add_map_x_209_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_209_moto_org = ((_net_7980)?data_in_org478:10'b0)|
    ((_net_3988)?data_in_org477:10'b0);
   assign  _add_map_x_209_sg_up = ((_net_7979)?sg_in477:2'b0)|
    ((_net_3987)?sg_in478:2'b0);
   assign  _add_map_x_209_sg_down = ((_net_7978)?3'b000:2'b0)|
    ((_net_3986)?sg_in476:2'b0);
   assign  _add_map_x_209_sg_left = 3'b000;
   assign  _add_map_x_209_sg_right = ((_net_7977)?sg_in446:2'b0)|
    ((_net_3985)?sg_in445:2'b0);
   assign  _add_map_x_209_wall_t_in = dig_w;
   assign  _add_map_x_209_moto = ((_net_7974)?data_in478:10'b0)|
    ((_net_3982)?data_in477:10'b0);
   assign  _add_map_x_209_up = ((_net_7973)?data_in477:10'b0)|
    ((_net_3981)?data_in478:10'b0);
   assign  _add_map_x_209_right = ((_net_7972)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_3980)?data_in476:10'b0);
   assign  _add_map_x_209_down = ((_net_7971)?data_in446:10'b0)|
    ((_net_3979)?data_in445:10'b0);
   assign  _add_map_x_209_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_209_start = start;
   assign  _add_map_x_209_goal = goal;
   assign  _add_map_x_209_now = ((_net_7967)?10'b0111011110:10'b0)|
    ((_net_3975)?10'b0111011101:10'b0);
   assign  _add_map_x_209_add_exe = (_net_7966|_net_3974);
   assign  _add_map_x_209_p_reset = p_reset;
   assign  _add_map_x_209_m_clock = m_clock;
   assign  _add_map_x_208_moto_org_near = ((_net_7965)?data_in_org475:10'b0)|
    ((_net_3973)?data_in_org476:10'b0);
   assign  _add_map_x_208_moto_org_near1 = ((_net_7964)?data_in_org477:10'b0)|
    ((_net_3972)?data_in_org474:10'b0);
   assign  _add_map_x_208_moto_org_near2 = ((_net_7963)?data_in_org444:10'b0)|
    ((_net_3971)?data_in_org443:10'b0);
   assign  _add_map_x_208_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_208_moto_org = ((_net_7961)?data_in_org476:10'b0)|
    ((_net_3969)?data_in_org475:10'b0);
   assign  _add_map_x_208_sg_up = ((_net_7960)?sg_in475:2'b0)|
    ((_net_3968)?sg_in476:2'b0);
   assign  _add_map_x_208_sg_down = ((_net_7959)?sg_in477:2'b0)|
    ((_net_3967)?sg_in474:2'b0);
   assign  _add_map_x_208_sg_left = 3'b000;
   assign  _add_map_x_208_sg_right = ((_net_7958)?sg_in444:2'b0)|
    ((_net_3966)?sg_in443:2'b0);
   assign  _add_map_x_208_wall_t_in = dig_w;
   assign  _add_map_x_208_moto = ((_net_7955)?data_in476:10'b0)|
    ((_net_3963)?data_in475:10'b0);
   assign  _add_map_x_208_up = ((_net_7954)?data_in475:10'b0)|
    ((_net_3962)?data_in476:10'b0);
   assign  _add_map_x_208_right = ((_net_7953)?data_in477:10'b0)|
    ((_net_3961)?data_in474:10'b0);
   assign  _add_map_x_208_down = ((_net_7952)?data_in444:10'b0)|
    ((_net_3960)?data_in443:10'b0);
   assign  _add_map_x_208_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_208_start = start;
   assign  _add_map_x_208_goal = goal;
   assign  _add_map_x_208_now = ((_net_7948)?10'b0111011100:10'b0)|
    ((_net_3956)?10'b0111011011:10'b0);
   assign  _add_map_x_208_add_exe = (_net_7947|_net_3955);
   assign  _add_map_x_208_p_reset = p_reset;
   assign  _add_map_x_208_m_clock = m_clock;
   assign  _add_map_x_207_moto_org_near = ((_net_7946)?data_in_org473:10'b0)|
    ((_net_3954)?data_in_org474:10'b0);
   assign  _add_map_x_207_moto_org_near1 = ((_net_7945)?data_in_org475:10'b0)|
    ((_net_3953)?data_in_org472:10'b0);
   assign  _add_map_x_207_moto_org_near2 = ((_net_7944)?data_in_org442:10'b0)|
    ((_net_3952)?data_in_org441:10'b0);
   assign  _add_map_x_207_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_207_moto_org = ((_net_7942)?data_in_org474:10'b0)|
    ((_net_3950)?data_in_org473:10'b0);
   assign  _add_map_x_207_sg_up = ((_net_7941)?sg_in473:2'b0)|
    ((_net_3949)?sg_in474:2'b0);
   assign  _add_map_x_207_sg_down = ((_net_7940)?sg_in475:2'b0)|
    ((_net_3948)?sg_in472:2'b0);
   assign  _add_map_x_207_sg_left = 3'b000;
   assign  _add_map_x_207_sg_right = ((_net_7939)?sg_in442:2'b0)|
    ((_net_3947)?sg_in441:2'b0);
   assign  _add_map_x_207_wall_t_in = dig_w;
   assign  _add_map_x_207_moto = ((_net_7936)?data_in474:10'b0)|
    ((_net_3944)?data_in473:10'b0);
   assign  _add_map_x_207_up = ((_net_7935)?data_in473:10'b0)|
    ((_net_3943)?data_in474:10'b0);
   assign  _add_map_x_207_right = ((_net_7934)?data_in475:10'b0)|
    ((_net_3942)?data_in472:10'b0);
   assign  _add_map_x_207_down = ((_net_7933)?data_in442:10'b0)|
    ((_net_3941)?data_in441:10'b0);
   assign  _add_map_x_207_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_207_start = start;
   assign  _add_map_x_207_goal = goal;
   assign  _add_map_x_207_now = ((_net_7929)?10'b0111011010:10'b0)|
    ((_net_3937)?10'b0111011001:10'b0);
   assign  _add_map_x_207_add_exe = (_net_7928|_net_3936);
   assign  _add_map_x_207_p_reset = p_reset;
   assign  _add_map_x_207_m_clock = m_clock;
   assign  _add_map_x_206_moto_org_near = ((_net_7927)?data_in_org471:10'b0)|
    ((_net_3935)?data_in_org472:10'b0);
   assign  _add_map_x_206_moto_org_near1 = ((_net_7926)?data_in_org473:10'b0)|
    ((_net_3934)?data_in_org470:10'b0);
   assign  _add_map_x_206_moto_org_near2 = ((_net_7925)?data_in_org440:10'b0)|
    ((_net_3933)?data_in_org439:10'b0);
   assign  _add_map_x_206_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_206_moto_org = ((_net_7923)?data_in_org472:10'b0)|
    ((_net_3931)?data_in_org471:10'b0);
   assign  _add_map_x_206_sg_up = ((_net_7922)?sg_in471:2'b0)|
    ((_net_3930)?sg_in472:2'b0);
   assign  _add_map_x_206_sg_down = ((_net_7921)?sg_in473:2'b0)|
    ((_net_3929)?sg_in470:2'b0);
   assign  _add_map_x_206_sg_left = 3'b000;
   assign  _add_map_x_206_sg_right = ((_net_7920)?sg_in440:2'b0)|
    ((_net_3928)?sg_in439:2'b0);
   assign  _add_map_x_206_wall_t_in = dig_w;
   assign  _add_map_x_206_moto = ((_net_7917)?data_in472:10'b0)|
    ((_net_3925)?data_in471:10'b0);
   assign  _add_map_x_206_up = ((_net_7916)?data_in471:10'b0)|
    ((_net_3924)?data_in472:10'b0);
   assign  _add_map_x_206_right = ((_net_7915)?data_in473:10'b0)|
    ((_net_3923)?data_in470:10'b0);
   assign  _add_map_x_206_down = ((_net_7914)?data_in440:10'b0)|
    ((_net_3922)?data_in439:10'b0);
   assign  _add_map_x_206_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_206_start = start;
   assign  _add_map_x_206_goal = goal;
   assign  _add_map_x_206_now = ((_net_7910)?10'b0111011000:10'b0)|
    ((_net_3918)?10'b0111010111:10'b0);
   assign  _add_map_x_206_add_exe = (_net_7909|_net_3917);
   assign  _add_map_x_206_p_reset = p_reset;
   assign  _add_map_x_206_m_clock = m_clock;
   assign  _add_map_x_205_moto_org_near = ((_net_7908)?data_in_org469:10'b0)|
    ((_net_3916)?data_in_org470:10'b0);
   assign  _add_map_x_205_moto_org_near1 = ((_net_7907)?data_in_org471:10'b0)|
    ((_net_3915)?data_in_org468:10'b0);
   assign  _add_map_x_205_moto_org_near2 = ((_net_7906)?data_in_org438:10'b0)|
    ((_net_3914)?data_in_org437:10'b0);
   assign  _add_map_x_205_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_205_moto_org = ((_net_7904)?data_in_org470:10'b0)|
    ((_net_3912)?data_in_org469:10'b0);
   assign  _add_map_x_205_sg_up = ((_net_7903)?sg_in469:2'b0)|
    ((_net_3911)?sg_in470:2'b0);
   assign  _add_map_x_205_sg_down = ((_net_7902)?sg_in471:2'b0)|
    ((_net_3910)?sg_in468:2'b0);
   assign  _add_map_x_205_sg_left = 3'b000;
   assign  _add_map_x_205_sg_right = ((_net_7901)?sg_in438:2'b0)|
    ((_net_3909)?sg_in437:2'b0);
   assign  _add_map_x_205_wall_t_in = dig_w;
   assign  _add_map_x_205_moto = ((_net_7898)?data_in470:10'b0)|
    ((_net_3906)?data_in469:10'b0);
   assign  _add_map_x_205_up = ((_net_7897)?data_in469:10'b0)|
    ((_net_3905)?data_in470:10'b0);
   assign  _add_map_x_205_right = ((_net_7896)?data_in471:10'b0)|
    ((_net_3904)?data_in468:10'b0);
   assign  _add_map_x_205_down = ((_net_7895)?data_in438:10'b0)|
    ((_net_3903)?data_in437:10'b0);
   assign  _add_map_x_205_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_205_start = start;
   assign  _add_map_x_205_goal = goal;
   assign  _add_map_x_205_now = ((_net_7891)?10'b0111010110:10'b0)|
    ((_net_3899)?10'b0111010101:10'b0);
   assign  _add_map_x_205_add_exe = (_net_7890|_net_3898);
   assign  _add_map_x_205_p_reset = p_reset;
   assign  _add_map_x_205_m_clock = m_clock;
   assign  _add_map_x_204_moto_org_near = ((_net_7889)?data_in_org467:10'b0)|
    ((_net_3897)?data_in_org468:10'b0);
   assign  _add_map_x_204_moto_org_near1 = ((_net_7888)?data_in_org469:10'b0)|
    ((_net_3896)?data_in_org466:10'b0);
   assign  _add_map_x_204_moto_org_near2 = ((_net_7887)?data_in_org436:10'b0)|
    ((_net_3895)?data_in_org435:10'b0);
   assign  _add_map_x_204_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_204_moto_org = ((_net_7885)?data_in_org468:10'b0)|
    ((_net_3893)?data_in_org467:10'b0);
   assign  _add_map_x_204_sg_up = ((_net_7884)?sg_in467:2'b0)|
    ((_net_3892)?sg_in468:2'b0);
   assign  _add_map_x_204_sg_down = ((_net_7883)?sg_in469:2'b0)|
    ((_net_3891)?sg_in466:2'b0);
   assign  _add_map_x_204_sg_left = 3'b000;
   assign  _add_map_x_204_sg_right = ((_net_7882)?sg_in436:2'b0)|
    ((_net_3890)?sg_in435:2'b0);
   assign  _add_map_x_204_wall_t_in = dig_w;
   assign  _add_map_x_204_moto = ((_net_7879)?data_in468:10'b0)|
    ((_net_3887)?data_in467:10'b0);
   assign  _add_map_x_204_up = ((_net_7878)?data_in467:10'b0)|
    ((_net_3886)?data_in468:10'b0);
   assign  _add_map_x_204_right = ((_net_7877)?data_in469:10'b0)|
    ((_net_3885)?data_in466:10'b0);
   assign  _add_map_x_204_down = ((_net_7876)?data_in436:10'b0)|
    ((_net_3884)?data_in435:10'b0);
   assign  _add_map_x_204_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_204_start = start;
   assign  _add_map_x_204_goal = goal;
   assign  _add_map_x_204_now = ((_net_7872)?10'b0111010100:10'b0)|
    ((_net_3880)?10'b0111010011:10'b0);
   assign  _add_map_x_204_add_exe = (_net_7871|_net_3879);
   assign  _add_map_x_204_p_reset = p_reset;
   assign  _add_map_x_204_m_clock = m_clock;
   assign  _add_map_x_203_moto_org_near = ((_net_7870)?data_in_org465:10'b0)|
    ((_net_3878)?data_in_org466:10'b0);
   assign  _add_map_x_203_moto_org_near1 = ((_net_7869)?data_in_org467:10'b0)|
    ((_net_3877)?data_in_org464:10'b0);
   assign  _add_map_x_203_moto_org_near2 = ((_net_7868)?data_in_org434:10'b0)|
    ((_net_3876)?data_in_org433:10'b0);
   assign  _add_map_x_203_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_203_moto_org = ((_net_7866)?data_in_org466:10'b0)|
    ((_net_3874)?data_in_org465:10'b0);
   assign  _add_map_x_203_sg_up = ((_net_7865)?sg_in465:2'b0)|
    ((_net_3873)?sg_in466:2'b0);
   assign  _add_map_x_203_sg_down = ((_net_7864)?sg_in467:2'b0)|
    ((_net_3872)?sg_in464:2'b0);
   assign  _add_map_x_203_sg_left = 3'b000;
   assign  _add_map_x_203_sg_right = ((_net_7863)?sg_in434:2'b0)|
    ((_net_3871)?sg_in433:2'b0);
   assign  _add_map_x_203_wall_t_in = dig_w;
   assign  _add_map_x_203_moto = ((_net_7860)?data_in466:10'b0)|
    ((_net_3868)?data_in465:10'b0);
   assign  _add_map_x_203_up = ((_net_7859)?data_in465:10'b0)|
    ((_net_3867)?data_in466:10'b0);
   assign  _add_map_x_203_right = ((_net_7858)?data_in467:10'b0)|
    ((_net_3866)?data_in464:10'b0);
   assign  _add_map_x_203_down = ((_net_7857)?data_in434:10'b0)|
    ((_net_3865)?data_in433:10'b0);
   assign  _add_map_x_203_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_203_start = start;
   assign  _add_map_x_203_goal = goal;
   assign  _add_map_x_203_now = ((_net_7853)?10'b0111010010:10'b0)|
    ((_net_3861)?10'b0111010001:10'b0);
   assign  _add_map_x_203_add_exe = (_net_7852|_net_3860);
   assign  _add_map_x_203_p_reset = p_reset;
   assign  _add_map_x_203_m_clock = m_clock;
   assign  _add_map_x_202_moto_org_near = ((_net_7851)?data_in_org463:10'b0)|
    ((_net_3859)?data_in_org464:10'b0);
   assign  _add_map_x_202_moto_org_near1 = ((_net_7850)?data_in_org465:10'b0)|
    ((_net_3858)?data_in_org462:10'b0);
   assign  _add_map_x_202_moto_org_near2 = ((_net_7849)?data_in_org432:10'b0)|
    ((_net_3857)?data_in_org431:10'b0);
   assign  _add_map_x_202_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_202_moto_org = ((_net_7847)?data_in_org464:10'b0)|
    ((_net_3855)?data_in_org463:10'b0);
   assign  _add_map_x_202_sg_up = ((_net_7846)?sg_in463:2'b0)|
    ((_net_3854)?sg_in464:2'b0);
   assign  _add_map_x_202_sg_down = ((_net_7845)?sg_in465:2'b0)|
    ((_net_3853)?sg_in462:2'b0);
   assign  _add_map_x_202_sg_left = 3'b000;
   assign  _add_map_x_202_sg_right = ((_net_7844)?sg_in432:2'b0)|
    ((_net_3852)?sg_in431:2'b0);
   assign  _add_map_x_202_wall_t_in = dig_w;
   assign  _add_map_x_202_moto = ((_net_7841)?data_in464:10'b0)|
    ((_net_3849)?data_in463:10'b0);
   assign  _add_map_x_202_up = ((_net_7840)?data_in463:10'b0)|
    ((_net_3848)?data_in464:10'b0);
   assign  _add_map_x_202_right = ((_net_7839)?data_in465:10'b0)|
    ((_net_3847)?data_in462:10'b0);
   assign  _add_map_x_202_down = ((_net_7838)?data_in432:10'b0)|
    ((_net_3846)?data_in431:10'b0);
   assign  _add_map_x_202_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_202_start = start;
   assign  _add_map_x_202_goal = goal;
   assign  _add_map_x_202_now = ((_net_7834)?10'b0111010000:10'b0)|
    ((_net_3842)?10'b0111001111:10'b0);
   assign  _add_map_x_202_add_exe = (_net_7833|_net_3841);
   assign  _add_map_x_202_p_reset = p_reset;
   assign  _add_map_x_202_m_clock = m_clock;
   assign  _add_map_x_201_moto_org_near = ((_net_7832)?data_in_org461:10'b0)|
    ((_net_3840)?data_in_org462:10'b0);
   assign  _add_map_x_201_moto_org_near1 = ((_net_7831)?data_in_org463:10'b0)|
    ((_net_3839)?data_in_org460:10'b0);
   assign  _add_map_x_201_moto_org_near2 = ((_net_7830)?data_in_org430:10'b0)|
    ((_net_3838)?data_in_org429:10'b0);
   assign  _add_map_x_201_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_201_moto_org = ((_net_7828)?data_in_org462:10'b0)|
    ((_net_3836)?data_in_org461:10'b0);
   assign  _add_map_x_201_sg_up = ((_net_7827)?sg_in461:2'b0)|
    ((_net_3835)?sg_in462:2'b0);
   assign  _add_map_x_201_sg_down = ((_net_7826)?sg_in463:2'b0)|
    ((_net_3834)?sg_in460:2'b0);
   assign  _add_map_x_201_sg_left = 3'b000;
   assign  _add_map_x_201_sg_right = ((_net_7825)?sg_in430:2'b0)|
    ((_net_3833)?sg_in429:2'b0);
   assign  _add_map_x_201_wall_t_in = dig_w;
   assign  _add_map_x_201_moto = ((_net_7822)?data_in462:10'b0)|
    ((_net_3830)?data_in461:10'b0);
   assign  _add_map_x_201_up = ((_net_7821)?data_in461:10'b0)|
    ((_net_3829)?data_in462:10'b0);
   assign  _add_map_x_201_right = ((_net_7820)?data_in463:10'b0)|
    ((_net_3828)?data_in460:10'b0);
   assign  _add_map_x_201_down = ((_net_7819)?data_in430:10'b0)|
    ((_net_3827)?data_in429:10'b0);
   assign  _add_map_x_201_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_201_start = start;
   assign  _add_map_x_201_goal = goal;
   assign  _add_map_x_201_now = ((_net_7815)?10'b0111001110:10'b0)|
    ((_net_3823)?10'b0111001101:10'b0);
   assign  _add_map_x_201_add_exe = (_net_7814|_net_3822);
   assign  _add_map_x_201_p_reset = p_reset;
   assign  _add_map_x_201_m_clock = m_clock;
   assign  _add_map_x_200_moto_org_near = ((_net_7813)?data_in_org459:10'b0)|
    ((_net_3821)?data_in_org460:10'b0);
   assign  _add_map_x_200_moto_org_near1 = ((_net_7812)?data_in_org461:10'b0)|
    ((_net_3820)?data_in_org458:10'b0);
   assign  _add_map_x_200_moto_org_near2 = ((_net_7811)?data_in_org428:10'b0)|
    ((_net_3819)?data_in_org427:10'b0);
   assign  _add_map_x_200_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_200_moto_org = ((_net_7809)?data_in_org460:10'b0)|
    ((_net_3817)?data_in_org459:10'b0);
   assign  _add_map_x_200_sg_up = ((_net_7808)?sg_in459:2'b0)|
    ((_net_3816)?sg_in460:2'b0);
   assign  _add_map_x_200_sg_down = ((_net_7807)?sg_in461:2'b0)|
    ((_net_3815)?sg_in458:2'b0);
   assign  _add_map_x_200_sg_left = 3'b000;
   assign  _add_map_x_200_sg_right = ((_net_7806)?sg_in428:2'b0)|
    ((_net_3814)?sg_in427:2'b0);
   assign  _add_map_x_200_wall_t_in = dig_w;
   assign  _add_map_x_200_moto = ((_net_7803)?data_in460:10'b0)|
    ((_net_3811)?data_in459:10'b0);
   assign  _add_map_x_200_up = ((_net_7802)?data_in459:10'b0)|
    ((_net_3810)?data_in460:10'b0);
   assign  _add_map_x_200_right = ((_net_7801)?data_in461:10'b0)|
    ((_net_3809)?data_in458:10'b0);
   assign  _add_map_x_200_down = ((_net_7800)?data_in428:10'b0)|
    ((_net_3808)?data_in427:10'b0);
   assign  _add_map_x_200_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_200_start = start;
   assign  _add_map_x_200_goal = goal;
   assign  _add_map_x_200_now = ((_net_7796)?10'b0111001100:10'b0)|
    ((_net_3804)?10'b0111001011:10'b0);
   assign  _add_map_x_200_add_exe = (_net_7795|_net_3803);
   assign  _add_map_x_200_p_reset = p_reset;
   assign  _add_map_x_200_m_clock = m_clock;
   assign  _add_map_x_199_moto_org_near = ((_net_7794)?data_in_org457:10'b0)|
    ((_net_3802)?data_in_org458:10'b0);
   assign  _add_map_x_199_moto_org_near1 = ((_net_7793)?data_in_org459:10'b0)|
    ((_net_3801)?data_in_org456:10'b0);
   assign  _add_map_x_199_moto_org_near2 = ((_net_7792)?data_in_org426:10'b0)|
    ((_net_3800)?data_in_org425:10'b0);
   assign  _add_map_x_199_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_199_moto_org = ((_net_7790)?data_in_org458:10'b0)|
    ((_net_3798)?data_in_org457:10'b0);
   assign  _add_map_x_199_sg_up = ((_net_7789)?sg_in457:2'b0)|
    ((_net_3797)?sg_in458:2'b0);
   assign  _add_map_x_199_sg_down = ((_net_7788)?sg_in459:2'b0)|
    ((_net_3796)?sg_in456:2'b0);
   assign  _add_map_x_199_sg_left = 3'b000;
   assign  _add_map_x_199_sg_right = ((_net_7787)?sg_in426:2'b0)|
    ((_net_3795)?sg_in425:2'b0);
   assign  _add_map_x_199_wall_t_in = dig_w;
   assign  _add_map_x_199_moto = ((_net_7784)?data_in458:10'b0)|
    ((_net_3792)?data_in457:10'b0);
   assign  _add_map_x_199_up = ((_net_7783)?data_in457:10'b0)|
    ((_net_3791)?data_in458:10'b0);
   assign  _add_map_x_199_right = ((_net_7782)?data_in459:10'b0)|
    ((_net_3790)?data_in456:10'b0);
   assign  _add_map_x_199_down = ((_net_7781)?data_in426:10'b0)|
    ((_net_3789)?data_in425:10'b0);
   assign  _add_map_x_199_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_199_start = start;
   assign  _add_map_x_199_goal = goal;
   assign  _add_map_x_199_now = ((_net_7777)?10'b0111001010:10'b0)|
    ((_net_3785)?10'b0111001001:10'b0);
   assign  _add_map_x_199_add_exe = (_net_7776|_net_3784);
   assign  _add_map_x_199_p_reset = p_reset;
   assign  _add_map_x_199_m_clock = m_clock;
   assign  _add_map_x_198_moto_org_near = ((_net_7775)?data_in_org455:10'b0)|
    ((_net_3783)?data_in_org456:10'b0);
   assign  _add_map_x_198_moto_org_near1 = ((_net_7774)?data_in_org457:10'b0)|
    ((_net_3782)?data_in_org454:10'b0);
   assign  _add_map_x_198_moto_org_near2 = ((_net_7773)?data_in_org424:10'b0)|
    ((_net_3781)?data_in_org423:10'b0);
   assign  _add_map_x_198_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_198_moto_org = ((_net_7771)?data_in_org456:10'b0)|
    ((_net_3779)?data_in_org455:10'b0);
   assign  _add_map_x_198_sg_up = ((_net_7770)?sg_in455:2'b0)|
    ((_net_3778)?sg_in456:2'b0);
   assign  _add_map_x_198_sg_down = ((_net_7769)?sg_in457:2'b0)|
    ((_net_3777)?sg_in454:2'b0);
   assign  _add_map_x_198_sg_left = 3'b000;
   assign  _add_map_x_198_sg_right = ((_net_7768)?sg_in424:2'b0)|
    ((_net_3776)?sg_in423:2'b0);
   assign  _add_map_x_198_wall_t_in = dig_w;
   assign  _add_map_x_198_moto = ((_net_7765)?data_in456:10'b0)|
    ((_net_3773)?data_in455:10'b0);
   assign  _add_map_x_198_up = ((_net_7764)?data_in455:10'b0)|
    ((_net_3772)?data_in456:10'b0);
   assign  _add_map_x_198_right = ((_net_7763)?data_in457:10'b0)|
    ((_net_3771)?data_in454:10'b0);
   assign  _add_map_x_198_down = ((_net_7762)?data_in424:10'b0)|
    ((_net_3770)?data_in423:10'b0);
   assign  _add_map_x_198_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_198_start = start;
   assign  _add_map_x_198_goal = goal;
   assign  _add_map_x_198_now = ((_net_7758)?10'b0111001000:10'b0)|
    ((_net_3766)?10'b0111000111:10'b0);
   assign  _add_map_x_198_add_exe = (_net_7757|_net_3765);
   assign  _add_map_x_198_p_reset = p_reset;
   assign  _add_map_x_198_m_clock = m_clock;
   assign  _add_map_x_197_moto_org_near = ((_net_7756)?data_in_org453:10'b0)|
    ((_net_3764)?data_in_org454:10'b0);
   assign  _add_map_x_197_moto_org_near1 = ((_net_7755)?data_in_org455:10'b0)|
    ((_net_3763)?data_in_org452:10'b0);
   assign  _add_map_x_197_moto_org_near2 = ((_net_7754)?data_in_org422:10'b0)|
    ((_net_3762)?data_in_org421:10'b0);
   assign  _add_map_x_197_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_197_moto_org = ((_net_7752)?data_in_org454:10'b0)|
    ((_net_3760)?data_in_org453:10'b0);
   assign  _add_map_x_197_sg_up = ((_net_7751)?sg_in453:2'b0)|
    ((_net_3759)?sg_in454:2'b0);
   assign  _add_map_x_197_sg_down = ((_net_7750)?sg_in455:2'b0)|
    ((_net_3758)?sg_in452:2'b0);
   assign  _add_map_x_197_sg_left = 3'b000;
   assign  _add_map_x_197_sg_right = ((_net_7749)?sg_in422:2'b0)|
    ((_net_3757)?sg_in421:2'b0);
   assign  _add_map_x_197_wall_t_in = dig_w;
   assign  _add_map_x_197_moto = ((_net_7746)?data_in454:10'b0)|
    ((_net_3754)?data_in453:10'b0);
   assign  _add_map_x_197_up = ((_net_7745)?data_in453:10'b0)|
    ((_net_3753)?data_in454:10'b0);
   assign  _add_map_x_197_right = ((_net_7744)?data_in455:10'b0)|
    ((_net_3752)?data_in452:10'b0);
   assign  _add_map_x_197_down = ((_net_7743)?data_in422:10'b0)|
    ((_net_3751)?data_in421:10'b0);
   assign  _add_map_x_197_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_197_start = start;
   assign  _add_map_x_197_goal = goal;
   assign  _add_map_x_197_now = ((_net_7739)?10'b0111000110:10'b0)|
    ((_net_3747)?10'b0111000101:10'b0);
   assign  _add_map_x_197_add_exe = (_net_7738|_net_3746);
   assign  _add_map_x_197_p_reset = p_reset;
   assign  _add_map_x_197_m_clock = m_clock;
   assign  _add_map_x_196_moto_org_near = ((_net_7737)?data_in_org451:10'b0)|
    ((_net_3745)?data_in_org452:10'b0);
   assign  _add_map_x_196_moto_org_near1 = ((_net_7736)?data_in_org453:10'b0)|
    ((_net_3744)?data_in_org450:10'b0);
   assign  _add_map_x_196_moto_org_near2 = ((_net_7735)?data_in_org420:10'b0)|
    ((_net_3743)?data_in_org419:10'b0);
   assign  _add_map_x_196_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_196_moto_org = ((_net_7733)?data_in_org452:10'b0)|
    ((_net_3741)?data_in_org451:10'b0);
   assign  _add_map_x_196_sg_up = ((_net_7732)?sg_in451:2'b0)|
    ((_net_3740)?sg_in452:2'b0);
   assign  _add_map_x_196_sg_down = ((_net_7731)?sg_in453:2'b0)|
    ((_net_3739)?sg_in450:2'b0);
   assign  _add_map_x_196_sg_left = 3'b000;
   assign  _add_map_x_196_sg_right = ((_net_7730)?sg_in420:2'b0)|
    ((_net_3738)?sg_in419:2'b0);
   assign  _add_map_x_196_wall_t_in = dig_w;
   assign  _add_map_x_196_moto = ((_net_7727)?data_in452:10'b0)|
    ((_net_3735)?data_in451:10'b0);
   assign  _add_map_x_196_up = ((_net_7726)?data_in451:10'b0)|
    ((_net_3734)?data_in452:10'b0);
   assign  _add_map_x_196_right = ((_net_7725)?data_in453:10'b0)|
    ((_net_3733)?data_in450:10'b0);
   assign  _add_map_x_196_down = ((_net_7724)?data_in420:10'b0)|
    ((_net_3732)?data_in419:10'b0);
   assign  _add_map_x_196_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_196_start = start;
   assign  _add_map_x_196_goal = goal;
   assign  _add_map_x_196_now = ((_net_7720)?10'b0111000100:10'b0)|
    ((_net_3728)?10'b0111000011:10'b0);
   assign  _add_map_x_196_add_exe = (_net_7719|_net_3727);
   assign  _add_map_x_196_p_reset = p_reset;
   assign  _add_map_x_196_m_clock = m_clock;
   assign  _add_map_x_195_moto_org_near = ((_net_7718)?data_in_org449:10'b0)|
    ((_net_3726)?data_in_org450:10'b0);
   assign  _add_map_x_195_moto_org_near1 = ((_net_7717)?data_in_org451:10'b0)|
    ((_net_3725)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_195_moto_org_near2 = ((_net_7716)?data_in_org418:10'b0)|
    ((_net_3724)?data_in_org417:10'b0);
   assign  _add_map_x_195_moto_org_near3 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_195_moto_org = ((_net_7714)?data_in_org450:10'b0)|
    ((_net_3722)?data_in_org449:10'b0);
   assign  _add_map_x_195_sg_up = ((_net_7713)?sg_in449:2'b0)|
    ((_net_3721)?sg_in450:2'b0);
   assign  _add_map_x_195_sg_down = ((_net_7712)?sg_in451:2'b0)|
    ((_net_3720)?3'b000:2'b0);
   assign  _add_map_x_195_sg_left = 3'b000;
   assign  _add_map_x_195_sg_right = ((_net_7711)?sg_in418:2'b0)|
    ((_net_3719)?sg_in417:2'b0);
   assign  _add_map_x_195_wall_t_in = dig_w;
   assign  _add_map_x_195_moto = ((_net_7708)?data_in450:10'b0)|
    ((_net_3716)?data_in449:10'b0);
   assign  _add_map_x_195_up = ((_net_7707)?data_in449:10'b0)|
    ((_net_3715)?data_in450:10'b0);
   assign  _add_map_x_195_right = ((_net_7706)?data_in451:10'b0)|
    ((_net_3714)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_195_down = ((_net_7705)?data_in418:10'b0)|
    ((_net_3713)?data_in417:10'b0);
   assign  _add_map_x_195_left = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_195_start = start;
   assign  _add_map_x_195_goal = goal;
   assign  _add_map_x_195_now = ((_net_7701)?10'b0111000010:10'b0)|
    ((_net_3709)?10'b0111000001:10'b0);
   assign  _add_map_x_195_add_exe = (_net_7700|_net_3708);
   assign  _add_map_x_195_p_reset = p_reset;
   assign  _add_map_x_195_m_clock = m_clock;
   assign  _add_map_x_194_moto_org_near = ((_net_7699)?data_in_org446:10'b0)|
    ((_net_3707)?data_in_org445:10'b0);
   assign  _add_map_x_194_moto_org_near1 = ((_net_7698)?data_in_org444:10'b0)|
    ((_net_3706)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_194_moto_org_near2 = ((_net_7697)?data_in_org413:10'b0)|
    ((_net_3705)?data_in_org414:10'b0);
   assign  _add_map_x_194_moto_org_near3 = ((_net_7696)?data_in_org477:10'b0)|
    ((_net_3704)?data_in_org478:10'b0);
   assign  _add_map_x_194_moto_org = ((_net_7695)?data_in_org445:10'b0)|
    ((_net_3703)?data_in_org446:10'b0);
   assign  _add_map_x_194_sg_up = ((_net_7694)?sg_in446:2'b0)|
    ((_net_3702)?sg_in445:2'b0);
   assign  _add_map_x_194_sg_down = ((_net_7693)?sg_in413:2'b0)|
    ((_net_3701)?3'b000:2'b0);
   assign  _add_map_x_194_sg_left = ((_net_7691)?sg_in477:2'b0)|
    ((_net_3699)?sg_in478:2'b0);
   assign  _add_map_x_194_sg_right = ((_net_7692)?sg_in444:2'b0)|
    ((_net_3700)?sg_in414:2'b0);
   assign  _add_map_x_194_wall_t_in = dig_w;
   assign  _add_map_x_194_moto = ((_net_7689)?data_in445:10'b0)|
    ((_net_3697)?data_in446:10'b0);
   assign  _add_map_x_194_up = ((_net_7688)?data_in446:10'b0)|
    ((_net_3696)?data_in445:10'b0);
   assign  _add_map_x_194_right = ((_net_7687)?data_in444:10'b0)|
    ((_net_3695)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_194_down = ((_net_7686)?data_in413:10'b0)|
    ((_net_3694)?data_in414:10'b0);
   assign  _add_map_x_194_left = ((_net_7685)?data_in477:10'b0)|
    ((_net_3693)?data_in478:10'b0);
   assign  _add_map_x_194_start = start;
   assign  _add_map_x_194_goal = goal;
   assign  _add_map_x_194_now = ((_net_7682)?10'b0110111101:10'b0)|
    ((_net_3690)?10'b0110111110:10'b0);
   assign  _add_map_x_194_add_exe = (_net_7681|_net_3689);
   assign  _add_map_x_194_p_reset = p_reset;
   assign  _add_map_x_194_m_clock = m_clock;
   assign  _add_map_x_193_moto_org_near = ((_net_7680)?data_in_org444:10'b0)|
    ((_net_3688)?data_in_org443:10'b0);
   assign  _add_map_x_193_moto_org_near1 = ((_net_7679)?data_in_org442:10'b0)|
    ((_net_3687)?data_in_org445:10'b0);
   assign  _add_map_x_193_moto_org_near2 = ((_net_7678)?data_in_org411:10'b0)|
    ((_net_3686)?data_in_org412:10'b0);
   assign  _add_map_x_193_moto_org_near3 = ((_net_7677)?data_in_org475:10'b0)|
    ((_net_3685)?data_in_org476:10'b0);
   assign  _add_map_x_193_moto_org = ((_net_7676)?data_in_org443:10'b0)|
    ((_net_3684)?data_in_org444:10'b0);
   assign  _add_map_x_193_sg_up = ((_net_7675)?sg_in444:2'b0)|
    ((_net_3683)?sg_in443:2'b0);
   assign  _add_map_x_193_sg_down = ((_net_7674)?sg_in411:2'b0)|
    ((_net_3682)?sg_in445:2'b0);
   assign  _add_map_x_193_sg_left = ((_net_7672)?sg_in475:2'b0)|
    ((_net_3680)?sg_in476:2'b0);
   assign  _add_map_x_193_sg_right = ((_net_7673)?sg_in442:2'b0)|
    ((_net_3681)?sg_in412:2'b0);
   assign  _add_map_x_193_wall_t_in = dig_w;
   assign  _add_map_x_193_moto = ((_net_7670)?data_in443:10'b0)|
    ((_net_3678)?data_in444:10'b0);
   assign  _add_map_x_193_up = ((_net_7669)?data_in444:10'b0)|
    ((_net_3677)?data_in443:10'b0);
   assign  _add_map_x_193_right = ((_net_7668)?data_in442:10'b0)|
    ((_net_3676)?data_in445:10'b0);
   assign  _add_map_x_193_down = ((_net_7667)?data_in411:10'b0)|
    ((_net_3675)?data_in412:10'b0);
   assign  _add_map_x_193_left = ((_net_7666)?data_in475:10'b0)|
    ((_net_3674)?data_in476:10'b0);
   assign  _add_map_x_193_start = start;
   assign  _add_map_x_193_goal = goal;
   assign  _add_map_x_193_now = ((_net_7663)?10'b0110111011:10'b0)|
    ((_net_3671)?10'b0110111100:10'b0);
   assign  _add_map_x_193_add_exe = (_net_7662|_net_3670);
   assign  _add_map_x_193_p_reset = p_reset;
   assign  _add_map_x_193_m_clock = m_clock;
   assign  _add_map_x_192_moto_org_near = ((_net_7661)?data_in_org442:10'b0)|
    ((_net_3669)?data_in_org441:10'b0);
   assign  _add_map_x_192_moto_org_near1 = ((_net_7660)?data_in_org440:10'b0)|
    ((_net_3668)?data_in_org443:10'b0);
   assign  _add_map_x_192_moto_org_near2 = ((_net_7659)?data_in_org409:10'b0)|
    ((_net_3667)?data_in_org410:10'b0);
   assign  _add_map_x_192_moto_org_near3 = ((_net_7658)?data_in_org473:10'b0)|
    ((_net_3666)?data_in_org474:10'b0);
   assign  _add_map_x_192_moto_org = ((_net_7657)?data_in_org441:10'b0)|
    ((_net_3665)?data_in_org442:10'b0);
   assign  _add_map_x_192_sg_up = ((_net_7656)?sg_in442:2'b0)|
    ((_net_3664)?sg_in441:2'b0);
   assign  _add_map_x_192_sg_down = ((_net_7655)?sg_in409:2'b0)|
    ((_net_3663)?sg_in443:2'b0);
   assign  _add_map_x_192_sg_left = ((_net_7653)?sg_in473:2'b0)|
    ((_net_3661)?sg_in474:2'b0);
   assign  _add_map_x_192_sg_right = ((_net_7654)?sg_in440:2'b0)|
    ((_net_3662)?sg_in410:2'b0);
   assign  _add_map_x_192_wall_t_in = dig_w;
   assign  _add_map_x_192_moto = ((_net_7651)?data_in441:10'b0)|
    ((_net_3659)?data_in442:10'b0);
   assign  _add_map_x_192_up = ((_net_7650)?data_in442:10'b0)|
    ((_net_3658)?data_in441:10'b0);
   assign  _add_map_x_192_right = ((_net_7649)?data_in440:10'b0)|
    ((_net_3657)?data_in443:10'b0);
   assign  _add_map_x_192_down = ((_net_7648)?data_in409:10'b0)|
    ((_net_3656)?data_in410:10'b0);
   assign  _add_map_x_192_left = ((_net_7647)?data_in473:10'b0)|
    ((_net_3655)?data_in474:10'b0);
   assign  _add_map_x_192_start = start;
   assign  _add_map_x_192_goal = goal;
   assign  _add_map_x_192_now = ((_net_7644)?10'b0110111001:10'b0)|
    ((_net_3652)?10'b0110111010:10'b0);
   assign  _add_map_x_192_add_exe = (_net_7643|_net_3651);
   assign  _add_map_x_192_p_reset = p_reset;
   assign  _add_map_x_192_m_clock = m_clock;
   assign  _add_map_x_191_moto_org_near = ((_net_7642)?data_in_org440:10'b0)|
    ((_net_3650)?data_in_org439:10'b0);
   assign  _add_map_x_191_moto_org_near1 = ((_net_7641)?data_in_org438:10'b0)|
    ((_net_3649)?data_in_org441:10'b0);
   assign  _add_map_x_191_moto_org_near2 = ((_net_7640)?data_in_org407:10'b0)|
    ((_net_3648)?data_in_org408:10'b0);
   assign  _add_map_x_191_moto_org_near3 = ((_net_7639)?data_in_org471:10'b0)|
    ((_net_3647)?data_in_org472:10'b0);
   assign  _add_map_x_191_moto_org = ((_net_7638)?data_in_org439:10'b0)|
    ((_net_3646)?data_in_org440:10'b0);
   assign  _add_map_x_191_sg_up = ((_net_7637)?sg_in440:2'b0)|
    ((_net_3645)?sg_in439:2'b0);
   assign  _add_map_x_191_sg_down = ((_net_7636)?sg_in407:2'b0)|
    ((_net_3644)?sg_in441:2'b0);
   assign  _add_map_x_191_sg_left = ((_net_7634)?sg_in471:2'b0)|
    ((_net_3642)?sg_in472:2'b0);
   assign  _add_map_x_191_sg_right = ((_net_7635)?sg_in438:2'b0)|
    ((_net_3643)?sg_in408:2'b0);
   assign  _add_map_x_191_wall_t_in = dig_w;
   assign  _add_map_x_191_moto = ((_net_7632)?data_in439:10'b0)|
    ((_net_3640)?data_in440:10'b0);
   assign  _add_map_x_191_up = ((_net_7631)?data_in440:10'b0)|
    ((_net_3639)?data_in439:10'b0);
   assign  _add_map_x_191_right = ((_net_7630)?data_in438:10'b0)|
    ((_net_3638)?data_in441:10'b0);
   assign  _add_map_x_191_down = ((_net_7629)?data_in407:10'b0)|
    ((_net_3637)?data_in408:10'b0);
   assign  _add_map_x_191_left = ((_net_7628)?data_in471:10'b0)|
    ((_net_3636)?data_in472:10'b0);
   assign  _add_map_x_191_start = start;
   assign  _add_map_x_191_goal = goal;
   assign  _add_map_x_191_now = ((_net_7625)?10'b0110110111:10'b0)|
    ((_net_3633)?10'b0110111000:10'b0);
   assign  _add_map_x_191_add_exe = (_net_7624|_net_3632);
   assign  _add_map_x_191_p_reset = p_reset;
   assign  _add_map_x_191_m_clock = m_clock;
   assign  _add_map_x_190_moto_org_near = ((_net_7623)?data_in_org438:10'b0)|
    ((_net_3631)?data_in_org437:10'b0);
   assign  _add_map_x_190_moto_org_near1 = ((_net_7622)?data_in_org436:10'b0)|
    ((_net_3630)?data_in_org439:10'b0);
   assign  _add_map_x_190_moto_org_near2 = ((_net_7621)?data_in_org405:10'b0)|
    ((_net_3629)?data_in_org406:10'b0);
   assign  _add_map_x_190_moto_org_near3 = ((_net_7620)?data_in_org469:10'b0)|
    ((_net_3628)?data_in_org470:10'b0);
   assign  _add_map_x_190_moto_org = ((_net_7619)?data_in_org437:10'b0)|
    ((_net_3627)?data_in_org438:10'b0);
   assign  _add_map_x_190_sg_up = ((_net_7618)?sg_in438:2'b0)|
    ((_net_3626)?sg_in437:2'b0);
   assign  _add_map_x_190_sg_down = ((_net_7617)?sg_in405:2'b0)|
    ((_net_3625)?sg_in439:2'b0);
   assign  _add_map_x_190_sg_left = ((_net_7615)?sg_in469:2'b0)|
    ((_net_3623)?sg_in470:2'b0);
   assign  _add_map_x_190_sg_right = ((_net_7616)?sg_in436:2'b0)|
    ((_net_3624)?sg_in406:2'b0);
   assign  _add_map_x_190_wall_t_in = dig_w;
   assign  _add_map_x_190_moto = ((_net_7613)?data_in437:10'b0)|
    ((_net_3621)?data_in438:10'b0);
   assign  _add_map_x_190_up = ((_net_7612)?data_in438:10'b0)|
    ((_net_3620)?data_in437:10'b0);
   assign  _add_map_x_190_right = ((_net_7611)?data_in436:10'b0)|
    ((_net_3619)?data_in439:10'b0);
   assign  _add_map_x_190_down = ((_net_7610)?data_in405:10'b0)|
    ((_net_3618)?data_in406:10'b0);
   assign  _add_map_x_190_left = ((_net_7609)?data_in469:10'b0)|
    ((_net_3617)?data_in470:10'b0);
   assign  _add_map_x_190_start = start;
   assign  _add_map_x_190_goal = goal;
   assign  _add_map_x_190_now = ((_net_7606)?10'b0110110101:10'b0)|
    ((_net_3614)?10'b0110110110:10'b0);
   assign  _add_map_x_190_add_exe = (_net_7605|_net_3613);
   assign  _add_map_x_190_p_reset = p_reset;
   assign  _add_map_x_190_m_clock = m_clock;
   assign  _add_map_x_189_moto_org_near = ((_net_7604)?data_in_org436:10'b0)|
    ((_net_3612)?data_in_org435:10'b0);
   assign  _add_map_x_189_moto_org_near1 = ((_net_7603)?data_in_org434:10'b0)|
    ((_net_3611)?data_in_org437:10'b0);
   assign  _add_map_x_189_moto_org_near2 = ((_net_7602)?data_in_org403:10'b0)|
    ((_net_3610)?data_in_org404:10'b0);
   assign  _add_map_x_189_moto_org_near3 = ((_net_7601)?data_in_org467:10'b0)|
    ((_net_3609)?data_in_org468:10'b0);
   assign  _add_map_x_189_moto_org = ((_net_7600)?data_in_org435:10'b0)|
    ((_net_3608)?data_in_org436:10'b0);
   assign  _add_map_x_189_sg_up = ((_net_7599)?sg_in436:2'b0)|
    ((_net_3607)?sg_in435:2'b0);
   assign  _add_map_x_189_sg_down = ((_net_7598)?sg_in403:2'b0)|
    ((_net_3606)?sg_in437:2'b0);
   assign  _add_map_x_189_sg_left = ((_net_7596)?sg_in467:2'b0)|
    ((_net_3604)?sg_in468:2'b0);
   assign  _add_map_x_189_sg_right = ((_net_7597)?sg_in434:2'b0)|
    ((_net_3605)?sg_in404:2'b0);
   assign  _add_map_x_189_wall_t_in = dig_w;
   assign  _add_map_x_189_moto = ((_net_7594)?data_in435:10'b0)|
    ((_net_3602)?data_in436:10'b0);
   assign  _add_map_x_189_up = ((_net_7593)?data_in436:10'b0)|
    ((_net_3601)?data_in435:10'b0);
   assign  _add_map_x_189_right = ((_net_7592)?data_in434:10'b0)|
    ((_net_3600)?data_in437:10'b0);
   assign  _add_map_x_189_down = ((_net_7591)?data_in403:10'b0)|
    ((_net_3599)?data_in404:10'b0);
   assign  _add_map_x_189_left = ((_net_7590)?data_in467:10'b0)|
    ((_net_3598)?data_in468:10'b0);
   assign  _add_map_x_189_start = start;
   assign  _add_map_x_189_goal = goal;
   assign  _add_map_x_189_now = ((_net_7587)?10'b0110110011:10'b0)|
    ((_net_3595)?10'b0110110100:10'b0);
   assign  _add_map_x_189_add_exe = (_net_7586|_net_3594);
   assign  _add_map_x_189_p_reset = p_reset;
   assign  _add_map_x_189_m_clock = m_clock;
   assign  _add_map_x_188_moto_org_near = ((_net_7585)?data_in_org434:10'b0)|
    ((_net_3593)?data_in_org433:10'b0);
   assign  _add_map_x_188_moto_org_near1 = ((_net_7584)?data_in_org432:10'b0)|
    ((_net_3592)?data_in_org435:10'b0);
   assign  _add_map_x_188_moto_org_near2 = ((_net_7583)?data_in_org401:10'b0)|
    ((_net_3591)?data_in_org402:10'b0);
   assign  _add_map_x_188_moto_org_near3 = ((_net_7582)?data_in_org465:10'b0)|
    ((_net_3590)?data_in_org466:10'b0);
   assign  _add_map_x_188_moto_org = ((_net_7581)?data_in_org433:10'b0)|
    ((_net_3589)?data_in_org434:10'b0);
   assign  _add_map_x_188_sg_up = ((_net_7580)?sg_in434:2'b0)|
    ((_net_3588)?sg_in433:2'b0);
   assign  _add_map_x_188_sg_down = ((_net_7579)?sg_in401:2'b0)|
    ((_net_3587)?sg_in435:2'b0);
   assign  _add_map_x_188_sg_left = ((_net_7577)?sg_in465:2'b0)|
    ((_net_3585)?sg_in466:2'b0);
   assign  _add_map_x_188_sg_right = ((_net_7578)?sg_in432:2'b0)|
    ((_net_3586)?sg_in402:2'b0);
   assign  _add_map_x_188_wall_t_in = dig_w;
   assign  _add_map_x_188_moto = ((_net_7575)?data_in433:10'b0)|
    ((_net_3583)?data_in434:10'b0);
   assign  _add_map_x_188_up = ((_net_7574)?data_in434:10'b0)|
    ((_net_3582)?data_in433:10'b0);
   assign  _add_map_x_188_right = ((_net_7573)?data_in432:10'b0)|
    ((_net_3581)?data_in435:10'b0);
   assign  _add_map_x_188_down = ((_net_7572)?data_in401:10'b0)|
    ((_net_3580)?data_in402:10'b0);
   assign  _add_map_x_188_left = ((_net_7571)?data_in465:10'b0)|
    ((_net_3579)?data_in466:10'b0);
   assign  _add_map_x_188_start = start;
   assign  _add_map_x_188_goal = goal;
   assign  _add_map_x_188_now = ((_net_7568)?10'b0110110001:10'b0)|
    ((_net_3576)?10'b0110110010:10'b0);
   assign  _add_map_x_188_add_exe = (_net_7567|_net_3575);
   assign  _add_map_x_188_p_reset = p_reset;
   assign  _add_map_x_188_m_clock = m_clock;
   assign  _add_map_x_187_moto_org_near = ((_net_7566)?data_in_org432:10'b0)|
    ((_net_3574)?data_in_org431:10'b0);
   assign  _add_map_x_187_moto_org_near1 = ((_net_7565)?data_in_org430:10'b0)|
    ((_net_3573)?data_in_org433:10'b0);
   assign  _add_map_x_187_moto_org_near2 = ((_net_7564)?data_in_org399:10'b0)|
    ((_net_3572)?data_in_org400:10'b0);
   assign  _add_map_x_187_moto_org_near3 = ((_net_7563)?data_in_org463:10'b0)|
    ((_net_3571)?data_in_org464:10'b0);
   assign  _add_map_x_187_moto_org = ((_net_7562)?data_in_org431:10'b0)|
    ((_net_3570)?data_in_org432:10'b0);
   assign  _add_map_x_187_sg_up = ((_net_7561)?sg_in432:2'b0)|
    ((_net_3569)?sg_in431:2'b0);
   assign  _add_map_x_187_sg_down = ((_net_7560)?sg_in399:2'b0)|
    ((_net_3568)?sg_in433:2'b0);
   assign  _add_map_x_187_sg_left = ((_net_7558)?sg_in463:2'b0)|
    ((_net_3566)?sg_in464:2'b0);
   assign  _add_map_x_187_sg_right = ((_net_7559)?sg_in430:2'b0)|
    ((_net_3567)?sg_in400:2'b0);
   assign  _add_map_x_187_wall_t_in = dig_w;
   assign  _add_map_x_187_moto = ((_net_7556)?data_in431:10'b0)|
    ((_net_3564)?data_in432:10'b0);
   assign  _add_map_x_187_up = ((_net_7555)?data_in432:10'b0)|
    ((_net_3563)?data_in431:10'b0);
   assign  _add_map_x_187_right = ((_net_7554)?data_in430:10'b0)|
    ((_net_3562)?data_in433:10'b0);
   assign  _add_map_x_187_down = ((_net_7553)?data_in399:10'b0)|
    ((_net_3561)?data_in400:10'b0);
   assign  _add_map_x_187_left = ((_net_7552)?data_in463:10'b0)|
    ((_net_3560)?data_in464:10'b0);
   assign  _add_map_x_187_start = start;
   assign  _add_map_x_187_goal = goal;
   assign  _add_map_x_187_now = ((_net_7549)?10'b0110101111:10'b0)|
    ((_net_3557)?10'b0110110000:10'b0);
   assign  _add_map_x_187_add_exe = (_net_7548|_net_3556);
   assign  _add_map_x_187_p_reset = p_reset;
   assign  _add_map_x_187_m_clock = m_clock;
   assign  _add_map_x_186_moto_org_near = ((_net_7547)?data_in_org430:10'b0)|
    ((_net_3555)?data_in_org429:10'b0);
   assign  _add_map_x_186_moto_org_near1 = ((_net_7546)?data_in_org428:10'b0)|
    ((_net_3554)?data_in_org431:10'b0);
   assign  _add_map_x_186_moto_org_near2 = ((_net_7545)?data_in_org397:10'b0)|
    ((_net_3553)?data_in_org398:10'b0);
   assign  _add_map_x_186_moto_org_near3 = ((_net_7544)?data_in_org461:10'b0)|
    ((_net_3552)?data_in_org462:10'b0);
   assign  _add_map_x_186_moto_org = ((_net_7543)?data_in_org429:10'b0)|
    ((_net_3551)?data_in_org430:10'b0);
   assign  _add_map_x_186_sg_up = ((_net_7542)?sg_in430:2'b0)|
    ((_net_3550)?sg_in429:2'b0);
   assign  _add_map_x_186_sg_down = ((_net_7541)?sg_in397:2'b0)|
    ((_net_3549)?sg_in431:2'b0);
   assign  _add_map_x_186_sg_left = ((_net_7539)?sg_in461:2'b0)|
    ((_net_3547)?sg_in462:2'b0);
   assign  _add_map_x_186_sg_right = ((_net_7540)?sg_in428:2'b0)|
    ((_net_3548)?sg_in398:2'b0);
   assign  _add_map_x_186_wall_t_in = dig_w;
   assign  _add_map_x_186_moto = ((_net_7537)?data_in429:10'b0)|
    ((_net_3545)?data_in430:10'b0);
   assign  _add_map_x_186_up = ((_net_7536)?data_in430:10'b0)|
    ((_net_3544)?data_in429:10'b0);
   assign  _add_map_x_186_right = ((_net_7535)?data_in428:10'b0)|
    ((_net_3543)?data_in431:10'b0);
   assign  _add_map_x_186_down = ((_net_7534)?data_in397:10'b0)|
    ((_net_3542)?data_in398:10'b0);
   assign  _add_map_x_186_left = ((_net_7533)?data_in461:10'b0)|
    ((_net_3541)?data_in462:10'b0);
   assign  _add_map_x_186_start = start;
   assign  _add_map_x_186_goal = goal;
   assign  _add_map_x_186_now = ((_net_7530)?10'b0110101101:10'b0)|
    ((_net_3538)?10'b0110101110:10'b0);
   assign  _add_map_x_186_add_exe = (_net_7529|_net_3537);
   assign  _add_map_x_186_p_reset = p_reset;
   assign  _add_map_x_186_m_clock = m_clock;
   assign  _add_map_x_185_moto_org_near = ((_net_7528)?data_in_org428:10'b0)|
    ((_net_3536)?data_in_org427:10'b0);
   assign  _add_map_x_185_moto_org_near1 = ((_net_7527)?data_in_org426:10'b0)|
    ((_net_3535)?data_in_org429:10'b0);
   assign  _add_map_x_185_moto_org_near2 = ((_net_7526)?data_in_org395:10'b0)|
    ((_net_3534)?data_in_org396:10'b0);
   assign  _add_map_x_185_moto_org_near3 = ((_net_7525)?data_in_org459:10'b0)|
    ((_net_3533)?data_in_org460:10'b0);
   assign  _add_map_x_185_moto_org = ((_net_7524)?data_in_org427:10'b0)|
    ((_net_3532)?data_in_org428:10'b0);
   assign  _add_map_x_185_sg_up = ((_net_7523)?sg_in428:2'b0)|
    ((_net_3531)?sg_in427:2'b0);
   assign  _add_map_x_185_sg_down = ((_net_7522)?sg_in395:2'b0)|
    ((_net_3530)?sg_in429:2'b0);
   assign  _add_map_x_185_sg_left = ((_net_7520)?sg_in459:2'b0)|
    ((_net_3528)?sg_in460:2'b0);
   assign  _add_map_x_185_sg_right = ((_net_7521)?sg_in426:2'b0)|
    ((_net_3529)?sg_in396:2'b0);
   assign  _add_map_x_185_wall_t_in = dig_w;
   assign  _add_map_x_185_moto = ((_net_7518)?data_in427:10'b0)|
    ((_net_3526)?data_in428:10'b0);
   assign  _add_map_x_185_up = ((_net_7517)?data_in428:10'b0)|
    ((_net_3525)?data_in427:10'b0);
   assign  _add_map_x_185_right = ((_net_7516)?data_in426:10'b0)|
    ((_net_3524)?data_in429:10'b0);
   assign  _add_map_x_185_down = ((_net_7515)?data_in395:10'b0)|
    ((_net_3523)?data_in396:10'b0);
   assign  _add_map_x_185_left = ((_net_7514)?data_in459:10'b0)|
    ((_net_3522)?data_in460:10'b0);
   assign  _add_map_x_185_start = start;
   assign  _add_map_x_185_goal = goal;
   assign  _add_map_x_185_now = ((_net_7511)?10'b0110101011:10'b0)|
    ((_net_3519)?10'b0110101100:10'b0);
   assign  _add_map_x_185_add_exe = (_net_7510|_net_3518);
   assign  _add_map_x_185_p_reset = p_reset;
   assign  _add_map_x_185_m_clock = m_clock;
   assign  _add_map_x_184_moto_org_near = ((_net_7509)?data_in_org426:10'b0)|
    ((_net_3517)?data_in_org425:10'b0);
   assign  _add_map_x_184_moto_org_near1 = ((_net_7508)?data_in_org424:10'b0)|
    ((_net_3516)?data_in_org427:10'b0);
   assign  _add_map_x_184_moto_org_near2 = ((_net_7507)?data_in_org393:10'b0)|
    ((_net_3515)?data_in_org394:10'b0);
   assign  _add_map_x_184_moto_org_near3 = ((_net_7506)?data_in_org457:10'b0)|
    ((_net_3514)?data_in_org458:10'b0);
   assign  _add_map_x_184_moto_org = ((_net_7505)?data_in_org425:10'b0)|
    ((_net_3513)?data_in_org426:10'b0);
   assign  _add_map_x_184_sg_up = ((_net_7504)?sg_in426:2'b0)|
    ((_net_3512)?sg_in425:2'b0);
   assign  _add_map_x_184_sg_down = ((_net_7503)?sg_in393:2'b0)|
    ((_net_3511)?sg_in427:2'b0);
   assign  _add_map_x_184_sg_left = ((_net_7501)?sg_in457:2'b0)|
    ((_net_3509)?sg_in458:2'b0);
   assign  _add_map_x_184_sg_right = ((_net_7502)?sg_in424:2'b0)|
    ((_net_3510)?sg_in394:2'b0);
   assign  _add_map_x_184_wall_t_in = dig_w;
   assign  _add_map_x_184_moto = ((_net_7499)?data_in425:10'b0)|
    ((_net_3507)?data_in426:10'b0);
   assign  _add_map_x_184_up = ((_net_7498)?data_in426:10'b0)|
    ((_net_3506)?data_in425:10'b0);
   assign  _add_map_x_184_right = ((_net_7497)?data_in424:10'b0)|
    ((_net_3505)?data_in427:10'b0);
   assign  _add_map_x_184_down = ((_net_7496)?data_in393:10'b0)|
    ((_net_3504)?data_in394:10'b0);
   assign  _add_map_x_184_left = ((_net_7495)?data_in457:10'b0)|
    ((_net_3503)?data_in458:10'b0);
   assign  _add_map_x_184_start = start;
   assign  _add_map_x_184_goal = goal;
   assign  _add_map_x_184_now = ((_net_7492)?10'b0110101001:10'b0)|
    ((_net_3500)?10'b0110101010:10'b0);
   assign  _add_map_x_184_add_exe = (_net_7491|_net_3499);
   assign  _add_map_x_184_p_reset = p_reset;
   assign  _add_map_x_184_m_clock = m_clock;
   assign  _add_map_x_183_moto_org_near = ((_net_7490)?data_in_org424:10'b0)|
    ((_net_3498)?data_in_org423:10'b0);
   assign  _add_map_x_183_moto_org_near1 = ((_net_7489)?data_in_org422:10'b0)|
    ((_net_3497)?data_in_org425:10'b0);
   assign  _add_map_x_183_moto_org_near2 = ((_net_7488)?data_in_org391:10'b0)|
    ((_net_3496)?data_in_org392:10'b0);
   assign  _add_map_x_183_moto_org_near3 = ((_net_7487)?data_in_org455:10'b0)|
    ((_net_3495)?data_in_org456:10'b0);
   assign  _add_map_x_183_moto_org = ((_net_7486)?data_in_org423:10'b0)|
    ((_net_3494)?data_in_org424:10'b0);
   assign  _add_map_x_183_sg_up = ((_net_7485)?sg_in424:2'b0)|
    ((_net_3493)?sg_in423:2'b0);
   assign  _add_map_x_183_sg_down = ((_net_7484)?sg_in391:2'b0)|
    ((_net_3492)?sg_in425:2'b0);
   assign  _add_map_x_183_sg_left = ((_net_7482)?sg_in455:2'b0)|
    ((_net_3490)?sg_in456:2'b0);
   assign  _add_map_x_183_sg_right = ((_net_7483)?sg_in422:2'b0)|
    ((_net_3491)?sg_in392:2'b0);
   assign  _add_map_x_183_wall_t_in = dig_w;
   assign  _add_map_x_183_moto = ((_net_7480)?data_in423:10'b0)|
    ((_net_3488)?data_in424:10'b0);
   assign  _add_map_x_183_up = ((_net_7479)?data_in424:10'b0)|
    ((_net_3487)?data_in423:10'b0);
   assign  _add_map_x_183_right = ((_net_7478)?data_in422:10'b0)|
    ((_net_3486)?data_in425:10'b0);
   assign  _add_map_x_183_down = ((_net_7477)?data_in391:10'b0)|
    ((_net_3485)?data_in392:10'b0);
   assign  _add_map_x_183_left = ((_net_7476)?data_in455:10'b0)|
    ((_net_3484)?data_in456:10'b0);
   assign  _add_map_x_183_start = start;
   assign  _add_map_x_183_goal = goal;
   assign  _add_map_x_183_now = ((_net_7473)?10'b0110100111:10'b0)|
    ((_net_3481)?10'b0110101000:10'b0);
   assign  _add_map_x_183_add_exe = (_net_7472|_net_3480);
   assign  _add_map_x_183_p_reset = p_reset;
   assign  _add_map_x_183_m_clock = m_clock;
   assign  _add_map_x_182_moto_org_near = ((_net_7471)?data_in_org422:10'b0)|
    ((_net_3479)?data_in_org421:10'b0);
   assign  _add_map_x_182_moto_org_near1 = ((_net_7470)?data_in_org420:10'b0)|
    ((_net_3478)?data_in_org423:10'b0);
   assign  _add_map_x_182_moto_org_near2 = ((_net_7469)?data_in_org389:10'b0)|
    ((_net_3477)?data_in_org390:10'b0);
   assign  _add_map_x_182_moto_org_near3 = ((_net_7468)?data_in_org453:10'b0)|
    ((_net_3476)?data_in_org454:10'b0);
   assign  _add_map_x_182_moto_org = ((_net_7467)?data_in_org421:10'b0)|
    ((_net_3475)?data_in_org422:10'b0);
   assign  _add_map_x_182_sg_up = ((_net_7466)?sg_in422:2'b0)|
    ((_net_3474)?sg_in421:2'b0);
   assign  _add_map_x_182_sg_down = ((_net_7465)?sg_in389:2'b0)|
    ((_net_3473)?sg_in423:2'b0);
   assign  _add_map_x_182_sg_left = ((_net_7463)?sg_in453:2'b0)|
    ((_net_3471)?sg_in454:2'b0);
   assign  _add_map_x_182_sg_right = ((_net_7464)?sg_in420:2'b0)|
    ((_net_3472)?sg_in390:2'b0);
   assign  _add_map_x_182_wall_t_in = dig_w;
   assign  _add_map_x_182_moto = ((_net_7461)?data_in421:10'b0)|
    ((_net_3469)?data_in422:10'b0);
   assign  _add_map_x_182_up = ((_net_7460)?data_in422:10'b0)|
    ((_net_3468)?data_in421:10'b0);
   assign  _add_map_x_182_right = ((_net_7459)?data_in420:10'b0)|
    ((_net_3467)?data_in423:10'b0);
   assign  _add_map_x_182_down = ((_net_7458)?data_in389:10'b0)|
    ((_net_3466)?data_in390:10'b0);
   assign  _add_map_x_182_left = ((_net_7457)?data_in453:10'b0)|
    ((_net_3465)?data_in454:10'b0);
   assign  _add_map_x_182_start = start;
   assign  _add_map_x_182_goal = goal;
   assign  _add_map_x_182_now = ((_net_7454)?10'b0110100101:10'b0)|
    ((_net_3462)?10'b0110100110:10'b0);
   assign  _add_map_x_182_add_exe = (_net_7453|_net_3461);
   assign  _add_map_x_182_p_reset = p_reset;
   assign  _add_map_x_182_m_clock = m_clock;
   assign  _add_map_x_181_moto_org_near = ((_net_7452)?data_in_org420:10'b0)|
    ((_net_3460)?data_in_org419:10'b0);
   assign  _add_map_x_181_moto_org_near1 = ((_net_7451)?data_in_org418:10'b0)|
    ((_net_3459)?data_in_org421:10'b0);
   assign  _add_map_x_181_moto_org_near2 = ((_net_7450)?data_in_org387:10'b0)|
    ((_net_3458)?data_in_org388:10'b0);
   assign  _add_map_x_181_moto_org_near3 = ((_net_7449)?data_in_org451:10'b0)|
    ((_net_3457)?data_in_org452:10'b0);
   assign  _add_map_x_181_moto_org = ((_net_7448)?data_in_org419:10'b0)|
    ((_net_3456)?data_in_org420:10'b0);
   assign  _add_map_x_181_sg_up = ((_net_7447)?sg_in420:2'b0)|
    ((_net_3455)?sg_in419:2'b0);
   assign  _add_map_x_181_sg_down = ((_net_7446)?sg_in387:2'b0)|
    ((_net_3454)?sg_in421:2'b0);
   assign  _add_map_x_181_sg_left = ((_net_7444)?sg_in451:2'b0)|
    ((_net_3452)?sg_in452:2'b0);
   assign  _add_map_x_181_sg_right = ((_net_7445)?sg_in418:2'b0)|
    ((_net_3453)?sg_in388:2'b0);
   assign  _add_map_x_181_wall_t_in = dig_w;
   assign  _add_map_x_181_moto = ((_net_7442)?data_in419:10'b0)|
    ((_net_3450)?data_in420:10'b0);
   assign  _add_map_x_181_up = ((_net_7441)?data_in420:10'b0)|
    ((_net_3449)?data_in419:10'b0);
   assign  _add_map_x_181_right = ((_net_7440)?data_in418:10'b0)|
    ((_net_3448)?data_in421:10'b0);
   assign  _add_map_x_181_down = ((_net_7439)?data_in387:10'b0)|
    ((_net_3447)?data_in388:10'b0);
   assign  _add_map_x_181_left = ((_net_7438)?data_in451:10'b0)|
    ((_net_3446)?data_in452:10'b0);
   assign  _add_map_x_181_start = start;
   assign  _add_map_x_181_goal = goal;
   assign  _add_map_x_181_now = ((_net_7435)?10'b0110100011:10'b0)|
    ((_net_3443)?10'b0110100100:10'b0);
   assign  _add_map_x_181_add_exe = (_net_7434|_net_3442);
   assign  _add_map_x_181_p_reset = p_reset;
   assign  _add_map_x_181_m_clock = m_clock;
   assign  _add_map_x_180_moto_org_near = ((_net_7433)?data_in_org418:10'b0)|
    ((_net_3441)?data_in_org417:10'b0);
   assign  _add_map_x_180_moto_org_near1 = ((_net_7432)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_3440)?data_in_org419:10'b0);
   assign  _add_map_x_180_moto_org_near2 = ((_net_7431)?data_in_org385:10'b0)|
    ((_net_3439)?data_in_org386:10'b0);
   assign  _add_map_x_180_moto_org_near3 = ((_net_7430)?data_in_org449:10'b0)|
    ((_net_3438)?data_in_org450:10'b0);
   assign  _add_map_x_180_moto_org = ((_net_7429)?data_in_org417:10'b0)|
    ((_net_3437)?data_in_org418:10'b0);
   assign  _add_map_x_180_sg_up = ((_net_7428)?sg_in418:2'b0)|
    ((_net_3436)?sg_in417:2'b0);
   assign  _add_map_x_180_sg_down = ((_net_7427)?sg_in385:2'b0)|
    ((_net_3435)?sg_in419:2'b0);
   assign  _add_map_x_180_sg_left = ((_net_7425)?sg_in449:2'b0)|
    ((_net_3433)?sg_in450:2'b0);
   assign  _add_map_x_180_sg_right = ((_net_7426)?3'b000:2'b0)|
    ((_net_3434)?sg_in386:2'b0);
   assign  _add_map_x_180_wall_t_in = dig_w;
   assign  _add_map_x_180_moto = ((_net_7423)?data_in417:10'b0)|
    ((_net_3431)?data_in418:10'b0);
   assign  _add_map_x_180_up = ((_net_7422)?data_in418:10'b0)|
    ((_net_3430)?data_in417:10'b0);
   assign  _add_map_x_180_right = ((_net_7421)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_3429)?data_in419:10'b0);
   assign  _add_map_x_180_down = ((_net_7420)?data_in385:10'b0)|
    ((_net_3428)?data_in386:10'b0);
   assign  _add_map_x_180_left = ((_net_7419)?data_in449:10'b0)|
    ((_net_3427)?data_in450:10'b0);
   assign  _add_map_x_180_start = start;
   assign  _add_map_x_180_goal = goal;
   assign  _add_map_x_180_now = ((_net_7416)?10'b0110100001:10'b0)|
    ((_net_3424)?10'b0110100010:10'b0);
   assign  _add_map_x_180_add_exe = (_net_7415|_net_3423);
   assign  _add_map_x_180_p_reset = p_reset;
   assign  _add_map_x_180_m_clock = m_clock;
   assign  _add_map_x_179_moto_org_near = ((_net_7414)?data_in_org413:10'b0)|
    ((_net_3422)?data_in_org414:10'b0);
   assign  _add_map_x_179_moto_org_near1 = ((_net_7413)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_3421)?data_in_org412:10'b0);
   assign  _add_map_x_179_moto_org_near2 = ((_net_7412)?data_in_org382:10'b0)|
    ((_net_3420)?data_in_org381:10'b0);
   assign  _add_map_x_179_moto_org_near3 = ((_net_7411)?data_in_org446:10'b0)|
    ((_net_3419)?data_in_org445:10'b0);
   assign  _add_map_x_179_moto_org = ((_net_7410)?data_in_org414:10'b0)|
    ((_net_3418)?data_in_org413:10'b0);
   assign  _add_map_x_179_sg_up = ((_net_7409)?sg_in413:2'b0)|
    ((_net_3417)?sg_in414:2'b0);
   assign  _add_map_x_179_sg_down = ((_net_7408)?3'b000:2'b0)|
    ((_net_3416)?sg_in412:2'b0);
   assign  _add_map_x_179_sg_left = ((_net_7406)?sg_in446:2'b0)|
    ((_net_3414)?sg_in445:2'b0);
   assign  _add_map_x_179_sg_right = ((_net_7407)?sg_in382:2'b0)|
    ((_net_3415)?sg_in381:2'b0);
   assign  _add_map_x_179_wall_t_in = dig_w;
   assign  _add_map_x_179_moto = ((_net_7404)?data_in414:10'b0)|
    ((_net_3412)?data_in413:10'b0);
   assign  _add_map_x_179_up = ((_net_7403)?data_in413:10'b0)|
    ((_net_3411)?data_in414:10'b0);
   assign  _add_map_x_179_right = ((_net_7402)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_3410)?data_in412:10'b0);
   assign  _add_map_x_179_down = ((_net_7401)?data_in382:10'b0)|
    ((_net_3409)?data_in381:10'b0);
   assign  _add_map_x_179_left = ((_net_7400)?data_in446:10'b0)|
    ((_net_3408)?data_in445:10'b0);
   assign  _add_map_x_179_start = start;
   assign  _add_map_x_179_goal = goal;
   assign  _add_map_x_179_now = ((_net_7397)?10'b0110011110:10'b0)|
    ((_net_3405)?10'b0110011101:10'b0);
   assign  _add_map_x_179_add_exe = (_net_7396|_net_3404);
   assign  _add_map_x_179_p_reset = p_reset;
   assign  _add_map_x_179_m_clock = m_clock;
   assign  _add_map_x_178_moto_org_near = ((_net_7395)?data_in_org411:10'b0)|
    ((_net_3403)?data_in_org412:10'b0);
   assign  _add_map_x_178_moto_org_near1 = ((_net_7394)?data_in_org413:10'b0)|
    ((_net_3402)?data_in_org410:10'b0);
   assign  _add_map_x_178_moto_org_near2 = ((_net_7393)?data_in_org380:10'b0)|
    ((_net_3401)?data_in_org379:10'b0);
   assign  _add_map_x_178_moto_org_near3 = ((_net_7392)?data_in_org444:10'b0)|
    ((_net_3400)?data_in_org443:10'b0);
   assign  _add_map_x_178_moto_org = ((_net_7391)?data_in_org412:10'b0)|
    ((_net_3399)?data_in_org411:10'b0);
   assign  _add_map_x_178_sg_up = ((_net_7390)?sg_in411:2'b0)|
    ((_net_3398)?sg_in412:2'b0);
   assign  _add_map_x_178_sg_down = ((_net_7389)?sg_in413:2'b0)|
    ((_net_3397)?sg_in410:2'b0);
   assign  _add_map_x_178_sg_left = ((_net_7387)?sg_in444:2'b0)|
    ((_net_3395)?sg_in443:2'b0);
   assign  _add_map_x_178_sg_right = ((_net_7388)?sg_in380:2'b0)|
    ((_net_3396)?sg_in379:2'b0);
   assign  _add_map_x_178_wall_t_in = dig_w;
   assign  _add_map_x_178_moto = ((_net_7385)?data_in412:10'b0)|
    ((_net_3393)?data_in411:10'b0);
   assign  _add_map_x_178_up = ((_net_7384)?data_in411:10'b0)|
    ((_net_3392)?data_in412:10'b0);
   assign  _add_map_x_178_right = ((_net_7383)?data_in413:10'b0)|
    ((_net_3391)?data_in410:10'b0);
   assign  _add_map_x_178_down = ((_net_7382)?data_in380:10'b0)|
    ((_net_3390)?data_in379:10'b0);
   assign  _add_map_x_178_left = ((_net_7381)?data_in444:10'b0)|
    ((_net_3389)?data_in443:10'b0);
   assign  _add_map_x_178_start = start;
   assign  _add_map_x_178_goal = goal;
   assign  _add_map_x_178_now = ((_net_7378)?10'b0110011100:10'b0)|
    ((_net_3386)?10'b0110011011:10'b0);
   assign  _add_map_x_178_add_exe = (_net_7377|_net_3385);
   assign  _add_map_x_178_p_reset = p_reset;
   assign  _add_map_x_178_m_clock = m_clock;
   assign  _add_map_x_177_moto_org_near = ((_net_7376)?data_in_org409:10'b0)|
    ((_net_3384)?data_in_org410:10'b0);
   assign  _add_map_x_177_moto_org_near1 = ((_net_7375)?data_in_org411:10'b0)|
    ((_net_3383)?data_in_org408:10'b0);
   assign  _add_map_x_177_moto_org_near2 = ((_net_7374)?data_in_org378:10'b0)|
    ((_net_3382)?data_in_org377:10'b0);
   assign  _add_map_x_177_moto_org_near3 = ((_net_7373)?data_in_org442:10'b0)|
    ((_net_3381)?data_in_org441:10'b0);
   assign  _add_map_x_177_moto_org = ((_net_7372)?data_in_org410:10'b0)|
    ((_net_3380)?data_in_org409:10'b0);
   assign  _add_map_x_177_sg_up = ((_net_7371)?sg_in409:2'b0)|
    ((_net_3379)?sg_in410:2'b0);
   assign  _add_map_x_177_sg_down = ((_net_7370)?sg_in411:2'b0)|
    ((_net_3378)?sg_in408:2'b0);
   assign  _add_map_x_177_sg_left = ((_net_7368)?sg_in442:2'b0)|
    ((_net_3376)?sg_in441:2'b0);
   assign  _add_map_x_177_sg_right = ((_net_7369)?sg_in378:2'b0)|
    ((_net_3377)?sg_in377:2'b0);
   assign  _add_map_x_177_wall_t_in = dig_w;
   assign  _add_map_x_177_moto = ((_net_7366)?data_in410:10'b0)|
    ((_net_3374)?data_in409:10'b0);
   assign  _add_map_x_177_up = ((_net_7365)?data_in409:10'b0)|
    ((_net_3373)?data_in410:10'b0);
   assign  _add_map_x_177_right = ((_net_7364)?data_in411:10'b0)|
    ((_net_3372)?data_in408:10'b0);
   assign  _add_map_x_177_down = ((_net_7363)?data_in378:10'b0)|
    ((_net_3371)?data_in377:10'b0);
   assign  _add_map_x_177_left = ((_net_7362)?data_in442:10'b0)|
    ((_net_3370)?data_in441:10'b0);
   assign  _add_map_x_177_start = start;
   assign  _add_map_x_177_goal = goal;
   assign  _add_map_x_177_now = ((_net_7359)?10'b0110011010:10'b0)|
    ((_net_3367)?10'b0110011001:10'b0);
   assign  _add_map_x_177_add_exe = (_net_7358|_net_3366);
   assign  _add_map_x_177_p_reset = p_reset;
   assign  _add_map_x_177_m_clock = m_clock;
   assign  _add_map_x_176_moto_org_near = ((_net_7357)?data_in_org407:10'b0)|
    ((_net_3365)?data_in_org408:10'b0);
   assign  _add_map_x_176_moto_org_near1 = ((_net_7356)?data_in_org409:10'b0)|
    ((_net_3364)?data_in_org406:10'b0);
   assign  _add_map_x_176_moto_org_near2 = ((_net_7355)?data_in_org376:10'b0)|
    ((_net_3363)?data_in_org375:10'b0);
   assign  _add_map_x_176_moto_org_near3 = ((_net_7354)?data_in_org440:10'b0)|
    ((_net_3362)?data_in_org439:10'b0);
   assign  _add_map_x_176_moto_org = ((_net_7353)?data_in_org408:10'b0)|
    ((_net_3361)?data_in_org407:10'b0);
   assign  _add_map_x_176_sg_up = ((_net_7352)?sg_in407:2'b0)|
    ((_net_3360)?sg_in408:2'b0);
   assign  _add_map_x_176_sg_down = ((_net_7351)?sg_in409:2'b0)|
    ((_net_3359)?sg_in406:2'b0);
   assign  _add_map_x_176_sg_left = ((_net_7349)?sg_in440:2'b0)|
    ((_net_3357)?sg_in439:2'b0);
   assign  _add_map_x_176_sg_right = ((_net_7350)?sg_in376:2'b0)|
    ((_net_3358)?sg_in375:2'b0);
   assign  _add_map_x_176_wall_t_in = dig_w;
   assign  _add_map_x_176_moto = ((_net_7347)?data_in408:10'b0)|
    ((_net_3355)?data_in407:10'b0);
   assign  _add_map_x_176_up = ((_net_7346)?data_in407:10'b0)|
    ((_net_3354)?data_in408:10'b0);
   assign  _add_map_x_176_right = ((_net_7345)?data_in409:10'b0)|
    ((_net_3353)?data_in406:10'b0);
   assign  _add_map_x_176_down = ((_net_7344)?data_in376:10'b0)|
    ((_net_3352)?data_in375:10'b0);
   assign  _add_map_x_176_left = ((_net_7343)?data_in440:10'b0)|
    ((_net_3351)?data_in439:10'b0);
   assign  _add_map_x_176_start = start;
   assign  _add_map_x_176_goal = goal;
   assign  _add_map_x_176_now = ((_net_7340)?10'b0110011000:10'b0)|
    ((_net_3348)?10'b0110010111:10'b0);
   assign  _add_map_x_176_add_exe = (_net_7339|_net_3347);
   assign  _add_map_x_176_p_reset = p_reset;
   assign  _add_map_x_176_m_clock = m_clock;
   assign  _add_map_x_175_moto_org_near = ((_net_7338)?data_in_org405:10'b0)|
    ((_net_3346)?data_in_org406:10'b0);
   assign  _add_map_x_175_moto_org_near1 = ((_net_7337)?data_in_org407:10'b0)|
    ((_net_3345)?data_in_org404:10'b0);
   assign  _add_map_x_175_moto_org_near2 = ((_net_7336)?data_in_org374:10'b0)|
    ((_net_3344)?data_in_org373:10'b0);
   assign  _add_map_x_175_moto_org_near3 = ((_net_7335)?data_in_org438:10'b0)|
    ((_net_3343)?data_in_org437:10'b0);
   assign  _add_map_x_175_moto_org = ((_net_7334)?data_in_org406:10'b0)|
    ((_net_3342)?data_in_org405:10'b0);
   assign  _add_map_x_175_sg_up = ((_net_7333)?sg_in405:2'b0)|
    ((_net_3341)?sg_in406:2'b0);
   assign  _add_map_x_175_sg_down = ((_net_7332)?sg_in407:2'b0)|
    ((_net_3340)?sg_in404:2'b0);
   assign  _add_map_x_175_sg_left = ((_net_7330)?sg_in438:2'b0)|
    ((_net_3338)?sg_in437:2'b0);
   assign  _add_map_x_175_sg_right = ((_net_7331)?sg_in374:2'b0)|
    ((_net_3339)?sg_in373:2'b0);
   assign  _add_map_x_175_wall_t_in = dig_w;
   assign  _add_map_x_175_moto = ((_net_7328)?data_in406:10'b0)|
    ((_net_3336)?data_in405:10'b0);
   assign  _add_map_x_175_up = ((_net_7327)?data_in405:10'b0)|
    ((_net_3335)?data_in406:10'b0);
   assign  _add_map_x_175_right = ((_net_7326)?data_in407:10'b0)|
    ((_net_3334)?data_in404:10'b0);
   assign  _add_map_x_175_down = ((_net_7325)?data_in374:10'b0)|
    ((_net_3333)?data_in373:10'b0);
   assign  _add_map_x_175_left = ((_net_7324)?data_in438:10'b0)|
    ((_net_3332)?data_in437:10'b0);
   assign  _add_map_x_175_start = start;
   assign  _add_map_x_175_goal = goal;
   assign  _add_map_x_175_now = ((_net_7321)?10'b0110010110:10'b0)|
    ((_net_3329)?10'b0110010101:10'b0);
   assign  _add_map_x_175_add_exe = (_net_7320|_net_3328);
   assign  _add_map_x_175_p_reset = p_reset;
   assign  _add_map_x_175_m_clock = m_clock;
   assign  _add_map_x_174_moto_org_near = ((_net_7319)?data_in_org403:10'b0)|
    ((_net_3327)?data_in_org404:10'b0);
   assign  _add_map_x_174_moto_org_near1 = ((_net_7318)?data_in_org405:10'b0)|
    ((_net_3326)?data_in_org402:10'b0);
   assign  _add_map_x_174_moto_org_near2 = ((_net_7317)?data_in_org372:10'b0)|
    ((_net_3325)?data_in_org371:10'b0);
   assign  _add_map_x_174_moto_org_near3 = ((_net_7316)?data_in_org436:10'b0)|
    ((_net_3324)?data_in_org435:10'b0);
   assign  _add_map_x_174_moto_org = ((_net_7315)?data_in_org404:10'b0)|
    ((_net_3323)?data_in_org403:10'b0);
   assign  _add_map_x_174_sg_up = ((_net_7314)?sg_in403:2'b0)|
    ((_net_3322)?sg_in404:2'b0);
   assign  _add_map_x_174_sg_down = ((_net_7313)?sg_in405:2'b0)|
    ((_net_3321)?sg_in402:2'b0);
   assign  _add_map_x_174_sg_left = ((_net_7311)?sg_in436:2'b0)|
    ((_net_3319)?sg_in435:2'b0);
   assign  _add_map_x_174_sg_right = ((_net_7312)?sg_in372:2'b0)|
    ((_net_3320)?sg_in371:2'b0);
   assign  _add_map_x_174_wall_t_in = dig_w;
   assign  _add_map_x_174_moto = ((_net_7309)?data_in404:10'b0)|
    ((_net_3317)?data_in403:10'b0);
   assign  _add_map_x_174_up = ((_net_7308)?data_in403:10'b0)|
    ((_net_3316)?data_in404:10'b0);
   assign  _add_map_x_174_right = ((_net_7307)?data_in405:10'b0)|
    ((_net_3315)?data_in402:10'b0);
   assign  _add_map_x_174_down = ((_net_7306)?data_in372:10'b0)|
    ((_net_3314)?data_in371:10'b0);
   assign  _add_map_x_174_left = ((_net_7305)?data_in436:10'b0)|
    ((_net_3313)?data_in435:10'b0);
   assign  _add_map_x_174_start = start;
   assign  _add_map_x_174_goal = goal;
   assign  _add_map_x_174_now = ((_net_7302)?10'b0110010100:10'b0)|
    ((_net_3310)?10'b0110010011:10'b0);
   assign  _add_map_x_174_add_exe = (_net_7301|_net_3309);
   assign  _add_map_x_174_p_reset = p_reset;
   assign  _add_map_x_174_m_clock = m_clock;
   assign  _add_map_x_173_moto_org_near = ((_net_7300)?data_in_org401:10'b0)|
    ((_net_3308)?data_in_org402:10'b0);
   assign  _add_map_x_173_moto_org_near1 = ((_net_7299)?data_in_org403:10'b0)|
    ((_net_3307)?data_in_org400:10'b0);
   assign  _add_map_x_173_moto_org_near2 = ((_net_7298)?data_in_org370:10'b0)|
    ((_net_3306)?data_in_org369:10'b0);
   assign  _add_map_x_173_moto_org_near3 = ((_net_7297)?data_in_org434:10'b0)|
    ((_net_3305)?data_in_org433:10'b0);
   assign  _add_map_x_173_moto_org = ((_net_7296)?data_in_org402:10'b0)|
    ((_net_3304)?data_in_org401:10'b0);
   assign  _add_map_x_173_sg_up = ((_net_7295)?sg_in401:2'b0)|
    ((_net_3303)?sg_in402:2'b0);
   assign  _add_map_x_173_sg_down = ((_net_7294)?sg_in403:2'b0)|
    ((_net_3302)?sg_in400:2'b0);
   assign  _add_map_x_173_sg_left = ((_net_7292)?sg_in434:2'b0)|
    ((_net_3300)?sg_in433:2'b0);
   assign  _add_map_x_173_sg_right = ((_net_7293)?sg_in370:2'b0)|
    ((_net_3301)?sg_in369:2'b0);
   assign  _add_map_x_173_wall_t_in = dig_w;
   assign  _add_map_x_173_moto = ((_net_7290)?data_in402:10'b0)|
    ((_net_3298)?data_in401:10'b0);
   assign  _add_map_x_173_up = ((_net_7289)?data_in401:10'b0)|
    ((_net_3297)?data_in402:10'b0);
   assign  _add_map_x_173_right = ((_net_7288)?data_in403:10'b0)|
    ((_net_3296)?data_in400:10'b0);
   assign  _add_map_x_173_down = ((_net_7287)?data_in370:10'b0)|
    ((_net_3295)?data_in369:10'b0);
   assign  _add_map_x_173_left = ((_net_7286)?data_in434:10'b0)|
    ((_net_3294)?data_in433:10'b0);
   assign  _add_map_x_173_start = start;
   assign  _add_map_x_173_goal = goal;
   assign  _add_map_x_173_now = ((_net_7283)?10'b0110010010:10'b0)|
    ((_net_3291)?10'b0110010001:10'b0);
   assign  _add_map_x_173_add_exe = (_net_7282|_net_3290);
   assign  _add_map_x_173_p_reset = p_reset;
   assign  _add_map_x_173_m_clock = m_clock;
   assign  _add_map_x_172_moto_org_near = ((_net_7281)?data_in_org399:10'b0)|
    ((_net_3289)?data_in_org400:10'b0);
   assign  _add_map_x_172_moto_org_near1 = ((_net_7280)?data_in_org401:10'b0)|
    ((_net_3288)?data_in_org398:10'b0);
   assign  _add_map_x_172_moto_org_near2 = ((_net_7279)?data_in_org368:10'b0)|
    ((_net_3287)?data_in_org367:10'b0);
   assign  _add_map_x_172_moto_org_near3 = ((_net_7278)?data_in_org432:10'b0)|
    ((_net_3286)?data_in_org431:10'b0);
   assign  _add_map_x_172_moto_org = ((_net_7277)?data_in_org400:10'b0)|
    ((_net_3285)?data_in_org399:10'b0);
   assign  _add_map_x_172_sg_up = ((_net_7276)?sg_in399:2'b0)|
    ((_net_3284)?sg_in400:2'b0);
   assign  _add_map_x_172_sg_down = ((_net_7275)?sg_in401:2'b0)|
    ((_net_3283)?sg_in398:2'b0);
   assign  _add_map_x_172_sg_left = ((_net_7273)?sg_in432:2'b0)|
    ((_net_3281)?sg_in431:2'b0);
   assign  _add_map_x_172_sg_right = ((_net_7274)?sg_in368:2'b0)|
    ((_net_3282)?sg_in367:2'b0);
   assign  _add_map_x_172_wall_t_in = dig_w;
   assign  _add_map_x_172_moto = ((_net_7271)?data_in400:10'b0)|
    ((_net_3279)?data_in399:10'b0);
   assign  _add_map_x_172_up = ((_net_7270)?data_in399:10'b0)|
    ((_net_3278)?data_in400:10'b0);
   assign  _add_map_x_172_right = ((_net_7269)?data_in401:10'b0)|
    ((_net_3277)?data_in398:10'b0);
   assign  _add_map_x_172_down = ((_net_7268)?data_in368:10'b0)|
    ((_net_3276)?data_in367:10'b0);
   assign  _add_map_x_172_left = ((_net_7267)?data_in432:10'b0)|
    ((_net_3275)?data_in431:10'b0);
   assign  _add_map_x_172_start = start;
   assign  _add_map_x_172_goal = goal;
   assign  _add_map_x_172_now = ((_net_7264)?10'b0110010000:10'b0)|
    ((_net_3272)?10'b0110001111:10'b0);
   assign  _add_map_x_172_add_exe = (_net_7263|_net_3271);
   assign  _add_map_x_172_p_reset = p_reset;
   assign  _add_map_x_172_m_clock = m_clock;
   assign  _add_map_x_171_moto_org_near = ((_net_7262)?data_in_org397:10'b0)|
    ((_net_3270)?data_in_org398:10'b0);
   assign  _add_map_x_171_moto_org_near1 = ((_net_7261)?data_in_org399:10'b0)|
    ((_net_3269)?data_in_org396:10'b0);
   assign  _add_map_x_171_moto_org_near2 = ((_net_7260)?data_in_org366:10'b0)|
    ((_net_3268)?data_in_org365:10'b0);
   assign  _add_map_x_171_moto_org_near3 = ((_net_7259)?data_in_org430:10'b0)|
    ((_net_3267)?data_in_org429:10'b0);
   assign  _add_map_x_171_moto_org = ((_net_7258)?data_in_org398:10'b0)|
    ((_net_3266)?data_in_org397:10'b0);
   assign  _add_map_x_171_sg_up = ((_net_7257)?sg_in397:2'b0)|
    ((_net_3265)?sg_in398:2'b0);
   assign  _add_map_x_171_sg_down = ((_net_7256)?sg_in399:2'b0)|
    ((_net_3264)?sg_in396:2'b0);
   assign  _add_map_x_171_sg_left = ((_net_7254)?sg_in430:2'b0)|
    ((_net_3262)?sg_in429:2'b0);
   assign  _add_map_x_171_sg_right = ((_net_7255)?sg_in366:2'b0)|
    ((_net_3263)?sg_in365:2'b0);
   assign  _add_map_x_171_wall_t_in = dig_w;
   assign  _add_map_x_171_moto = ((_net_7252)?data_in398:10'b0)|
    ((_net_3260)?data_in397:10'b0);
   assign  _add_map_x_171_up = ((_net_7251)?data_in397:10'b0)|
    ((_net_3259)?data_in398:10'b0);
   assign  _add_map_x_171_right = ((_net_7250)?data_in399:10'b0)|
    ((_net_3258)?data_in396:10'b0);
   assign  _add_map_x_171_down = ((_net_7249)?data_in366:10'b0)|
    ((_net_3257)?data_in365:10'b0);
   assign  _add_map_x_171_left = ((_net_7248)?data_in430:10'b0)|
    ((_net_3256)?data_in429:10'b0);
   assign  _add_map_x_171_start = start;
   assign  _add_map_x_171_goal = goal;
   assign  _add_map_x_171_now = ((_net_7245)?10'b0110001110:10'b0)|
    ((_net_3253)?10'b0110001101:10'b0);
   assign  _add_map_x_171_add_exe = (_net_7244|_net_3252);
   assign  _add_map_x_171_p_reset = p_reset;
   assign  _add_map_x_171_m_clock = m_clock;
   assign  _add_map_x_170_moto_org_near = ((_net_7243)?data_in_org395:10'b0)|
    ((_net_3251)?data_in_org396:10'b0);
   assign  _add_map_x_170_moto_org_near1 = ((_net_7242)?data_in_org397:10'b0)|
    ((_net_3250)?data_in_org394:10'b0);
   assign  _add_map_x_170_moto_org_near2 = ((_net_7241)?data_in_org364:10'b0)|
    ((_net_3249)?data_in_org363:10'b0);
   assign  _add_map_x_170_moto_org_near3 = ((_net_7240)?data_in_org428:10'b0)|
    ((_net_3248)?data_in_org427:10'b0);
   assign  _add_map_x_170_moto_org = ((_net_7239)?data_in_org396:10'b0)|
    ((_net_3247)?data_in_org395:10'b0);
   assign  _add_map_x_170_sg_up = ((_net_7238)?sg_in395:2'b0)|
    ((_net_3246)?sg_in396:2'b0);
   assign  _add_map_x_170_sg_down = ((_net_7237)?sg_in397:2'b0)|
    ((_net_3245)?sg_in394:2'b0);
   assign  _add_map_x_170_sg_left = ((_net_7235)?sg_in428:2'b0)|
    ((_net_3243)?sg_in427:2'b0);
   assign  _add_map_x_170_sg_right = ((_net_7236)?sg_in364:2'b0)|
    ((_net_3244)?sg_in363:2'b0);
   assign  _add_map_x_170_wall_t_in = dig_w;
   assign  _add_map_x_170_moto = ((_net_7233)?data_in396:10'b0)|
    ((_net_3241)?data_in395:10'b0);
   assign  _add_map_x_170_up = ((_net_7232)?data_in395:10'b0)|
    ((_net_3240)?data_in396:10'b0);
   assign  _add_map_x_170_right = ((_net_7231)?data_in397:10'b0)|
    ((_net_3239)?data_in394:10'b0);
   assign  _add_map_x_170_down = ((_net_7230)?data_in364:10'b0)|
    ((_net_3238)?data_in363:10'b0);
   assign  _add_map_x_170_left = ((_net_7229)?data_in428:10'b0)|
    ((_net_3237)?data_in427:10'b0);
   assign  _add_map_x_170_start = start;
   assign  _add_map_x_170_goal = goal;
   assign  _add_map_x_170_now = ((_net_7226)?10'b0110001100:10'b0)|
    ((_net_3234)?10'b0110001011:10'b0);
   assign  _add_map_x_170_add_exe = (_net_7225|_net_3233);
   assign  _add_map_x_170_p_reset = p_reset;
   assign  _add_map_x_170_m_clock = m_clock;
   assign  _add_map_x_169_moto_org_near = ((_net_7224)?data_in_org393:10'b0)|
    ((_net_3232)?data_in_org394:10'b0);
   assign  _add_map_x_169_moto_org_near1 = ((_net_7223)?data_in_org395:10'b0)|
    ((_net_3231)?data_in_org392:10'b0);
   assign  _add_map_x_169_moto_org_near2 = ((_net_7222)?data_in_org362:10'b0)|
    ((_net_3230)?data_in_org361:10'b0);
   assign  _add_map_x_169_moto_org_near3 = ((_net_7221)?data_in_org426:10'b0)|
    ((_net_3229)?data_in_org425:10'b0);
   assign  _add_map_x_169_moto_org = ((_net_7220)?data_in_org394:10'b0)|
    ((_net_3228)?data_in_org393:10'b0);
   assign  _add_map_x_169_sg_up = ((_net_7219)?sg_in393:2'b0)|
    ((_net_3227)?sg_in394:2'b0);
   assign  _add_map_x_169_sg_down = ((_net_7218)?sg_in395:2'b0)|
    ((_net_3226)?sg_in392:2'b0);
   assign  _add_map_x_169_sg_left = ((_net_7216)?sg_in426:2'b0)|
    ((_net_3224)?sg_in425:2'b0);
   assign  _add_map_x_169_sg_right = ((_net_7217)?sg_in362:2'b0)|
    ((_net_3225)?sg_in361:2'b0);
   assign  _add_map_x_169_wall_t_in = dig_w;
   assign  _add_map_x_169_moto = ((_net_7214)?data_in394:10'b0)|
    ((_net_3222)?data_in393:10'b0);
   assign  _add_map_x_169_up = ((_net_7213)?data_in393:10'b0)|
    ((_net_3221)?data_in394:10'b0);
   assign  _add_map_x_169_right = ((_net_7212)?data_in395:10'b0)|
    ((_net_3220)?data_in392:10'b0);
   assign  _add_map_x_169_down = ((_net_7211)?data_in362:10'b0)|
    ((_net_3219)?data_in361:10'b0);
   assign  _add_map_x_169_left = ((_net_7210)?data_in426:10'b0)|
    ((_net_3218)?data_in425:10'b0);
   assign  _add_map_x_169_start = start;
   assign  _add_map_x_169_goal = goal;
   assign  _add_map_x_169_now = ((_net_7207)?10'b0110001010:10'b0)|
    ((_net_3215)?10'b0110001001:10'b0);
   assign  _add_map_x_169_add_exe = (_net_7206|_net_3214);
   assign  _add_map_x_169_p_reset = p_reset;
   assign  _add_map_x_169_m_clock = m_clock;
   assign  _add_map_x_168_moto_org_near = ((_net_7205)?data_in_org391:10'b0)|
    ((_net_3213)?data_in_org392:10'b0);
   assign  _add_map_x_168_moto_org_near1 = ((_net_7204)?data_in_org393:10'b0)|
    ((_net_3212)?data_in_org390:10'b0);
   assign  _add_map_x_168_moto_org_near2 = ((_net_7203)?data_in_org360:10'b0)|
    ((_net_3211)?data_in_org359:10'b0);
   assign  _add_map_x_168_moto_org_near3 = ((_net_7202)?data_in_org424:10'b0)|
    ((_net_3210)?data_in_org423:10'b0);
   assign  _add_map_x_168_moto_org = ((_net_7201)?data_in_org392:10'b0)|
    ((_net_3209)?data_in_org391:10'b0);
   assign  _add_map_x_168_sg_up = ((_net_7200)?sg_in391:2'b0)|
    ((_net_3208)?sg_in392:2'b0);
   assign  _add_map_x_168_sg_down = ((_net_7199)?sg_in393:2'b0)|
    ((_net_3207)?sg_in390:2'b0);
   assign  _add_map_x_168_sg_left = ((_net_7197)?sg_in424:2'b0)|
    ((_net_3205)?sg_in423:2'b0);
   assign  _add_map_x_168_sg_right = ((_net_7198)?sg_in360:2'b0)|
    ((_net_3206)?sg_in359:2'b0);
   assign  _add_map_x_168_wall_t_in = dig_w;
   assign  _add_map_x_168_moto = ((_net_7195)?data_in392:10'b0)|
    ((_net_3203)?data_in391:10'b0);
   assign  _add_map_x_168_up = ((_net_7194)?data_in391:10'b0)|
    ((_net_3202)?data_in392:10'b0);
   assign  _add_map_x_168_right = ((_net_7193)?data_in393:10'b0)|
    ((_net_3201)?data_in390:10'b0);
   assign  _add_map_x_168_down = ((_net_7192)?data_in360:10'b0)|
    ((_net_3200)?data_in359:10'b0);
   assign  _add_map_x_168_left = ((_net_7191)?data_in424:10'b0)|
    ((_net_3199)?data_in423:10'b0);
   assign  _add_map_x_168_start = start;
   assign  _add_map_x_168_goal = goal;
   assign  _add_map_x_168_now = ((_net_7188)?10'b0110001000:10'b0)|
    ((_net_3196)?10'b0110000111:10'b0);
   assign  _add_map_x_168_add_exe = (_net_7187|_net_3195);
   assign  _add_map_x_168_p_reset = p_reset;
   assign  _add_map_x_168_m_clock = m_clock;
   assign  _add_map_x_167_moto_org_near = ((_net_7186)?data_in_org389:10'b0)|
    ((_net_3194)?data_in_org390:10'b0);
   assign  _add_map_x_167_moto_org_near1 = ((_net_7185)?data_in_org391:10'b0)|
    ((_net_3193)?data_in_org388:10'b0);
   assign  _add_map_x_167_moto_org_near2 = ((_net_7184)?data_in_org358:10'b0)|
    ((_net_3192)?data_in_org357:10'b0);
   assign  _add_map_x_167_moto_org_near3 = ((_net_7183)?data_in_org422:10'b0)|
    ((_net_3191)?data_in_org421:10'b0);
   assign  _add_map_x_167_moto_org = ((_net_7182)?data_in_org390:10'b0)|
    ((_net_3190)?data_in_org389:10'b0);
   assign  _add_map_x_167_sg_up = ((_net_7181)?sg_in389:2'b0)|
    ((_net_3189)?sg_in390:2'b0);
   assign  _add_map_x_167_sg_down = ((_net_7180)?sg_in391:2'b0)|
    ((_net_3188)?sg_in388:2'b0);
   assign  _add_map_x_167_sg_left = ((_net_7178)?sg_in422:2'b0)|
    ((_net_3186)?sg_in421:2'b0);
   assign  _add_map_x_167_sg_right = ((_net_7179)?sg_in358:2'b0)|
    ((_net_3187)?sg_in357:2'b0);
   assign  _add_map_x_167_wall_t_in = dig_w;
   assign  _add_map_x_167_moto = ((_net_7176)?data_in390:10'b0)|
    ((_net_3184)?data_in389:10'b0);
   assign  _add_map_x_167_up = ((_net_7175)?data_in389:10'b0)|
    ((_net_3183)?data_in390:10'b0);
   assign  _add_map_x_167_right = ((_net_7174)?data_in391:10'b0)|
    ((_net_3182)?data_in388:10'b0);
   assign  _add_map_x_167_down = ((_net_7173)?data_in358:10'b0)|
    ((_net_3181)?data_in357:10'b0);
   assign  _add_map_x_167_left = ((_net_7172)?data_in422:10'b0)|
    ((_net_3180)?data_in421:10'b0);
   assign  _add_map_x_167_start = start;
   assign  _add_map_x_167_goal = goal;
   assign  _add_map_x_167_now = ((_net_7169)?10'b0110000110:10'b0)|
    ((_net_3177)?10'b0110000101:10'b0);
   assign  _add_map_x_167_add_exe = (_net_7168|_net_3176);
   assign  _add_map_x_167_p_reset = p_reset;
   assign  _add_map_x_167_m_clock = m_clock;
   assign  _add_map_x_166_moto_org_near = ((_net_7167)?data_in_org387:10'b0)|
    ((_net_3175)?data_in_org388:10'b0);
   assign  _add_map_x_166_moto_org_near1 = ((_net_7166)?data_in_org389:10'b0)|
    ((_net_3174)?data_in_org386:10'b0);
   assign  _add_map_x_166_moto_org_near2 = ((_net_7165)?data_in_org356:10'b0)|
    ((_net_3173)?data_in_org355:10'b0);
   assign  _add_map_x_166_moto_org_near3 = ((_net_7164)?data_in_org420:10'b0)|
    ((_net_3172)?data_in_org419:10'b0);
   assign  _add_map_x_166_moto_org = ((_net_7163)?data_in_org388:10'b0)|
    ((_net_3171)?data_in_org387:10'b0);
   assign  _add_map_x_166_sg_up = ((_net_7162)?sg_in387:2'b0)|
    ((_net_3170)?sg_in388:2'b0);
   assign  _add_map_x_166_sg_down = ((_net_7161)?sg_in389:2'b0)|
    ((_net_3169)?sg_in386:2'b0);
   assign  _add_map_x_166_sg_left = ((_net_7159)?sg_in420:2'b0)|
    ((_net_3167)?sg_in419:2'b0);
   assign  _add_map_x_166_sg_right = ((_net_7160)?sg_in356:2'b0)|
    ((_net_3168)?sg_in355:2'b0);
   assign  _add_map_x_166_wall_t_in = dig_w;
   assign  _add_map_x_166_moto = ((_net_7157)?data_in388:10'b0)|
    ((_net_3165)?data_in387:10'b0);
   assign  _add_map_x_166_up = ((_net_7156)?data_in387:10'b0)|
    ((_net_3164)?data_in388:10'b0);
   assign  _add_map_x_166_right = ((_net_7155)?data_in389:10'b0)|
    ((_net_3163)?data_in386:10'b0);
   assign  _add_map_x_166_down = ((_net_7154)?data_in356:10'b0)|
    ((_net_3162)?data_in355:10'b0);
   assign  _add_map_x_166_left = ((_net_7153)?data_in420:10'b0)|
    ((_net_3161)?data_in419:10'b0);
   assign  _add_map_x_166_start = start;
   assign  _add_map_x_166_goal = goal;
   assign  _add_map_x_166_now = ((_net_7150)?10'b0110000100:10'b0)|
    ((_net_3158)?10'b0110000011:10'b0);
   assign  _add_map_x_166_add_exe = (_net_7149|_net_3157);
   assign  _add_map_x_166_p_reset = p_reset;
   assign  _add_map_x_166_m_clock = m_clock;
   assign  _add_map_x_165_moto_org_near = ((_net_7148)?data_in_org385:10'b0)|
    ((_net_3156)?data_in_org386:10'b0);
   assign  _add_map_x_165_moto_org_near1 = ((_net_7147)?data_in_org387:10'b0)|
    ((_net_3155)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_165_moto_org_near2 = ((_net_7146)?data_in_org354:10'b0)|
    ((_net_3154)?data_in_org353:10'b0);
   assign  _add_map_x_165_moto_org_near3 = ((_net_7145)?data_in_org418:10'b0)|
    ((_net_3153)?data_in_org417:10'b0);
   assign  _add_map_x_165_moto_org = ((_net_7144)?data_in_org386:10'b0)|
    ((_net_3152)?data_in_org385:10'b0);
   assign  _add_map_x_165_sg_up = ((_net_7143)?sg_in385:2'b0)|
    ((_net_3151)?sg_in386:2'b0);
   assign  _add_map_x_165_sg_down = ((_net_7142)?sg_in387:2'b0)|
    ((_net_3150)?3'b000:2'b0);
   assign  _add_map_x_165_sg_left = ((_net_7140)?sg_in418:2'b0)|
    ((_net_3148)?sg_in417:2'b0);
   assign  _add_map_x_165_sg_right = ((_net_7141)?sg_in354:2'b0)|
    ((_net_3149)?sg_in353:2'b0);
   assign  _add_map_x_165_wall_t_in = dig_w;
   assign  _add_map_x_165_moto = ((_net_7138)?data_in386:10'b0)|
    ((_net_3146)?data_in385:10'b0);
   assign  _add_map_x_165_up = ((_net_7137)?data_in385:10'b0)|
    ((_net_3145)?data_in386:10'b0);
   assign  _add_map_x_165_right = ((_net_7136)?data_in387:10'b0)|
    ((_net_3144)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_165_down = ((_net_7135)?data_in354:10'b0)|
    ((_net_3143)?data_in353:10'b0);
   assign  _add_map_x_165_left = ((_net_7134)?data_in418:10'b0)|
    ((_net_3142)?data_in417:10'b0);
   assign  _add_map_x_165_start = start;
   assign  _add_map_x_165_goal = goal;
   assign  _add_map_x_165_now = ((_net_7131)?10'b0110000010:10'b0)|
    ((_net_3139)?10'b0110000001:10'b0);
   assign  _add_map_x_165_add_exe = (_net_7130|_net_3138);
   assign  _add_map_x_165_p_reset = p_reset;
   assign  _add_map_x_165_m_clock = m_clock;
   assign  _add_map_x_164_moto_org_near = ((_net_7129)?data_in_org382:10'b0)|
    ((_net_3137)?data_in_org381:10'b0);
   assign  _add_map_x_164_moto_org_near1 = ((_net_7128)?data_in_org380:10'b0)|
    ((_net_3136)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_164_moto_org_near2 = ((_net_7127)?data_in_org349:10'b0)|
    ((_net_3135)?data_in_org350:10'b0);
   assign  _add_map_x_164_moto_org_near3 = ((_net_7126)?data_in_org413:10'b0)|
    ((_net_3134)?data_in_org414:10'b0);
   assign  _add_map_x_164_moto_org = ((_net_7125)?data_in_org381:10'b0)|
    ((_net_3133)?data_in_org382:10'b0);
   assign  _add_map_x_164_sg_up = ((_net_7124)?sg_in382:2'b0)|
    ((_net_3132)?sg_in381:2'b0);
   assign  _add_map_x_164_sg_down = ((_net_7123)?sg_in349:2'b0)|
    ((_net_3131)?3'b000:2'b0);
   assign  _add_map_x_164_sg_left = ((_net_7121)?sg_in413:2'b0)|
    ((_net_3129)?sg_in414:2'b0);
   assign  _add_map_x_164_sg_right = ((_net_7122)?sg_in380:2'b0)|
    ((_net_3130)?sg_in350:2'b0);
   assign  _add_map_x_164_wall_t_in = dig_w;
   assign  _add_map_x_164_moto = ((_net_7119)?data_in381:10'b0)|
    ((_net_3127)?data_in382:10'b0);
   assign  _add_map_x_164_up = ((_net_7118)?data_in382:10'b0)|
    ((_net_3126)?data_in381:10'b0);
   assign  _add_map_x_164_right = ((_net_7117)?data_in380:10'b0)|
    ((_net_3125)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_164_down = ((_net_7116)?data_in349:10'b0)|
    ((_net_3124)?data_in350:10'b0);
   assign  _add_map_x_164_left = ((_net_7115)?data_in413:10'b0)|
    ((_net_3123)?data_in414:10'b0);
   assign  _add_map_x_164_start = start;
   assign  _add_map_x_164_goal = goal;
   assign  _add_map_x_164_now = ((_net_7112)?10'b0101111101:10'b0)|
    ((_net_3120)?10'b0101111110:10'b0);
   assign  _add_map_x_164_add_exe = (_net_7111|_net_3119);
   assign  _add_map_x_164_p_reset = p_reset;
   assign  _add_map_x_164_m_clock = m_clock;
   assign  _add_map_x_163_moto_org_near = ((_net_7110)?data_in_org380:10'b0)|
    ((_net_3118)?data_in_org379:10'b0);
   assign  _add_map_x_163_moto_org_near1 = ((_net_7109)?data_in_org378:10'b0)|
    ((_net_3117)?data_in_org381:10'b0);
   assign  _add_map_x_163_moto_org_near2 = ((_net_7108)?data_in_org347:10'b0)|
    ((_net_3116)?data_in_org348:10'b0);
   assign  _add_map_x_163_moto_org_near3 = ((_net_7107)?data_in_org411:10'b0)|
    ((_net_3115)?data_in_org412:10'b0);
   assign  _add_map_x_163_moto_org = ((_net_7106)?data_in_org379:10'b0)|
    ((_net_3114)?data_in_org380:10'b0);
   assign  _add_map_x_163_sg_up = ((_net_7105)?sg_in380:2'b0)|
    ((_net_3113)?sg_in379:2'b0);
   assign  _add_map_x_163_sg_down = ((_net_7104)?sg_in347:2'b0)|
    ((_net_3112)?sg_in381:2'b0);
   assign  _add_map_x_163_sg_left = ((_net_7102)?sg_in411:2'b0)|
    ((_net_3110)?sg_in412:2'b0);
   assign  _add_map_x_163_sg_right = ((_net_7103)?sg_in378:2'b0)|
    ((_net_3111)?sg_in348:2'b0);
   assign  _add_map_x_163_wall_t_in = dig_w;
   assign  _add_map_x_163_moto = ((_net_7100)?data_in379:10'b0)|
    ((_net_3108)?data_in380:10'b0);
   assign  _add_map_x_163_up = ((_net_7099)?data_in380:10'b0)|
    ((_net_3107)?data_in379:10'b0);
   assign  _add_map_x_163_right = ((_net_7098)?data_in378:10'b0)|
    ((_net_3106)?data_in381:10'b0);
   assign  _add_map_x_163_down = ((_net_7097)?data_in347:10'b0)|
    ((_net_3105)?data_in348:10'b0);
   assign  _add_map_x_163_left = ((_net_7096)?data_in411:10'b0)|
    ((_net_3104)?data_in412:10'b0);
   assign  _add_map_x_163_start = start;
   assign  _add_map_x_163_goal = goal;
   assign  _add_map_x_163_now = ((_net_7093)?10'b0101111011:10'b0)|
    ((_net_3101)?10'b0101111100:10'b0);
   assign  _add_map_x_163_add_exe = (_net_7092|_net_3100);
   assign  _add_map_x_163_p_reset = p_reset;
   assign  _add_map_x_163_m_clock = m_clock;
   assign  _add_map_x_162_moto_org_near = ((_net_7091)?data_in_org378:10'b0)|
    ((_net_3099)?data_in_org377:10'b0);
   assign  _add_map_x_162_moto_org_near1 = ((_net_7090)?data_in_org376:10'b0)|
    ((_net_3098)?data_in_org379:10'b0);
   assign  _add_map_x_162_moto_org_near2 = ((_net_7089)?data_in_org345:10'b0)|
    ((_net_3097)?data_in_org346:10'b0);
   assign  _add_map_x_162_moto_org_near3 = ((_net_7088)?data_in_org409:10'b0)|
    ((_net_3096)?data_in_org410:10'b0);
   assign  _add_map_x_162_moto_org = ((_net_7087)?data_in_org377:10'b0)|
    ((_net_3095)?data_in_org378:10'b0);
   assign  _add_map_x_162_sg_up = ((_net_7086)?sg_in378:2'b0)|
    ((_net_3094)?sg_in377:2'b0);
   assign  _add_map_x_162_sg_down = ((_net_7085)?sg_in345:2'b0)|
    ((_net_3093)?sg_in379:2'b0);
   assign  _add_map_x_162_sg_left = ((_net_7083)?sg_in409:2'b0)|
    ((_net_3091)?sg_in410:2'b0);
   assign  _add_map_x_162_sg_right = ((_net_7084)?sg_in376:2'b0)|
    ((_net_3092)?sg_in346:2'b0);
   assign  _add_map_x_162_wall_t_in = dig_w;
   assign  _add_map_x_162_moto = ((_net_7081)?data_in377:10'b0)|
    ((_net_3089)?data_in378:10'b0);
   assign  _add_map_x_162_up = ((_net_7080)?data_in378:10'b0)|
    ((_net_3088)?data_in377:10'b0);
   assign  _add_map_x_162_right = ((_net_7079)?data_in376:10'b0)|
    ((_net_3087)?data_in379:10'b0);
   assign  _add_map_x_162_down = ((_net_7078)?data_in345:10'b0)|
    ((_net_3086)?data_in346:10'b0);
   assign  _add_map_x_162_left = ((_net_7077)?data_in409:10'b0)|
    ((_net_3085)?data_in410:10'b0);
   assign  _add_map_x_162_start = start;
   assign  _add_map_x_162_goal = goal;
   assign  _add_map_x_162_now = ((_net_7074)?10'b0101111001:10'b0)|
    ((_net_3082)?10'b0101111010:10'b0);
   assign  _add_map_x_162_add_exe = (_net_7073|_net_3081);
   assign  _add_map_x_162_p_reset = p_reset;
   assign  _add_map_x_162_m_clock = m_clock;
   assign  _add_map_x_161_moto_org_near = ((_net_7072)?data_in_org376:10'b0)|
    ((_net_3080)?data_in_org375:10'b0);
   assign  _add_map_x_161_moto_org_near1 = ((_net_7071)?data_in_org374:10'b0)|
    ((_net_3079)?data_in_org377:10'b0);
   assign  _add_map_x_161_moto_org_near2 = ((_net_7070)?data_in_org343:10'b0)|
    ((_net_3078)?data_in_org344:10'b0);
   assign  _add_map_x_161_moto_org_near3 = ((_net_7069)?data_in_org407:10'b0)|
    ((_net_3077)?data_in_org408:10'b0);
   assign  _add_map_x_161_moto_org = ((_net_7068)?data_in_org375:10'b0)|
    ((_net_3076)?data_in_org376:10'b0);
   assign  _add_map_x_161_sg_up = ((_net_7067)?sg_in376:2'b0)|
    ((_net_3075)?sg_in375:2'b0);
   assign  _add_map_x_161_sg_down = ((_net_7066)?sg_in343:2'b0)|
    ((_net_3074)?sg_in377:2'b0);
   assign  _add_map_x_161_sg_left = ((_net_7064)?sg_in407:2'b0)|
    ((_net_3072)?sg_in408:2'b0);
   assign  _add_map_x_161_sg_right = ((_net_7065)?sg_in374:2'b0)|
    ((_net_3073)?sg_in344:2'b0);
   assign  _add_map_x_161_wall_t_in = dig_w;
   assign  _add_map_x_161_moto = ((_net_7062)?data_in375:10'b0)|
    ((_net_3070)?data_in376:10'b0);
   assign  _add_map_x_161_up = ((_net_7061)?data_in376:10'b0)|
    ((_net_3069)?data_in375:10'b0);
   assign  _add_map_x_161_right = ((_net_7060)?data_in374:10'b0)|
    ((_net_3068)?data_in377:10'b0);
   assign  _add_map_x_161_down = ((_net_7059)?data_in343:10'b0)|
    ((_net_3067)?data_in344:10'b0);
   assign  _add_map_x_161_left = ((_net_7058)?data_in407:10'b0)|
    ((_net_3066)?data_in408:10'b0);
   assign  _add_map_x_161_start = start;
   assign  _add_map_x_161_goal = goal;
   assign  _add_map_x_161_now = ((_net_7055)?10'b0101110111:10'b0)|
    ((_net_3063)?10'b0101111000:10'b0);
   assign  _add_map_x_161_add_exe = (_net_7054|_net_3062);
   assign  _add_map_x_161_p_reset = p_reset;
   assign  _add_map_x_161_m_clock = m_clock;
   assign  _add_map_x_160_moto_org_near = ((_net_7053)?data_in_org374:10'b0)|
    ((_net_3061)?data_in_org373:10'b0);
   assign  _add_map_x_160_moto_org_near1 = ((_net_7052)?data_in_org372:10'b0)|
    ((_net_3060)?data_in_org375:10'b0);
   assign  _add_map_x_160_moto_org_near2 = ((_net_7051)?data_in_org341:10'b0)|
    ((_net_3059)?data_in_org342:10'b0);
   assign  _add_map_x_160_moto_org_near3 = ((_net_7050)?data_in_org405:10'b0)|
    ((_net_3058)?data_in_org406:10'b0);
   assign  _add_map_x_160_moto_org = ((_net_7049)?data_in_org373:10'b0)|
    ((_net_3057)?data_in_org374:10'b0);
   assign  _add_map_x_160_sg_up = ((_net_7048)?sg_in374:2'b0)|
    ((_net_3056)?sg_in373:2'b0);
   assign  _add_map_x_160_sg_down = ((_net_7047)?sg_in341:2'b0)|
    ((_net_3055)?sg_in375:2'b0);
   assign  _add_map_x_160_sg_left = ((_net_7045)?sg_in405:2'b0)|
    ((_net_3053)?sg_in406:2'b0);
   assign  _add_map_x_160_sg_right = ((_net_7046)?sg_in372:2'b0)|
    ((_net_3054)?sg_in342:2'b0);
   assign  _add_map_x_160_wall_t_in = dig_w;
   assign  _add_map_x_160_moto = ((_net_7043)?data_in373:10'b0)|
    ((_net_3051)?data_in374:10'b0);
   assign  _add_map_x_160_up = ((_net_7042)?data_in374:10'b0)|
    ((_net_3050)?data_in373:10'b0);
   assign  _add_map_x_160_right = ((_net_7041)?data_in372:10'b0)|
    ((_net_3049)?data_in375:10'b0);
   assign  _add_map_x_160_down = ((_net_7040)?data_in341:10'b0)|
    ((_net_3048)?data_in342:10'b0);
   assign  _add_map_x_160_left = ((_net_7039)?data_in405:10'b0)|
    ((_net_3047)?data_in406:10'b0);
   assign  _add_map_x_160_start = start;
   assign  _add_map_x_160_goal = goal;
   assign  _add_map_x_160_now = ((_net_7036)?10'b0101110101:10'b0)|
    ((_net_3044)?10'b0101110110:10'b0);
   assign  _add_map_x_160_add_exe = (_net_7035|_net_3043);
   assign  _add_map_x_160_p_reset = p_reset;
   assign  _add_map_x_160_m_clock = m_clock;
   assign  _add_map_x_159_moto_org_near = ((_net_7034)?data_in_org372:10'b0)|
    ((_net_3042)?data_in_org371:10'b0);
   assign  _add_map_x_159_moto_org_near1 = ((_net_7033)?data_in_org370:10'b0)|
    ((_net_3041)?data_in_org373:10'b0);
   assign  _add_map_x_159_moto_org_near2 = ((_net_7032)?data_in_org339:10'b0)|
    ((_net_3040)?data_in_org340:10'b0);
   assign  _add_map_x_159_moto_org_near3 = ((_net_7031)?data_in_org403:10'b0)|
    ((_net_3039)?data_in_org404:10'b0);
   assign  _add_map_x_159_moto_org = ((_net_7030)?data_in_org371:10'b0)|
    ((_net_3038)?data_in_org372:10'b0);
   assign  _add_map_x_159_sg_up = ((_net_7029)?sg_in372:2'b0)|
    ((_net_3037)?sg_in371:2'b0);
   assign  _add_map_x_159_sg_down = ((_net_7028)?sg_in339:2'b0)|
    ((_net_3036)?sg_in373:2'b0);
   assign  _add_map_x_159_sg_left = ((_net_7026)?sg_in403:2'b0)|
    ((_net_3034)?sg_in404:2'b0);
   assign  _add_map_x_159_sg_right = ((_net_7027)?sg_in370:2'b0)|
    ((_net_3035)?sg_in340:2'b0);
   assign  _add_map_x_159_wall_t_in = dig_w;
   assign  _add_map_x_159_moto = ((_net_7024)?data_in371:10'b0)|
    ((_net_3032)?data_in372:10'b0);
   assign  _add_map_x_159_up = ((_net_7023)?data_in372:10'b0)|
    ((_net_3031)?data_in371:10'b0);
   assign  _add_map_x_159_right = ((_net_7022)?data_in370:10'b0)|
    ((_net_3030)?data_in373:10'b0);
   assign  _add_map_x_159_down = ((_net_7021)?data_in339:10'b0)|
    ((_net_3029)?data_in340:10'b0);
   assign  _add_map_x_159_left = ((_net_7020)?data_in403:10'b0)|
    ((_net_3028)?data_in404:10'b0);
   assign  _add_map_x_159_start = start;
   assign  _add_map_x_159_goal = goal;
   assign  _add_map_x_159_now = ((_net_7017)?10'b0101110011:10'b0)|
    ((_net_3025)?10'b0101110100:10'b0);
   assign  _add_map_x_159_add_exe = (_net_7016|_net_3024);
   assign  _add_map_x_159_p_reset = p_reset;
   assign  _add_map_x_159_m_clock = m_clock;
   assign  _add_map_x_158_moto_org_near = ((_net_7015)?data_in_org370:10'b0)|
    ((_net_3023)?data_in_org369:10'b0);
   assign  _add_map_x_158_moto_org_near1 = ((_net_7014)?data_in_org368:10'b0)|
    ((_net_3022)?data_in_org371:10'b0);
   assign  _add_map_x_158_moto_org_near2 = ((_net_7013)?data_in_org337:10'b0)|
    ((_net_3021)?data_in_org338:10'b0);
   assign  _add_map_x_158_moto_org_near3 = ((_net_7012)?data_in_org401:10'b0)|
    ((_net_3020)?data_in_org402:10'b0);
   assign  _add_map_x_158_moto_org = ((_net_7011)?data_in_org369:10'b0)|
    ((_net_3019)?data_in_org370:10'b0);
   assign  _add_map_x_158_sg_up = ((_net_7010)?sg_in370:2'b0)|
    ((_net_3018)?sg_in369:2'b0);
   assign  _add_map_x_158_sg_down = ((_net_7009)?sg_in337:2'b0)|
    ((_net_3017)?sg_in371:2'b0);
   assign  _add_map_x_158_sg_left = ((_net_7007)?sg_in401:2'b0)|
    ((_net_3015)?sg_in402:2'b0);
   assign  _add_map_x_158_sg_right = ((_net_7008)?sg_in368:2'b0)|
    ((_net_3016)?sg_in338:2'b0);
   assign  _add_map_x_158_wall_t_in = dig_w;
   assign  _add_map_x_158_moto = ((_net_7005)?data_in369:10'b0)|
    ((_net_3013)?data_in370:10'b0);
   assign  _add_map_x_158_up = ((_net_7004)?data_in370:10'b0)|
    ((_net_3012)?data_in369:10'b0);
   assign  _add_map_x_158_right = ((_net_7003)?data_in368:10'b0)|
    ((_net_3011)?data_in371:10'b0);
   assign  _add_map_x_158_down = ((_net_7002)?data_in337:10'b0)|
    ((_net_3010)?data_in338:10'b0);
   assign  _add_map_x_158_left = ((_net_7001)?data_in401:10'b0)|
    ((_net_3009)?data_in402:10'b0);
   assign  _add_map_x_158_start = start;
   assign  _add_map_x_158_goal = goal;
   assign  _add_map_x_158_now = ((_net_6998)?10'b0101110001:10'b0)|
    ((_net_3006)?10'b0101110010:10'b0);
   assign  _add_map_x_158_add_exe = (_net_6997|_net_3005);
   assign  _add_map_x_158_p_reset = p_reset;
   assign  _add_map_x_158_m_clock = m_clock;
   assign  _add_map_x_157_moto_org_near = ((_net_6996)?data_in_org368:10'b0)|
    ((_net_3004)?data_in_org367:10'b0);
   assign  _add_map_x_157_moto_org_near1 = ((_net_6995)?data_in_org366:10'b0)|
    ((_net_3003)?data_in_org369:10'b0);
   assign  _add_map_x_157_moto_org_near2 = ((_net_6994)?data_in_org335:10'b0)|
    ((_net_3002)?data_in_org336:10'b0);
   assign  _add_map_x_157_moto_org_near3 = ((_net_6993)?data_in_org399:10'b0)|
    ((_net_3001)?data_in_org400:10'b0);
   assign  _add_map_x_157_moto_org = ((_net_6992)?data_in_org367:10'b0)|
    ((_net_3000)?data_in_org368:10'b0);
   assign  _add_map_x_157_sg_up = ((_net_6991)?sg_in368:2'b0)|
    ((_net_2999)?sg_in367:2'b0);
   assign  _add_map_x_157_sg_down = ((_net_6990)?sg_in335:2'b0)|
    ((_net_2998)?sg_in369:2'b0);
   assign  _add_map_x_157_sg_left = ((_net_6988)?sg_in399:2'b0)|
    ((_net_2996)?sg_in400:2'b0);
   assign  _add_map_x_157_sg_right = ((_net_6989)?sg_in366:2'b0)|
    ((_net_2997)?sg_in336:2'b0);
   assign  _add_map_x_157_wall_t_in = dig_w;
   assign  _add_map_x_157_moto = ((_net_6986)?data_in367:10'b0)|
    ((_net_2994)?data_in368:10'b0);
   assign  _add_map_x_157_up = ((_net_6985)?data_in368:10'b0)|
    ((_net_2993)?data_in367:10'b0);
   assign  _add_map_x_157_right = ((_net_6984)?data_in366:10'b0)|
    ((_net_2992)?data_in369:10'b0);
   assign  _add_map_x_157_down = ((_net_6983)?data_in335:10'b0)|
    ((_net_2991)?data_in336:10'b0);
   assign  _add_map_x_157_left = ((_net_6982)?data_in399:10'b0)|
    ((_net_2990)?data_in400:10'b0);
   assign  _add_map_x_157_start = start;
   assign  _add_map_x_157_goal = goal;
   assign  _add_map_x_157_now = ((_net_6979)?10'b0101101111:10'b0)|
    ((_net_2987)?10'b0101110000:10'b0);
   assign  _add_map_x_157_add_exe = (_net_6978|_net_2986);
   assign  _add_map_x_157_p_reset = p_reset;
   assign  _add_map_x_157_m_clock = m_clock;
   assign  _add_map_x_156_moto_org_near = ((_net_6977)?data_in_org366:10'b0)|
    ((_net_2985)?data_in_org365:10'b0);
   assign  _add_map_x_156_moto_org_near1 = ((_net_6976)?data_in_org364:10'b0)|
    ((_net_2984)?data_in_org367:10'b0);
   assign  _add_map_x_156_moto_org_near2 = ((_net_6975)?data_in_org333:10'b0)|
    ((_net_2983)?data_in_org334:10'b0);
   assign  _add_map_x_156_moto_org_near3 = ((_net_6974)?data_in_org397:10'b0)|
    ((_net_2982)?data_in_org398:10'b0);
   assign  _add_map_x_156_moto_org = ((_net_6973)?data_in_org365:10'b0)|
    ((_net_2981)?data_in_org366:10'b0);
   assign  _add_map_x_156_sg_up = ((_net_6972)?sg_in366:2'b0)|
    ((_net_2980)?sg_in365:2'b0);
   assign  _add_map_x_156_sg_down = ((_net_6971)?sg_in333:2'b0)|
    ((_net_2979)?sg_in367:2'b0);
   assign  _add_map_x_156_sg_left = ((_net_6969)?sg_in397:2'b0)|
    ((_net_2977)?sg_in398:2'b0);
   assign  _add_map_x_156_sg_right = ((_net_6970)?sg_in364:2'b0)|
    ((_net_2978)?sg_in334:2'b0);
   assign  _add_map_x_156_wall_t_in = dig_w;
   assign  _add_map_x_156_moto = ((_net_6967)?data_in365:10'b0)|
    ((_net_2975)?data_in366:10'b0);
   assign  _add_map_x_156_up = ((_net_6966)?data_in366:10'b0)|
    ((_net_2974)?data_in365:10'b0);
   assign  _add_map_x_156_right = ((_net_6965)?data_in364:10'b0)|
    ((_net_2973)?data_in367:10'b0);
   assign  _add_map_x_156_down = ((_net_6964)?data_in333:10'b0)|
    ((_net_2972)?data_in334:10'b0);
   assign  _add_map_x_156_left = ((_net_6963)?data_in397:10'b0)|
    ((_net_2971)?data_in398:10'b0);
   assign  _add_map_x_156_start = start;
   assign  _add_map_x_156_goal = goal;
   assign  _add_map_x_156_now = ((_net_6960)?10'b0101101101:10'b0)|
    ((_net_2968)?10'b0101101110:10'b0);
   assign  _add_map_x_156_add_exe = (_net_6959|_net_2967);
   assign  _add_map_x_156_p_reset = p_reset;
   assign  _add_map_x_156_m_clock = m_clock;
   assign  _add_map_x_155_moto_org_near = ((_net_6958)?data_in_org364:10'b0)|
    ((_net_2966)?data_in_org363:10'b0);
   assign  _add_map_x_155_moto_org_near1 = ((_net_6957)?data_in_org362:10'b0)|
    ((_net_2965)?data_in_org365:10'b0);
   assign  _add_map_x_155_moto_org_near2 = ((_net_6956)?data_in_org331:10'b0)|
    ((_net_2964)?data_in_org332:10'b0);
   assign  _add_map_x_155_moto_org_near3 = ((_net_6955)?data_in_org395:10'b0)|
    ((_net_2963)?data_in_org396:10'b0);
   assign  _add_map_x_155_moto_org = ((_net_6954)?data_in_org363:10'b0)|
    ((_net_2962)?data_in_org364:10'b0);
   assign  _add_map_x_155_sg_up = ((_net_6953)?sg_in364:2'b0)|
    ((_net_2961)?sg_in363:2'b0);
   assign  _add_map_x_155_sg_down = ((_net_6952)?sg_in331:2'b0)|
    ((_net_2960)?sg_in365:2'b0);
   assign  _add_map_x_155_sg_left = ((_net_6950)?sg_in395:2'b0)|
    ((_net_2958)?sg_in396:2'b0);
   assign  _add_map_x_155_sg_right = ((_net_6951)?sg_in362:2'b0)|
    ((_net_2959)?sg_in332:2'b0);
   assign  _add_map_x_155_wall_t_in = dig_w;
   assign  _add_map_x_155_moto = ((_net_6948)?data_in363:10'b0)|
    ((_net_2956)?data_in364:10'b0);
   assign  _add_map_x_155_up = ((_net_6947)?data_in364:10'b0)|
    ((_net_2955)?data_in363:10'b0);
   assign  _add_map_x_155_right = ((_net_6946)?data_in362:10'b0)|
    ((_net_2954)?data_in365:10'b0);
   assign  _add_map_x_155_down = ((_net_6945)?data_in331:10'b0)|
    ((_net_2953)?data_in332:10'b0);
   assign  _add_map_x_155_left = ((_net_6944)?data_in395:10'b0)|
    ((_net_2952)?data_in396:10'b0);
   assign  _add_map_x_155_start = start;
   assign  _add_map_x_155_goal = goal;
   assign  _add_map_x_155_now = ((_net_6941)?10'b0101101011:10'b0)|
    ((_net_2949)?10'b0101101100:10'b0);
   assign  _add_map_x_155_add_exe = (_net_6940|_net_2948);
   assign  _add_map_x_155_p_reset = p_reset;
   assign  _add_map_x_155_m_clock = m_clock;
   assign  _add_map_x_154_moto_org_near = ((_net_6939)?data_in_org362:10'b0)|
    ((_net_2947)?data_in_org361:10'b0);
   assign  _add_map_x_154_moto_org_near1 = ((_net_6938)?data_in_org360:10'b0)|
    ((_net_2946)?data_in_org363:10'b0);
   assign  _add_map_x_154_moto_org_near2 = ((_net_6937)?data_in_org329:10'b0)|
    ((_net_2945)?data_in_org330:10'b0);
   assign  _add_map_x_154_moto_org_near3 = ((_net_6936)?data_in_org393:10'b0)|
    ((_net_2944)?data_in_org394:10'b0);
   assign  _add_map_x_154_moto_org = ((_net_6935)?data_in_org361:10'b0)|
    ((_net_2943)?data_in_org362:10'b0);
   assign  _add_map_x_154_sg_up = ((_net_6934)?sg_in362:2'b0)|
    ((_net_2942)?sg_in361:2'b0);
   assign  _add_map_x_154_sg_down = ((_net_6933)?sg_in329:2'b0)|
    ((_net_2941)?sg_in363:2'b0);
   assign  _add_map_x_154_sg_left = ((_net_6931)?sg_in393:2'b0)|
    ((_net_2939)?sg_in394:2'b0);
   assign  _add_map_x_154_sg_right = ((_net_6932)?sg_in360:2'b0)|
    ((_net_2940)?sg_in330:2'b0);
   assign  _add_map_x_154_wall_t_in = dig_w;
   assign  _add_map_x_154_moto = ((_net_6929)?data_in361:10'b0)|
    ((_net_2937)?data_in362:10'b0);
   assign  _add_map_x_154_up = ((_net_6928)?data_in362:10'b0)|
    ((_net_2936)?data_in361:10'b0);
   assign  _add_map_x_154_right = ((_net_6927)?data_in360:10'b0)|
    ((_net_2935)?data_in363:10'b0);
   assign  _add_map_x_154_down = ((_net_6926)?data_in329:10'b0)|
    ((_net_2934)?data_in330:10'b0);
   assign  _add_map_x_154_left = ((_net_6925)?data_in393:10'b0)|
    ((_net_2933)?data_in394:10'b0);
   assign  _add_map_x_154_start = start;
   assign  _add_map_x_154_goal = goal;
   assign  _add_map_x_154_now = ((_net_6922)?10'b0101101001:10'b0)|
    ((_net_2930)?10'b0101101010:10'b0);
   assign  _add_map_x_154_add_exe = (_net_6921|_net_2929);
   assign  _add_map_x_154_p_reset = p_reset;
   assign  _add_map_x_154_m_clock = m_clock;
   assign  _add_map_x_153_moto_org_near = ((_net_6920)?data_in_org360:10'b0)|
    ((_net_2928)?data_in_org359:10'b0);
   assign  _add_map_x_153_moto_org_near1 = ((_net_6919)?data_in_org358:10'b0)|
    ((_net_2927)?data_in_org361:10'b0);
   assign  _add_map_x_153_moto_org_near2 = ((_net_6918)?data_in_org327:10'b0)|
    ((_net_2926)?data_in_org328:10'b0);
   assign  _add_map_x_153_moto_org_near3 = ((_net_6917)?data_in_org391:10'b0)|
    ((_net_2925)?data_in_org392:10'b0);
   assign  _add_map_x_153_moto_org = ((_net_6916)?data_in_org359:10'b0)|
    ((_net_2924)?data_in_org360:10'b0);
   assign  _add_map_x_153_sg_up = ((_net_6915)?sg_in360:2'b0)|
    ((_net_2923)?sg_in359:2'b0);
   assign  _add_map_x_153_sg_down = ((_net_6914)?sg_in327:2'b0)|
    ((_net_2922)?sg_in361:2'b0);
   assign  _add_map_x_153_sg_left = ((_net_6912)?sg_in391:2'b0)|
    ((_net_2920)?sg_in392:2'b0);
   assign  _add_map_x_153_sg_right = ((_net_6913)?sg_in358:2'b0)|
    ((_net_2921)?sg_in328:2'b0);
   assign  _add_map_x_153_wall_t_in = dig_w;
   assign  _add_map_x_153_moto = ((_net_6910)?data_in359:10'b0)|
    ((_net_2918)?data_in360:10'b0);
   assign  _add_map_x_153_up = ((_net_6909)?data_in360:10'b0)|
    ((_net_2917)?data_in359:10'b0);
   assign  _add_map_x_153_right = ((_net_6908)?data_in358:10'b0)|
    ((_net_2916)?data_in361:10'b0);
   assign  _add_map_x_153_down = ((_net_6907)?data_in327:10'b0)|
    ((_net_2915)?data_in328:10'b0);
   assign  _add_map_x_153_left = ((_net_6906)?data_in391:10'b0)|
    ((_net_2914)?data_in392:10'b0);
   assign  _add_map_x_153_start = start;
   assign  _add_map_x_153_goal = goal;
   assign  _add_map_x_153_now = ((_net_6903)?10'b0101100111:10'b0)|
    ((_net_2911)?10'b0101101000:10'b0);
   assign  _add_map_x_153_add_exe = (_net_6902|_net_2910);
   assign  _add_map_x_153_p_reset = p_reset;
   assign  _add_map_x_153_m_clock = m_clock;
   assign  _add_map_x_152_moto_org_near = ((_net_6901)?data_in_org358:10'b0)|
    ((_net_2909)?data_in_org357:10'b0);
   assign  _add_map_x_152_moto_org_near1 = ((_net_6900)?data_in_org356:10'b0)|
    ((_net_2908)?data_in_org359:10'b0);
   assign  _add_map_x_152_moto_org_near2 = ((_net_6899)?data_in_org325:10'b0)|
    ((_net_2907)?data_in_org326:10'b0);
   assign  _add_map_x_152_moto_org_near3 = ((_net_6898)?data_in_org389:10'b0)|
    ((_net_2906)?data_in_org390:10'b0);
   assign  _add_map_x_152_moto_org = ((_net_6897)?data_in_org357:10'b0)|
    ((_net_2905)?data_in_org358:10'b0);
   assign  _add_map_x_152_sg_up = ((_net_6896)?sg_in358:2'b0)|
    ((_net_2904)?sg_in357:2'b0);
   assign  _add_map_x_152_sg_down = ((_net_6895)?sg_in325:2'b0)|
    ((_net_2903)?sg_in359:2'b0);
   assign  _add_map_x_152_sg_left = ((_net_6893)?sg_in389:2'b0)|
    ((_net_2901)?sg_in390:2'b0);
   assign  _add_map_x_152_sg_right = ((_net_6894)?sg_in356:2'b0)|
    ((_net_2902)?sg_in326:2'b0);
   assign  _add_map_x_152_wall_t_in = dig_w;
   assign  _add_map_x_152_moto = ((_net_6891)?data_in357:10'b0)|
    ((_net_2899)?data_in358:10'b0);
   assign  _add_map_x_152_up = ((_net_6890)?data_in358:10'b0)|
    ((_net_2898)?data_in357:10'b0);
   assign  _add_map_x_152_right = ((_net_6889)?data_in356:10'b0)|
    ((_net_2897)?data_in359:10'b0);
   assign  _add_map_x_152_down = ((_net_6888)?data_in325:10'b0)|
    ((_net_2896)?data_in326:10'b0);
   assign  _add_map_x_152_left = ((_net_6887)?data_in389:10'b0)|
    ((_net_2895)?data_in390:10'b0);
   assign  _add_map_x_152_start = start;
   assign  _add_map_x_152_goal = goal;
   assign  _add_map_x_152_now = ((_net_6884)?10'b0101100101:10'b0)|
    ((_net_2892)?10'b0101100110:10'b0);
   assign  _add_map_x_152_add_exe = (_net_6883|_net_2891);
   assign  _add_map_x_152_p_reset = p_reset;
   assign  _add_map_x_152_m_clock = m_clock;
   assign  _add_map_x_151_moto_org_near = ((_net_6882)?data_in_org356:10'b0)|
    ((_net_2890)?data_in_org355:10'b0);
   assign  _add_map_x_151_moto_org_near1 = ((_net_6881)?data_in_org354:10'b0)|
    ((_net_2889)?data_in_org357:10'b0);
   assign  _add_map_x_151_moto_org_near2 = ((_net_6880)?data_in_org323:10'b0)|
    ((_net_2888)?data_in_org324:10'b0);
   assign  _add_map_x_151_moto_org_near3 = ((_net_6879)?data_in_org387:10'b0)|
    ((_net_2887)?data_in_org388:10'b0);
   assign  _add_map_x_151_moto_org = ((_net_6878)?data_in_org355:10'b0)|
    ((_net_2886)?data_in_org356:10'b0);
   assign  _add_map_x_151_sg_up = ((_net_6877)?sg_in356:2'b0)|
    ((_net_2885)?sg_in355:2'b0);
   assign  _add_map_x_151_sg_down = ((_net_6876)?sg_in323:2'b0)|
    ((_net_2884)?sg_in357:2'b0);
   assign  _add_map_x_151_sg_left = ((_net_6874)?sg_in387:2'b0)|
    ((_net_2882)?sg_in388:2'b0);
   assign  _add_map_x_151_sg_right = ((_net_6875)?sg_in354:2'b0)|
    ((_net_2883)?sg_in324:2'b0);
   assign  _add_map_x_151_wall_t_in = dig_w;
   assign  _add_map_x_151_moto = ((_net_6872)?data_in355:10'b0)|
    ((_net_2880)?data_in356:10'b0);
   assign  _add_map_x_151_up = ((_net_6871)?data_in356:10'b0)|
    ((_net_2879)?data_in355:10'b0);
   assign  _add_map_x_151_right = ((_net_6870)?data_in354:10'b0)|
    ((_net_2878)?data_in357:10'b0);
   assign  _add_map_x_151_down = ((_net_6869)?data_in323:10'b0)|
    ((_net_2877)?data_in324:10'b0);
   assign  _add_map_x_151_left = ((_net_6868)?data_in387:10'b0)|
    ((_net_2876)?data_in388:10'b0);
   assign  _add_map_x_151_start = start;
   assign  _add_map_x_151_goal = goal;
   assign  _add_map_x_151_now = ((_net_6865)?10'b0101100011:10'b0)|
    ((_net_2873)?10'b0101100100:10'b0);
   assign  _add_map_x_151_add_exe = (_net_6864|_net_2872);
   assign  _add_map_x_151_p_reset = p_reset;
   assign  _add_map_x_151_m_clock = m_clock;
   assign  _add_map_x_150_moto_org_near = ((_net_6863)?data_in_org354:10'b0)|
    ((_net_2871)?data_in_org353:10'b0);
   assign  _add_map_x_150_moto_org_near1 = ((_net_6862)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2870)?data_in_org355:10'b0);
   assign  _add_map_x_150_moto_org_near2 = ((_net_6861)?data_in_org321:10'b0)|
    ((_net_2869)?data_in_org322:10'b0);
   assign  _add_map_x_150_moto_org_near3 = ((_net_6860)?data_in_org385:10'b0)|
    ((_net_2868)?data_in_org386:10'b0);
   assign  _add_map_x_150_moto_org = ((_net_6859)?data_in_org353:10'b0)|
    ((_net_2867)?data_in_org354:10'b0);
   assign  _add_map_x_150_sg_up = ((_net_6858)?sg_in354:2'b0)|
    ((_net_2866)?sg_in353:2'b0);
   assign  _add_map_x_150_sg_down = ((_net_6857)?sg_in321:2'b0)|
    ((_net_2865)?sg_in355:2'b0);
   assign  _add_map_x_150_sg_left = ((_net_6855)?sg_in385:2'b0)|
    ((_net_2863)?sg_in386:2'b0);
   assign  _add_map_x_150_sg_right = ((_net_6856)?3'b000:2'b0)|
    ((_net_2864)?sg_in322:2'b0);
   assign  _add_map_x_150_wall_t_in = dig_w;
   assign  _add_map_x_150_moto = ((_net_6853)?data_in353:10'b0)|
    ((_net_2861)?data_in354:10'b0);
   assign  _add_map_x_150_up = ((_net_6852)?data_in354:10'b0)|
    ((_net_2860)?data_in353:10'b0);
   assign  _add_map_x_150_right = ((_net_6851)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2859)?data_in355:10'b0);
   assign  _add_map_x_150_down = ((_net_6850)?data_in321:10'b0)|
    ((_net_2858)?data_in322:10'b0);
   assign  _add_map_x_150_left = ((_net_6849)?data_in385:10'b0)|
    ((_net_2857)?data_in386:10'b0);
   assign  _add_map_x_150_start = start;
   assign  _add_map_x_150_goal = goal;
   assign  _add_map_x_150_now = ((_net_6846)?10'b0101100001:10'b0)|
    ((_net_2854)?10'b0101100010:10'b0);
   assign  _add_map_x_150_add_exe = (_net_6845|_net_2853);
   assign  _add_map_x_150_p_reset = p_reset;
   assign  _add_map_x_150_m_clock = m_clock;
   assign  _add_map_x_149_moto_org_near = ((_net_6844)?data_in_org349:10'b0)|
    ((_net_2852)?data_in_org350:10'b0);
   assign  _add_map_x_149_moto_org_near1 = ((_net_6843)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2851)?data_in_org348:10'b0);
   assign  _add_map_x_149_moto_org_near2 = ((_net_6842)?data_in_org318:10'b0)|
    ((_net_2850)?data_in_org317:10'b0);
   assign  _add_map_x_149_moto_org_near3 = ((_net_6841)?data_in_org382:10'b0)|
    ((_net_2849)?data_in_org381:10'b0);
   assign  _add_map_x_149_moto_org = ((_net_6840)?data_in_org350:10'b0)|
    ((_net_2848)?data_in_org349:10'b0);
   assign  _add_map_x_149_sg_up = ((_net_6839)?sg_in349:2'b0)|
    ((_net_2847)?sg_in350:2'b0);
   assign  _add_map_x_149_sg_down = ((_net_6838)?3'b000:2'b0)|
    ((_net_2846)?sg_in348:2'b0);
   assign  _add_map_x_149_sg_left = ((_net_6836)?sg_in382:2'b0)|
    ((_net_2844)?sg_in381:2'b0);
   assign  _add_map_x_149_sg_right = ((_net_6837)?sg_in318:2'b0)|
    ((_net_2845)?sg_in317:2'b0);
   assign  _add_map_x_149_wall_t_in = dig_w;
   assign  _add_map_x_149_moto = ((_net_6834)?data_in350:10'b0)|
    ((_net_2842)?data_in349:10'b0);
   assign  _add_map_x_149_up = ((_net_6833)?data_in349:10'b0)|
    ((_net_2841)?data_in350:10'b0);
   assign  _add_map_x_149_right = ((_net_6832)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2840)?data_in348:10'b0);
   assign  _add_map_x_149_down = ((_net_6831)?data_in318:10'b0)|
    ((_net_2839)?data_in317:10'b0);
   assign  _add_map_x_149_left = ((_net_6830)?data_in382:10'b0)|
    ((_net_2838)?data_in381:10'b0);
   assign  _add_map_x_149_start = start;
   assign  _add_map_x_149_goal = goal;
   assign  _add_map_x_149_now = ((_net_6827)?10'b0101011110:10'b0)|
    ((_net_2835)?10'b0101011101:10'b0);
   assign  _add_map_x_149_add_exe = (_net_6826|_net_2834);
   assign  _add_map_x_149_p_reset = p_reset;
   assign  _add_map_x_149_m_clock = m_clock;
   assign  _add_map_x_148_moto_org_near = ((_net_6825)?data_in_org347:10'b0)|
    ((_net_2833)?data_in_org348:10'b0);
   assign  _add_map_x_148_moto_org_near1 = ((_net_6824)?data_in_org349:10'b0)|
    ((_net_2832)?data_in_org346:10'b0);
   assign  _add_map_x_148_moto_org_near2 = ((_net_6823)?data_in_org316:10'b0)|
    ((_net_2831)?data_in_org315:10'b0);
   assign  _add_map_x_148_moto_org_near3 = ((_net_6822)?data_in_org380:10'b0)|
    ((_net_2830)?data_in_org379:10'b0);
   assign  _add_map_x_148_moto_org = ((_net_6821)?data_in_org348:10'b0)|
    ((_net_2829)?data_in_org347:10'b0);
   assign  _add_map_x_148_sg_up = ((_net_6820)?sg_in347:2'b0)|
    ((_net_2828)?sg_in348:2'b0);
   assign  _add_map_x_148_sg_down = ((_net_6819)?sg_in349:2'b0)|
    ((_net_2827)?sg_in346:2'b0);
   assign  _add_map_x_148_sg_left = ((_net_6817)?sg_in380:2'b0)|
    ((_net_2825)?sg_in379:2'b0);
   assign  _add_map_x_148_sg_right = ((_net_6818)?sg_in316:2'b0)|
    ((_net_2826)?sg_in315:2'b0);
   assign  _add_map_x_148_wall_t_in = dig_w;
   assign  _add_map_x_148_moto = ((_net_6815)?data_in348:10'b0)|
    ((_net_2823)?data_in347:10'b0);
   assign  _add_map_x_148_up = ((_net_6814)?data_in347:10'b0)|
    ((_net_2822)?data_in348:10'b0);
   assign  _add_map_x_148_right = ((_net_6813)?data_in349:10'b0)|
    ((_net_2821)?data_in346:10'b0);
   assign  _add_map_x_148_down = ((_net_6812)?data_in316:10'b0)|
    ((_net_2820)?data_in315:10'b0);
   assign  _add_map_x_148_left = ((_net_6811)?data_in380:10'b0)|
    ((_net_2819)?data_in379:10'b0);
   assign  _add_map_x_148_start = start;
   assign  _add_map_x_148_goal = goal;
   assign  _add_map_x_148_now = ((_net_6808)?10'b0101011100:10'b0)|
    ((_net_2816)?10'b0101011011:10'b0);
   assign  _add_map_x_148_add_exe = (_net_6807|_net_2815);
   assign  _add_map_x_148_p_reset = p_reset;
   assign  _add_map_x_148_m_clock = m_clock;
   assign  _add_map_x_147_moto_org_near = ((_net_6806)?data_in_org345:10'b0)|
    ((_net_2814)?data_in_org346:10'b0);
   assign  _add_map_x_147_moto_org_near1 = ((_net_6805)?data_in_org347:10'b0)|
    ((_net_2813)?data_in_org344:10'b0);
   assign  _add_map_x_147_moto_org_near2 = ((_net_6804)?data_in_org314:10'b0)|
    ((_net_2812)?data_in_org313:10'b0);
   assign  _add_map_x_147_moto_org_near3 = ((_net_6803)?data_in_org378:10'b0)|
    ((_net_2811)?data_in_org377:10'b0);
   assign  _add_map_x_147_moto_org = ((_net_6802)?data_in_org346:10'b0)|
    ((_net_2810)?data_in_org345:10'b0);
   assign  _add_map_x_147_sg_up = ((_net_6801)?sg_in345:2'b0)|
    ((_net_2809)?sg_in346:2'b0);
   assign  _add_map_x_147_sg_down = ((_net_6800)?sg_in347:2'b0)|
    ((_net_2808)?sg_in344:2'b0);
   assign  _add_map_x_147_sg_left = ((_net_6798)?sg_in378:2'b0)|
    ((_net_2806)?sg_in377:2'b0);
   assign  _add_map_x_147_sg_right = ((_net_6799)?sg_in314:2'b0)|
    ((_net_2807)?sg_in313:2'b0);
   assign  _add_map_x_147_wall_t_in = dig_w;
   assign  _add_map_x_147_moto = ((_net_6796)?data_in346:10'b0)|
    ((_net_2804)?data_in345:10'b0);
   assign  _add_map_x_147_up = ((_net_6795)?data_in345:10'b0)|
    ((_net_2803)?data_in346:10'b0);
   assign  _add_map_x_147_right = ((_net_6794)?data_in347:10'b0)|
    ((_net_2802)?data_in344:10'b0);
   assign  _add_map_x_147_down = ((_net_6793)?data_in314:10'b0)|
    ((_net_2801)?data_in313:10'b0);
   assign  _add_map_x_147_left = ((_net_6792)?data_in378:10'b0)|
    ((_net_2800)?data_in377:10'b0);
   assign  _add_map_x_147_start = start;
   assign  _add_map_x_147_goal = goal;
   assign  _add_map_x_147_now = ((_net_6789)?10'b0101011010:10'b0)|
    ((_net_2797)?10'b0101011001:10'b0);
   assign  _add_map_x_147_add_exe = (_net_6788|_net_2796);
   assign  _add_map_x_147_p_reset = p_reset;
   assign  _add_map_x_147_m_clock = m_clock;
   assign  _add_map_x_146_moto_org_near = ((_net_6787)?data_in_org343:10'b0)|
    ((_net_2795)?data_in_org344:10'b0);
   assign  _add_map_x_146_moto_org_near1 = ((_net_6786)?data_in_org345:10'b0)|
    ((_net_2794)?data_in_org342:10'b0);
   assign  _add_map_x_146_moto_org_near2 = ((_net_6785)?data_in_org312:10'b0)|
    ((_net_2793)?data_in_org311:10'b0);
   assign  _add_map_x_146_moto_org_near3 = ((_net_6784)?data_in_org376:10'b0)|
    ((_net_2792)?data_in_org375:10'b0);
   assign  _add_map_x_146_moto_org = ((_net_6783)?data_in_org344:10'b0)|
    ((_net_2791)?data_in_org343:10'b0);
   assign  _add_map_x_146_sg_up = ((_net_6782)?sg_in343:2'b0)|
    ((_net_2790)?sg_in344:2'b0);
   assign  _add_map_x_146_sg_down = ((_net_6781)?sg_in345:2'b0)|
    ((_net_2789)?sg_in342:2'b0);
   assign  _add_map_x_146_sg_left = ((_net_6779)?sg_in376:2'b0)|
    ((_net_2787)?sg_in375:2'b0);
   assign  _add_map_x_146_sg_right = ((_net_6780)?sg_in312:2'b0)|
    ((_net_2788)?sg_in311:2'b0);
   assign  _add_map_x_146_wall_t_in = dig_w;
   assign  _add_map_x_146_moto = ((_net_6777)?data_in344:10'b0)|
    ((_net_2785)?data_in343:10'b0);
   assign  _add_map_x_146_up = ((_net_6776)?data_in343:10'b0)|
    ((_net_2784)?data_in344:10'b0);
   assign  _add_map_x_146_right = ((_net_6775)?data_in345:10'b0)|
    ((_net_2783)?data_in342:10'b0);
   assign  _add_map_x_146_down = ((_net_6774)?data_in312:10'b0)|
    ((_net_2782)?data_in311:10'b0);
   assign  _add_map_x_146_left = ((_net_6773)?data_in376:10'b0)|
    ((_net_2781)?data_in375:10'b0);
   assign  _add_map_x_146_start = start;
   assign  _add_map_x_146_goal = goal;
   assign  _add_map_x_146_now = ((_net_6770)?10'b0101011000:10'b0)|
    ((_net_2778)?10'b0101010111:10'b0);
   assign  _add_map_x_146_add_exe = (_net_6769|_net_2777);
   assign  _add_map_x_146_p_reset = p_reset;
   assign  _add_map_x_146_m_clock = m_clock;
   assign  _add_map_x_145_moto_org_near = ((_net_6768)?data_in_org341:10'b0)|
    ((_net_2776)?data_in_org342:10'b0);
   assign  _add_map_x_145_moto_org_near1 = ((_net_6767)?data_in_org343:10'b0)|
    ((_net_2775)?data_in_org340:10'b0);
   assign  _add_map_x_145_moto_org_near2 = ((_net_6766)?data_in_org310:10'b0)|
    ((_net_2774)?data_in_org309:10'b0);
   assign  _add_map_x_145_moto_org_near3 = ((_net_6765)?data_in_org374:10'b0)|
    ((_net_2773)?data_in_org373:10'b0);
   assign  _add_map_x_145_moto_org = ((_net_6764)?data_in_org342:10'b0)|
    ((_net_2772)?data_in_org341:10'b0);
   assign  _add_map_x_145_sg_up = ((_net_6763)?sg_in341:2'b0)|
    ((_net_2771)?sg_in342:2'b0);
   assign  _add_map_x_145_sg_down = ((_net_6762)?sg_in343:2'b0)|
    ((_net_2770)?sg_in340:2'b0);
   assign  _add_map_x_145_sg_left = ((_net_6760)?sg_in374:2'b0)|
    ((_net_2768)?sg_in373:2'b0);
   assign  _add_map_x_145_sg_right = ((_net_6761)?sg_in310:2'b0)|
    ((_net_2769)?sg_in309:2'b0);
   assign  _add_map_x_145_wall_t_in = dig_w;
   assign  _add_map_x_145_moto = ((_net_6758)?data_in342:10'b0)|
    ((_net_2766)?data_in341:10'b0);
   assign  _add_map_x_145_up = ((_net_6757)?data_in341:10'b0)|
    ((_net_2765)?data_in342:10'b0);
   assign  _add_map_x_145_right = ((_net_6756)?data_in343:10'b0)|
    ((_net_2764)?data_in340:10'b0);
   assign  _add_map_x_145_down = ((_net_6755)?data_in310:10'b0)|
    ((_net_2763)?data_in309:10'b0);
   assign  _add_map_x_145_left = ((_net_6754)?data_in374:10'b0)|
    ((_net_2762)?data_in373:10'b0);
   assign  _add_map_x_145_start = start;
   assign  _add_map_x_145_goal = goal;
   assign  _add_map_x_145_now = ((_net_6751)?10'b0101010110:10'b0)|
    ((_net_2759)?10'b0101010101:10'b0);
   assign  _add_map_x_145_add_exe = (_net_6750|_net_2758);
   assign  _add_map_x_145_p_reset = p_reset;
   assign  _add_map_x_145_m_clock = m_clock;
   assign  _add_map_x_144_moto_org_near = ((_net_6749)?data_in_org339:10'b0)|
    ((_net_2757)?data_in_org340:10'b0);
   assign  _add_map_x_144_moto_org_near1 = ((_net_6748)?data_in_org341:10'b0)|
    ((_net_2756)?data_in_org338:10'b0);
   assign  _add_map_x_144_moto_org_near2 = ((_net_6747)?data_in_org308:10'b0)|
    ((_net_2755)?data_in_org307:10'b0);
   assign  _add_map_x_144_moto_org_near3 = ((_net_6746)?data_in_org372:10'b0)|
    ((_net_2754)?data_in_org371:10'b0);
   assign  _add_map_x_144_moto_org = ((_net_6745)?data_in_org340:10'b0)|
    ((_net_2753)?data_in_org339:10'b0);
   assign  _add_map_x_144_sg_up = ((_net_6744)?sg_in339:2'b0)|
    ((_net_2752)?sg_in340:2'b0);
   assign  _add_map_x_144_sg_down = ((_net_6743)?sg_in341:2'b0)|
    ((_net_2751)?sg_in338:2'b0);
   assign  _add_map_x_144_sg_left = ((_net_6741)?sg_in372:2'b0)|
    ((_net_2749)?sg_in371:2'b0);
   assign  _add_map_x_144_sg_right = ((_net_6742)?sg_in308:2'b0)|
    ((_net_2750)?sg_in307:2'b0);
   assign  _add_map_x_144_wall_t_in = dig_w;
   assign  _add_map_x_144_moto = ((_net_6739)?data_in340:10'b0)|
    ((_net_2747)?data_in339:10'b0);
   assign  _add_map_x_144_up = ((_net_6738)?data_in339:10'b0)|
    ((_net_2746)?data_in340:10'b0);
   assign  _add_map_x_144_right = ((_net_6737)?data_in341:10'b0)|
    ((_net_2745)?data_in338:10'b0);
   assign  _add_map_x_144_down = ((_net_6736)?data_in308:10'b0)|
    ((_net_2744)?data_in307:10'b0);
   assign  _add_map_x_144_left = ((_net_6735)?data_in372:10'b0)|
    ((_net_2743)?data_in371:10'b0);
   assign  _add_map_x_144_start = start;
   assign  _add_map_x_144_goal = goal;
   assign  _add_map_x_144_now = ((_net_6732)?10'b0101010100:10'b0)|
    ((_net_2740)?10'b0101010011:10'b0);
   assign  _add_map_x_144_add_exe = (_net_6731|_net_2739);
   assign  _add_map_x_144_p_reset = p_reset;
   assign  _add_map_x_144_m_clock = m_clock;
   assign  _add_map_x_143_moto_org_near = ((_net_6730)?data_in_org337:10'b0)|
    ((_net_2738)?data_in_org338:10'b0);
   assign  _add_map_x_143_moto_org_near1 = ((_net_6729)?data_in_org339:10'b0)|
    ((_net_2737)?data_in_org336:10'b0);
   assign  _add_map_x_143_moto_org_near2 = ((_net_6728)?data_in_org306:10'b0)|
    ((_net_2736)?data_in_org305:10'b0);
   assign  _add_map_x_143_moto_org_near3 = ((_net_6727)?data_in_org370:10'b0)|
    ((_net_2735)?data_in_org369:10'b0);
   assign  _add_map_x_143_moto_org = ((_net_6726)?data_in_org338:10'b0)|
    ((_net_2734)?data_in_org337:10'b0);
   assign  _add_map_x_143_sg_up = ((_net_6725)?sg_in337:2'b0)|
    ((_net_2733)?sg_in338:2'b0);
   assign  _add_map_x_143_sg_down = ((_net_6724)?sg_in339:2'b0)|
    ((_net_2732)?sg_in336:2'b0);
   assign  _add_map_x_143_sg_left = ((_net_6722)?sg_in370:2'b0)|
    ((_net_2730)?sg_in369:2'b0);
   assign  _add_map_x_143_sg_right = ((_net_6723)?sg_in306:2'b0)|
    ((_net_2731)?sg_in305:2'b0);
   assign  _add_map_x_143_wall_t_in = dig_w;
   assign  _add_map_x_143_moto = ((_net_6720)?data_in338:10'b0)|
    ((_net_2728)?data_in337:10'b0);
   assign  _add_map_x_143_up = ((_net_6719)?data_in337:10'b0)|
    ((_net_2727)?data_in338:10'b0);
   assign  _add_map_x_143_right = ((_net_6718)?data_in339:10'b0)|
    ((_net_2726)?data_in336:10'b0);
   assign  _add_map_x_143_down = ((_net_6717)?data_in306:10'b0)|
    ((_net_2725)?data_in305:10'b0);
   assign  _add_map_x_143_left = ((_net_6716)?data_in370:10'b0)|
    ((_net_2724)?data_in369:10'b0);
   assign  _add_map_x_143_start = start;
   assign  _add_map_x_143_goal = goal;
   assign  _add_map_x_143_now = ((_net_6713)?10'b0101010010:10'b0)|
    ((_net_2721)?10'b0101010001:10'b0);
   assign  _add_map_x_143_add_exe = (_net_6712|_net_2720);
   assign  _add_map_x_143_p_reset = p_reset;
   assign  _add_map_x_143_m_clock = m_clock;
   assign  _add_map_x_142_moto_org_near = ((_net_6711)?data_in_org335:10'b0)|
    ((_net_2719)?data_in_org336:10'b0);
   assign  _add_map_x_142_moto_org_near1 = ((_net_6710)?data_in_org337:10'b0)|
    ((_net_2718)?data_in_org334:10'b0);
   assign  _add_map_x_142_moto_org_near2 = ((_net_6709)?data_in_org304:10'b0)|
    ((_net_2717)?data_in_org303:10'b0);
   assign  _add_map_x_142_moto_org_near3 = ((_net_6708)?data_in_org368:10'b0)|
    ((_net_2716)?data_in_org367:10'b0);
   assign  _add_map_x_142_moto_org = ((_net_6707)?data_in_org336:10'b0)|
    ((_net_2715)?data_in_org335:10'b0);
   assign  _add_map_x_142_sg_up = ((_net_6706)?sg_in335:2'b0)|
    ((_net_2714)?sg_in336:2'b0);
   assign  _add_map_x_142_sg_down = ((_net_6705)?sg_in337:2'b0)|
    ((_net_2713)?sg_in334:2'b0);
   assign  _add_map_x_142_sg_left = ((_net_6703)?sg_in368:2'b0)|
    ((_net_2711)?sg_in367:2'b0);
   assign  _add_map_x_142_sg_right = ((_net_6704)?sg_in304:2'b0)|
    ((_net_2712)?sg_in303:2'b0);
   assign  _add_map_x_142_wall_t_in = dig_w;
   assign  _add_map_x_142_moto = ((_net_6701)?data_in336:10'b0)|
    ((_net_2709)?data_in335:10'b0);
   assign  _add_map_x_142_up = ((_net_6700)?data_in335:10'b0)|
    ((_net_2708)?data_in336:10'b0);
   assign  _add_map_x_142_right = ((_net_6699)?data_in337:10'b0)|
    ((_net_2707)?data_in334:10'b0);
   assign  _add_map_x_142_down = ((_net_6698)?data_in304:10'b0)|
    ((_net_2706)?data_in303:10'b0);
   assign  _add_map_x_142_left = ((_net_6697)?data_in368:10'b0)|
    ((_net_2705)?data_in367:10'b0);
   assign  _add_map_x_142_start = start;
   assign  _add_map_x_142_goal = goal;
   assign  _add_map_x_142_now = ((_net_6694)?10'b0101010000:10'b0)|
    ((_net_2702)?10'b0101001111:10'b0);
   assign  _add_map_x_142_add_exe = (_net_6693|_net_2701);
   assign  _add_map_x_142_p_reset = p_reset;
   assign  _add_map_x_142_m_clock = m_clock;
   assign  _add_map_x_141_moto_org_near = ((_net_6692)?data_in_org333:10'b0)|
    ((_net_2700)?data_in_org334:10'b0);
   assign  _add_map_x_141_moto_org_near1 = ((_net_6691)?data_in_org335:10'b0)|
    ((_net_2699)?data_in_org332:10'b0);
   assign  _add_map_x_141_moto_org_near2 = ((_net_6690)?data_in_org302:10'b0)|
    ((_net_2698)?data_in_org301:10'b0);
   assign  _add_map_x_141_moto_org_near3 = ((_net_6689)?data_in_org366:10'b0)|
    ((_net_2697)?data_in_org365:10'b0);
   assign  _add_map_x_141_moto_org = ((_net_6688)?data_in_org334:10'b0)|
    ((_net_2696)?data_in_org333:10'b0);
   assign  _add_map_x_141_sg_up = ((_net_6687)?sg_in333:2'b0)|
    ((_net_2695)?sg_in334:2'b0);
   assign  _add_map_x_141_sg_down = ((_net_6686)?sg_in335:2'b0)|
    ((_net_2694)?sg_in332:2'b0);
   assign  _add_map_x_141_sg_left = ((_net_6684)?sg_in366:2'b0)|
    ((_net_2692)?sg_in365:2'b0);
   assign  _add_map_x_141_sg_right = ((_net_6685)?sg_in302:2'b0)|
    ((_net_2693)?sg_in301:2'b0);
   assign  _add_map_x_141_wall_t_in = dig_w;
   assign  _add_map_x_141_moto = ((_net_6682)?data_in334:10'b0)|
    ((_net_2690)?data_in333:10'b0);
   assign  _add_map_x_141_up = ((_net_6681)?data_in333:10'b0)|
    ((_net_2689)?data_in334:10'b0);
   assign  _add_map_x_141_right = ((_net_6680)?data_in335:10'b0)|
    ((_net_2688)?data_in332:10'b0);
   assign  _add_map_x_141_down = ((_net_6679)?data_in302:10'b0)|
    ((_net_2687)?data_in301:10'b0);
   assign  _add_map_x_141_left = ((_net_6678)?data_in366:10'b0)|
    ((_net_2686)?data_in365:10'b0);
   assign  _add_map_x_141_start = start;
   assign  _add_map_x_141_goal = goal;
   assign  _add_map_x_141_now = ((_net_6675)?10'b0101001110:10'b0)|
    ((_net_2683)?10'b0101001101:10'b0);
   assign  _add_map_x_141_add_exe = (_net_6674|_net_2682);
   assign  _add_map_x_141_p_reset = p_reset;
   assign  _add_map_x_141_m_clock = m_clock;
   assign  _add_map_x_140_moto_org_near = ((_net_6673)?data_in_org331:10'b0)|
    ((_net_2681)?data_in_org332:10'b0);
   assign  _add_map_x_140_moto_org_near1 = ((_net_6672)?data_in_org333:10'b0)|
    ((_net_2680)?data_in_org330:10'b0);
   assign  _add_map_x_140_moto_org_near2 = ((_net_6671)?data_in_org300:10'b0)|
    ((_net_2679)?data_in_org299:10'b0);
   assign  _add_map_x_140_moto_org_near3 = ((_net_6670)?data_in_org364:10'b0)|
    ((_net_2678)?data_in_org363:10'b0);
   assign  _add_map_x_140_moto_org = ((_net_6669)?data_in_org332:10'b0)|
    ((_net_2677)?data_in_org331:10'b0);
   assign  _add_map_x_140_sg_up = ((_net_6668)?sg_in331:2'b0)|
    ((_net_2676)?sg_in332:2'b0);
   assign  _add_map_x_140_sg_down = ((_net_6667)?sg_in333:2'b0)|
    ((_net_2675)?sg_in330:2'b0);
   assign  _add_map_x_140_sg_left = ((_net_6665)?sg_in364:2'b0)|
    ((_net_2673)?sg_in363:2'b0);
   assign  _add_map_x_140_sg_right = ((_net_6666)?sg_in300:2'b0)|
    ((_net_2674)?sg_in299:2'b0);
   assign  _add_map_x_140_wall_t_in = dig_w;
   assign  _add_map_x_140_moto = ((_net_6663)?data_in332:10'b0)|
    ((_net_2671)?data_in331:10'b0);
   assign  _add_map_x_140_up = ((_net_6662)?data_in331:10'b0)|
    ((_net_2670)?data_in332:10'b0);
   assign  _add_map_x_140_right = ((_net_6661)?data_in333:10'b0)|
    ((_net_2669)?data_in330:10'b0);
   assign  _add_map_x_140_down = ((_net_6660)?data_in300:10'b0)|
    ((_net_2668)?data_in299:10'b0);
   assign  _add_map_x_140_left = ((_net_6659)?data_in364:10'b0)|
    ((_net_2667)?data_in363:10'b0);
   assign  _add_map_x_140_start = start;
   assign  _add_map_x_140_goal = goal;
   assign  _add_map_x_140_now = ((_net_6656)?10'b0101001100:10'b0)|
    ((_net_2664)?10'b0101001011:10'b0);
   assign  _add_map_x_140_add_exe = (_net_6655|_net_2663);
   assign  _add_map_x_140_p_reset = p_reset;
   assign  _add_map_x_140_m_clock = m_clock;
   assign  _add_map_x_139_moto_org_near = ((_net_6654)?data_in_org329:10'b0)|
    ((_net_2662)?data_in_org330:10'b0);
   assign  _add_map_x_139_moto_org_near1 = ((_net_6653)?data_in_org331:10'b0)|
    ((_net_2661)?data_in_org328:10'b0);
   assign  _add_map_x_139_moto_org_near2 = ((_net_6652)?data_in_org298:10'b0)|
    ((_net_2660)?data_in_org297:10'b0);
   assign  _add_map_x_139_moto_org_near3 = ((_net_6651)?data_in_org362:10'b0)|
    ((_net_2659)?data_in_org361:10'b0);
   assign  _add_map_x_139_moto_org = ((_net_6650)?data_in_org330:10'b0)|
    ((_net_2658)?data_in_org329:10'b0);
   assign  _add_map_x_139_sg_up = ((_net_6649)?sg_in329:2'b0)|
    ((_net_2657)?sg_in330:2'b0);
   assign  _add_map_x_139_sg_down = ((_net_6648)?sg_in331:2'b0)|
    ((_net_2656)?sg_in328:2'b0);
   assign  _add_map_x_139_sg_left = ((_net_6646)?sg_in362:2'b0)|
    ((_net_2654)?sg_in361:2'b0);
   assign  _add_map_x_139_sg_right = ((_net_6647)?sg_in298:2'b0)|
    ((_net_2655)?sg_in297:2'b0);
   assign  _add_map_x_139_wall_t_in = dig_w;
   assign  _add_map_x_139_moto = ((_net_6644)?data_in330:10'b0)|
    ((_net_2652)?data_in329:10'b0);
   assign  _add_map_x_139_up = ((_net_6643)?data_in329:10'b0)|
    ((_net_2651)?data_in330:10'b0);
   assign  _add_map_x_139_right = ((_net_6642)?data_in331:10'b0)|
    ((_net_2650)?data_in328:10'b0);
   assign  _add_map_x_139_down = ((_net_6641)?data_in298:10'b0)|
    ((_net_2649)?data_in297:10'b0);
   assign  _add_map_x_139_left = ((_net_6640)?data_in362:10'b0)|
    ((_net_2648)?data_in361:10'b0);
   assign  _add_map_x_139_start = start;
   assign  _add_map_x_139_goal = goal;
   assign  _add_map_x_139_now = ((_net_6637)?10'b0101001010:10'b0)|
    ((_net_2645)?10'b0101001001:10'b0);
   assign  _add_map_x_139_add_exe = (_net_6636|_net_2644);
   assign  _add_map_x_139_p_reset = p_reset;
   assign  _add_map_x_139_m_clock = m_clock;
   assign  _add_map_x_138_moto_org_near = ((_net_6635)?data_in_org327:10'b0)|
    ((_net_2643)?data_in_org328:10'b0);
   assign  _add_map_x_138_moto_org_near1 = ((_net_6634)?data_in_org329:10'b0)|
    ((_net_2642)?data_in_org326:10'b0);
   assign  _add_map_x_138_moto_org_near2 = ((_net_6633)?data_in_org296:10'b0)|
    ((_net_2641)?data_in_org295:10'b0);
   assign  _add_map_x_138_moto_org_near3 = ((_net_6632)?data_in_org360:10'b0)|
    ((_net_2640)?data_in_org359:10'b0);
   assign  _add_map_x_138_moto_org = ((_net_6631)?data_in_org328:10'b0)|
    ((_net_2639)?data_in_org327:10'b0);
   assign  _add_map_x_138_sg_up = ((_net_6630)?sg_in327:2'b0)|
    ((_net_2638)?sg_in328:2'b0);
   assign  _add_map_x_138_sg_down = ((_net_6629)?sg_in329:2'b0)|
    ((_net_2637)?sg_in326:2'b0);
   assign  _add_map_x_138_sg_left = ((_net_6627)?sg_in360:2'b0)|
    ((_net_2635)?sg_in359:2'b0);
   assign  _add_map_x_138_sg_right = ((_net_6628)?sg_in296:2'b0)|
    ((_net_2636)?sg_in295:2'b0);
   assign  _add_map_x_138_wall_t_in = dig_w;
   assign  _add_map_x_138_moto = ((_net_6625)?data_in328:10'b0)|
    ((_net_2633)?data_in327:10'b0);
   assign  _add_map_x_138_up = ((_net_6624)?data_in327:10'b0)|
    ((_net_2632)?data_in328:10'b0);
   assign  _add_map_x_138_right = ((_net_6623)?data_in329:10'b0)|
    ((_net_2631)?data_in326:10'b0);
   assign  _add_map_x_138_down = ((_net_6622)?data_in296:10'b0)|
    ((_net_2630)?data_in295:10'b0);
   assign  _add_map_x_138_left = ((_net_6621)?data_in360:10'b0)|
    ((_net_2629)?data_in359:10'b0);
   assign  _add_map_x_138_start = start;
   assign  _add_map_x_138_goal = goal;
   assign  _add_map_x_138_now = ((_net_6618)?10'b0101001000:10'b0)|
    ((_net_2626)?10'b0101000111:10'b0);
   assign  _add_map_x_138_add_exe = (_net_6617|_net_2625);
   assign  _add_map_x_138_p_reset = p_reset;
   assign  _add_map_x_138_m_clock = m_clock;
   assign  _add_map_x_137_moto_org_near = ((_net_6616)?data_in_org325:10'b0)|
    ((_net_2624)?data_in_org326:10'b0);
   assign  _add_map_x_137_moto_org_near1 = ((_net_6615)?data_in_org327:10'b0)|
    ((_net_2623)?data_in_org324:10'b0);
   assign  _add_map_x_137_moto_org_near2 = ((_net_6614)?data_in_org294:10'b0)|
    ((_net_2622)?data_in_org293:10'b0);
   assign  _add_map_x_137_moto_org_near3 = ((_net_6613)?data_in_org358:10'b0)|
    ((_net_2621)?data_in_org357:10'b0);
   assign  _add_map_x_137_moto_org = ((_net_6612)?data_in_org326:10'b0)|
    ((_net_2620)?data_in_org325:10'b0);
   assign  _add_map_x_137_sg_up = ((_net_6611)?sg_in325:2'b0)|
    ((_net_2619)?sg_in326:2'b0);
   assign  _add_map_x_137_sg_down = ((_net_6610)?sg_in327:2'b0)|
    ((_net_2618)?sg_in324:2'b0);
   assign  _add_map_x_137_sg_left = ((_net_6608)?sg_in358:2'b0)|
    ((_net_2616)?sg_in357:2'b0);
   assign  _add_map_x_137_sg_right = ((_net_6609)?sg_in294:2'b0)|
    ((_net_2617)?sg_in293:2'b0);
   assign  _add_map_x_137_wall_t_in = dig_w;
   assign  _add_map_x_137_moto = ((_net_6606)?data_in326:10'b0)|
    ((_net_2614)?data_in325:10'b0);
   assign  _add_map_x_137_up = ((_net_6605)?data_in325:10'b0)|
    ((_net_2613)?data_in326:10'b0);
   assign  _add_map_x_137_right = ((_net_6604)?data_in327:10'b0)|
    ((_net_2612)?data_in324:10'b0);
   assign  _add_map_x_137_down = ((_net_6603)?data_in294:10'b0)|
    ((_net_2611)?data_in293:10'b0);
   assign  _add_map_x_137_left = ((_net_6602)?data_in358:10'b0)|
    ((_net_2610)?data_in357:10'b0);
   assign  _add_map_x_137_start = start;
   assign  _add_map_x_137_goal = goal;
   assign  _add_map_x_137_now = ((_net_6599)?10'b0101000110:10'b0)|
    ((_net_2607)?10'b0101000101:10'b0);
   assign  _add_map_x_137_add_exe = (_net_6598|_net_2606);
   assign  _add_map_x_137_p_reset = p_reset;
   assign  _add_map_x_137_m_clock = m_clock;
   assign  _add_map_x_136_moto_org_near = ((_net_6597)?data_in_org323:10'b0)|
    ((_net_2605)?data_in_org324:10'b0);
   assign  _add_map_x_136_moto_org_near1 = ((_net_6596)?data_in_org325:10'b0)|
    ((_net_2604)?data_in_org322:10'b0);
   assign  _add_map_x_136_moto_org_near2 = ((_net_6595)?data_in_org292:10'b0)|
    ((_net_2603)?data_in_org291:10'b0);
   assign  _add_map_x_136_moto_org_near3 = ((_net_6594)?data_in_org356:10'b0)|
    ((_net_2602)?data_in_org355:10'b0);
   assign  _add_map_x_136_moto_org = ((_net_6593)?data_in_org324:10'b0)|
    ((_net_2601)?data_in_org323:10'b0);
   assign  _add_map_x_136_sg_up = ((_net_6592)?sg_in323:2'b0)|
    ((_net_2600)?sg_in324:2'b0);
   assign  _add_map_x_136_sg_down = ((_net_6591)?sg_in325:2'b0)|
    ((_net_2599)?sg_in322:2'b0);
   assign  _add_map_x_136_sg_left = ((_net_6589)?sg_in356:2'b0)|
    ((_net_2597)?sg_in355:2'b0);
   assign  _add_map_x_136_sg_right = ((_net_6590)?sg_in292:2'b0)|
    ((_net_2598)?sg_in291:2'b0);
   assign  _add_map_x_136_wall_t_in = dig_w;
   assign  _add_map_x_136_moto = ((_net_6587)?data_in324:10'b0)|
    ((_net_2595)?data_in323:10'b0);
   assign  _add_map_x_136_up = ((_net_6586)?data_in323:10'b0)|
    ((_net_2594)?data_in324:10'b0);
   assign  _add_map_x_136_right = ((_net_6585)?data_in325:10'b0)|
    ((_net_2593)?data_in322:10'b0);
   assign  _add_map_x_136_down = ((_net_6584)?data_in292:10'b0)|
    ((_net_2592)?data_in291:10'b0);
   assign  _add_map_x_136_left = ((_net_6583)?data_in356:10'b0)|
    ((_net_2591)?data_in355:10'b0);
   assign  _add_map_x_136_start = start;
   assign  _add_map_x_136_goal = goal;
   assign  _add_map_x_136_now = ((_net_6580)?10'b0101000100:10'b0)|
    ((_net_2588)?10'b0101000011:10'b0);
   assign  _add_map_x_136_add_exe = (_net_6579|_net_2587);
   assign  _add_map_x_136_p_reset = p_reset;
   assign  _add_map_x_136_m_clock = m_clock;
   assign  _add_map_x_135_moto_org_near = ((_net_6578)?data_in_org321:10'b0)|
    ((_net_2586)?data_in_org322:10'b0);
   assign  _add_map_x_135_moto_org_near1 = ((_net_6577)?data_in_org323:10'b0)|
    ((_net_2585)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_135_moto_org_near2 = ((_net_6576)?data_in_org290:10'b0)|
    ((_net_2584)?data_in_org289:10'b0);
   assign  _add_map_x_135_moto_org_near3 = ((_net_6575)?data_in_org354:10'b0)|
    ((_net_2583)?data_in_org353:10'b0);
   assign  _add_map_x_135_moto_org = ((_net_6574)?data_in_org322:10'b0)|
    ((_net_2582)?data_in_org321:10'b0);
   assign  _add_map_x_135_sg_up = ((_net_6573)?sg_in321:2'b0)|
    ((_net_2581)?sg_in322:2'b0);
   assign  _add_map_x_135_sg_down = ((_net_6572)?sg_in323:2'b0)|
    ((_net_2580)?3'b000:2'b0);
   assign  _add_map_x_135_sg_left = ((_net_6570)?sg_in354:2'b0)|
    ((_net_2578)?sg_in353:2'b0);
   assign  _add_map_x_135_sg_right = ((_net_6571)?sg_in290:2'b0)|
    ((_net_2579)?sg_in289:2'b0);
   assign  _add_map_x_135_wall_t_in = dig_w;
   assign  _add_map_x_135_moto = ((_net_6568)?data_in322:10'b0)|
    ((_net_2576)?data_in321:10'b0);
   assign  _add_map_x_135_up = ((_net_6567)?data_in321:10'b0)|
    ((_net_2575)?data_in322:10'b0);
   assign  _add_map_x_135_right = ((_net_6566)?data_in323:10'b0)|
    ((_net_2574)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_135_down = ((_net_6565)?data_in290:10'b0)|
    ((_net_2573)?data_in289:10'b0);
   assign  _add_map_x_135_left = ((_net_6564)?data_in354:10'b0)|
    ((_net_2572)?data_in353:10'b0);
   assign  _add_map_x_135_start = start;
   assign  _add_map_x_135_goal = goal;
   assign  _add_map_x_135_now = ((_net_6561)?10'b0101000010:10'b0)|
    ((_net_2569)?10'b0101000001:10'b0);
   assign  _add_map_x_135_add_exe = (_net_6560|_net_2568);
   assign  _add_map_x_135_p_reset = p_reset;
   assign  _add_map_x_135_m_clock = m_clock;
   assign  _add_map_x_134_moto_org_near = ((_net_6559)?data_in_org318:10'b0)|
    ((_net_2567)?data_in_org317:10'b0);
   assign  _add_map_x_134_moto_org_near1 = ((_net_6558)?data_in_org316:10'b0)|
    ((_net_2566)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_134_moto_org_near2 = ((_net_6557)?data_in_org285:10'b0)|
    ((_net_2565)?data_in_org286:10'b0);
   assign  _add_map_x_134_moto_org_near3 = ((_net_6556)?data_in_org349:10'b0)|
    ((_net_2564)?data_in_org350:10'b0);
   assign  _add_map_x_134_moto_org = ((_net_6555)?data_in_org317:10'b0)|
    ((_net_2563)?data_in_org318:10'b0);
   assign  _add_map_x_134_sg_up = ((_net_6554)?sg_in318:2'b0)|
    ((_net_2562)?sg_in317:2'b0);
   assign  _add_map_x_134_sg_down = ((_net_6553)?sg_in285:2'b0)|
    ((_net_2561)?3'b000:2'b0);
   assign  _add_map_x_134_sg_left = ((_net_6551)?sg_in349:2'b0)|
    ((_net_2559)?sg_in350:2'b0);
   assign  _add_map_x_134_sg_right = ((_net_6552)?sg_in316:2'b0)|
    ((_net_2560)?sg_in286:2'b0);
   assign  _add_map_x_134_wall_t_in = dig_w;
   assign  _add_map_x_134_moto = ((_net_6549)?data_in317:10'b0)|
    ((_net_2557)?data_in318:10'b0);
   assign  _add_map_x_134_up = ((_net_6548)?data_in318:10'b0)|
    ((_net_2556)?data_in317:10'b0);
   assign  _add_map_x_134_right = ((_net_6547)?data_in316:10'b0)|
    ((_net_2555)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_134_down = ((_net_6546)?data_in285:10'b0)|
    ((_net_2554)?data_in286:10'b0);
   assign  _add_map_x_134_left = ((_net_6545)?data_in349:10'b0)|
    ((_net_2553)?data_in350:10'b0);
   assign  _add_map_x_134_start = start;
   assign  _add_map_x_134_goal = goal;
   assign  _add_map_x_134_now = ((_net_6542)?10'b0100111101:10'b0)|
    ((_net_2550)?10'b0100111110:10'b0);
   assign  _add_map_x_134_add_exe = (_net_6541|_net_2549);
   assign  _add_map_x_134_p_reset = p_reset;
   assign  _add_map_x_134_m_clock = m_clock;
   assign  _add_map_x_133_moto_org_near = ((_net_6540)?data_in_org316:10'b0)|
    ((_net_2548)?data_in_org315:10'b0);
   assign  _add_map_x_133_moto_org_near1 = ((_net_6539)?data_in_org314:10'b0)|
    ((_net_2547)?data_in_org317:10'b0);
   assign  _add_map_x_133_moto_org_near2 = ((_net_6538)?data_in_org283:10'b0)|
    ((_net_2546)?data_in_org284:10'b0);
   assign  _add_map_x_133_moto_org_near3 = ((_net_6537)?data_in_org347:10'b0)|
    ((_net_2545)?data_in_org348:10'b0);
   assign  _add_map_x_133_moto_org = ((_net_6536)?data_in_org315:10'b0)|
    ((_net_2544)?data_in_org316:10'b0);
   assign  _add_map_x_133_sg_up = ((_net_6535)?sg_in316:2'b0)|
    ((_net_2543)?sg_in315:2'b0);
   assign  _add_map_x_133_sg_down = ((_net_6534)?sg_in283:2'b0)|
    ((_net_2542)?sg_in317:2'b0);
   assign  _add_map_x_133_sg_left = ((_net_6532)?sg_in347:2'b0)|
    ((_net_2540)?sg_in348:2'b0);
   assign  _add_map_x_133_sg_right = ((_net_6533)?sg_in314:2'b0)|
    ((_net_2541)?sg_in284:2'b0);
   assign  _add_map_x_133_wall_t_in = dig_w;
   assign  _add_map_x_133_moto = ((_net_6530)?data_in315:10'b0)|
    ((_net_2538)?data_in316:10'b0);
   assign  _add_map_x_133_up = ((_net_6529)?data_in316:10'b0)|
    ((_net_2537)?data_in315:10'b0);
   assign  _add_map_x_133_right = ((_net_6528)?data_in314:10'b0)|
    ((_net_2536)?data_in317:10'b0);
   assign  _add_map_x_133_down = ((_net_6527)?data_in283:10'b0)|
    ((_net_2535)?data_in284:10'b0);
   assign  _add_map_x_133_left = ((_net_6526)?data_in347:10'b0)|
    ((_net_2534)?data_in348:10'b0);
   assign  _add_map_x_133_start = start;
   assign  _add_map_x_133_goal = goal;
   assign  _add_map_x_133_now = ((_net_6523)?10'b0100111011:10'b0)|
    ((_net_2531)?10'b0100111100:10'b0);
   assign  _add_map_x_133_add_exe = (_net_6522|_net_2530);
   assign  _add_map_x_133_p_reset = p_reset;
   assign  _add_map_x_133_m_clock = m_clock;
   assign  _add_map_x_132_moto_org_near = ((_net_6521)?data_in_org314:10'b0)|
    ((_net_2529)?data_in_org313:10'b0);
   assign  _add_map_x_132_moto_org_near1 = ((_net_6520)?data_in_org312:10'b0)|
    ((_net_2528)?data_in_org315:10'b0);
   assign  _add_map_x_132_moto_org_near2 = ((_net_6519)?data_in_org281:10'b0)|
    ((_net_2527)?data_in_org282:10'b0);
   assign  _add_map_x_132_moto_org_near3 = ((_net_6518)?data_in_org345:10'b0)|
    ((_net_2526)?data_in_org346:10'b0);
   assign  _add_map_x_132_moto_org = ((_net_6517)?data_in_org313:10'b0)|
    ((_net_2525)?data_in_org314:10'b0);
   assign  _add_map_x_132_sg_up = ((_net_6516)?sg_in314:2'b0)|
    ((_net_2524)?sg_in313:2'b0);
   assign  _add_map_x_132_sg_down = ((_net_6515)?sg_in281:2'b0)|
    ((_net_2523)?sg_in315:2'b0);
   assign  _add_map_x_132_sg_left = ((_net_6513)?sg_in345:2'b0)|
    ((_net_2521)?sg_in346:2'b0);
   assign  _add_map_x_132_sg_right = ((_net_6514)?sg_in312:2'b0)|
    ((_net_2522)?sg_in282:2'b0);
   assign  _add_map_x_132_wall_t_in = dig_w;
   assign  _add_map_x_132_moto = ((_net_6511)?data_in313:10'b0)|
    ((_net_2519)?data_in314:10'b0);
   assign  _add_map_x_132_up = ((_net_6510)?data_in314:10'b0)|
    ((_net_2518)?data_in313:10'b0);
   assign  _add_map_x_132_right = ((_net_6509)?data_in312:10'b0)|
    ((_net_2517)?data_in315:10'b0);
   assign  _add_map_x_132_down = ((_net_6508)?data_in281:10'b0)|
    ((_net_2516)?data_in282:10'b0);
   assign  _add_map_x_132_left = ((_net_6507)?data_in345:10'b0)|
    ((_net_2515)?data_in346:10'b0);
   assign  _add_map_x_132_start = start;
   assign  _add_map_x_132_goal = goal;
   assign  _add_map_x_132_now = ((_net_6504)?10'b0100111001:10'b0)|
    ((_net_2512)?10'b0100111010:10'b0);
   assign  _add_map_x_132_add_exe = (_net_6503|_net_2511);
   assign  _add_map_x_132_p_reset = p_reset;
   assign  _add_map_x_132_m_clock = m_clock;
   assign  _add_map_x_131_moto_org_near = ((_net_6502)?data_in_org312:10'b0)|
    ((_net_2510)?data_in_org311:10'b0);
   assign  _add_map_x_131_moto_org_near1 = ((_net_6501)?data_in_org310:10'b0)|
    ((_net_2509)?data_in_org313:10'b0);
   assign  _add_map_x_131_moto_org_near2 = ((_net_6500)?data_in_org279:10'b0)|
    ((_net_2508)?data_in_org280:10'b0);
   assign  _add_map_x_131_moto_org_near3 = ((_net_6499)?data_in_org343:10'b0)|
    ((_net_2507)?data_in_org344:10'b0);
   assign  _add_map_x_131_moto_org = ((_net_6498)?data_in_org311:10'b0)|
    ((_net_2506)?data_in_org312:10'b0);
   assign  _add_map_x_131_sg_up = ((_net_6497)?sg_in312:2'b0)|
    ((_net_2505)?sg_in311:2'b0);
   assign  _add_map_x_131_sg_down = ((_net_6496)?sg_in279:2'b0)|
    ((_net_2504)?sg_in313:2'b0);
   assign  _add_map_x_131_sg_left = ((_net_6494)?sg_in343:2'b0)|
    ((_net_2502)?sg_in344:2'b0);
   assign  _add_map_x_131_sg_right = ((_net_6495)?sg_in310:2'b0)|
    ((_net_2503)?sg_in280:2'b0);
   assign  _add_map_x_131_wall_t_in = dig_w;
   assign  _add_map_x_131_moto = ((_net_6492)?data_in311:10'b0)|
    ((_net_2500)?data_in312:10'b0);
   assign  _add_map_x_131_up = ((_net_6491)?data_in312:10'b0)|
    ((_net_2499)?data_in311:10'b0);
   assign  _add_map_x_131_right = ((_net_6490)?data_in310:10'b0)|
    ((_net_2498)?data_in313:10'b0);
   assign  _add_map_x_131_down = ((_net_6489)?data_in279:10'b0)|
    ((_net_2497)?data_in280:10'b0);
   assign  _add_map_x_131_left = ((_net_6488)?data_in343:10'b0)|
    ((_net_2496)?data_in344:10'b0);
   assign  _add_map_x_131_start = start;
   assign  _add_map_x_131_goal = goal;
   assign  _add_map_x_131_now = ((_net_6485)?10'b0100110111:10'b0)|
    ((_net_2493)?10'b0100111000:10'b0);
   assign  _add_map_x_131_add_exe = (_net_6484|_net_2492);
   assign  _add_map_x_131_p_reset = p_reset;
   assign  _add_map_x_131_m_clock = m_clock;
   assign  _add_map_x_130_moto_org_near = ((_net_6483)?data_in_org310:10'b0)|
    ((_net_2491)?data_in_org309:10'b0);
   assign  _add_map_x_130_moto_org_near1 = ((_net_6482)?data_in_org308:10'b0)|
    ((_net_2490)?data_in_org311:10'b0);
   assign  _add_map_x_130_moto_org_near2 = ((_net_6481)?data_in_org277:10'b0)|
    ((_net_2489)?data_in_org278:10'b0);
   assign  _add_map_x_130_moto_org_near3 = ((_net_6480)?data_in_org341:10'b0)|
    ((_net_2488)?data_in_org342:10'b0);
   assign  _add_map_x_130_moto_org = ((_net_6479)?data_in_org309:10'b0)|
    ((_net_2487)?data_in_org310:10'b0);
   assign  _add_map_x_130_sg_up = ((_net_6478)?sg_in310:2'b0)|
    ((_net_2486)?sg_in309:2'b0);
   assign  _add_map_x_130_sg_down = ((_net_6477)?sg_in277:2'b0)|
    ((_net_2485)?sg_in311:2'b0);
   assign  _add_map_x_130_sg_left = ((_net_6475)?sg_in341:2'b0)|
    ((_net_2483)?sg_in342:2'b0);
   assign  _add_map_x_130_sg_right = ((_net_6476)?sg_in308:2'b0)|
    ((_net_2484)?sg_in278:2'b0);
   assign  _add_map_x_130_wall_t_in = dig_w;
   assign  _add_map_x_130_moto = ((_net_6473)?data_in309:10'b0)|
    ((_net_2481)?data_in310:10'b0);
   assign  _add_map_x_130_up = ((_net_6472)?data_in310:10'b0)|
    ((_net_2480)?data_in309:10'b0);
   assign  _add_map_x_130_right = ((_net_6471)?data_in308:10'b0)|
    ((_net_2479)?data_in311:10'b0);
   assign  _add_map_x_130_down = ((_net_6470)?data_in277:10'b0)|
    ((_net_2478)?data_in278:10'b0);
   assign  _add_map_x_130_left = ((_net_6469)?data_in341:10'b0)|
    ((_net_2477)?data_in342:10'b0);
   assign  _add_map_x_130_start = start;
   assign  _add_map_x_130_goal = goal;
   assign  _add_map_x_130_now = ((_net_6466)?10'b0100110101:10'b0)|
    ((_net_2474)?10'b0100110110:10'b0);
   assign  _add_map_x_130_add_exe = (_net_6465|_net_2473);
   assign  _add_map_x_130_p_reset = p_reset;
   assign  _add_map_x_130_m_clock = m_clock;
   assign  _add_map_x_129_moto_org_near = ((_net_6464)?data_in_org308:10'b0)|
    ((_net_2472)?data_in_org307:10'b0);
   assign  _add_map_x_129_moto_org_near1 = ((_net_6463)?data_in_org306:10'b0)|
    ((_net_2471)?data_in_org309:10'b0);
   assign  _add_map_x_129_moto_org_near2 = ((_net_6462)?data_in_org275:10'b0)|
    ((_net_2470)?data_in_org276:10'b0);
   assign  _add_map_x_129_moto_org_near3 = ((_net_6461)?data_in_org339:10'b0)|
    ((_net_2469)?data_in_org340:10'b0);
   assign  _add_map_x_129_moto_org = ((_net_6460)?data_in_org307:10'b0)|
    ((_net_2468)?data_in_org308:10'b0);
   assign  _add_map_x_129_sg_up = ((_net_6459)?sg_in308:2'b0)|
    ((_net_2467)?sg_in307:2'b0);
   assign  _add_map_x_129_sg_down = ((_net_6458)?sg_in275:2'b0)|
    ((_net_2466)?sg_in309:2'b0);
   assign  _add_map_x_129_sg_left = ((_net_6456)?sg_in339:2'b0)|
    ((_net_2464)?sg_in340:2'b0);
   assign  _add_map_x_129_sg_right = ((_net_6457)?sg_in306:2'b0)|
    ((_net_2465)?sg_in276:2'b0);
   assign  _add_map_x_129_wall_t_in = dig_w;
   assign  _add_map_x_129_moto = ((_net_6454)?data_in307:10'b0)|
    ((_net_2462)?data_in308:10'b0);
   assign  _add_map_x_129_up = ((_net_6453)?data_in308:10'b0)|
    ((_net_2461)?data_in307:10'b0);
   assign  _add_map_x_129_right = ((_net_6452)?data_in306:10'b0)|
    ((_net_2460)?data_in309:10'b0);
   assign  _add_map_x_129_down = ((_net_6451)?data_in275:10'b0)|
    ((_net_2459)?data_in276:10'b0);
   assign  _add_map_x_129_left = ((_net_6450)?data_in339:10'b0)|
    ((_net_2458)?data_in340:10'b0);
   assign  _add_map_x_129_start = start;
   assign  _add_map_x_129_goal = goal;
   assign  _add_map_x_129_now = ((_net_6447)?10'b0100110011:10'b0)|
    ((_net_2455)?10'b0100110100:10'b0);
   assign  _add_map_x_129_add_exe = (_net_6446|_net_2454);
   assign  _add_map_x_129_p_reset = p_reset;
   assign  _add_map_x_129_m_clock = m_clock;
   assign  _add_map_x_128_moto_org_near = ((_net_6445)?data_in_org306:10'b0)|
    ((_net_2453)?data_in_org305:10'b0);
   assign  _add_map_x_128_moto_org_near1 = ((_net_6444)?data_in_org304:10'b0)|
    ((_net_2452)?data_in_org307:10'b0);
   assign  _add_map_x_128_moto_org_near2 = ((_net_6443)?data_in_org273:10'b0)|
    ((_net_2451)?data_in_org274:10'b0);
   assign  _add_map_x_128_moto_org_near3 = ((_net_6442)?data_in_org337:10'b0)|
    ((_net_2450)?data_in_org338:10'b0);
   assign  _add_map_x_128_moto_org = ((_net_6441)?data_in_org305:10'b0)|
    ((_net_2449)?data_in_org306:10'b0);
   assign  _add_map_x_128_sg_up = ((_net_6440)?sg_in306:2'b0)|
    ((_net_2448)?sg_in305:2'b0);
   assign  _add_map_x_128_sg_down = ((_net_6439)?sg_in273:2'b0)|
    ((_net_2447)?sg_in307:2'b0);
   assign  _add_map_x_128_sg_left = ((_net_6437)?sg_in337:2'b0)|
    ((_net_2445)?sg_in338:2'b0);
   assign  _add_map_x_128_sg_right = ((_net_6438)?sg_in304:2'b0)|
    ((_net_2446)?sg_in274:2'b0);
   assign  _add_map_x_128_wall_t_in = dig_w;
   assign  _add_map_x_128_moto = ((_net_6435)?data_in305:10'b0)|
    ((_net_2443)?data_in306:10'b0);
   assign  _add_map_x_128_up = ((_net_6434)?data_in306:10'b0)|
    ((_net_2442)?data_in305:10'b0);
   assign  _add_map_x_128_right = ((_net_6433)?data_in304:10'b0)|
    ((_net_2441)?data_in307:10'b0);
   assign  _add_map_x_128_down = ((_net_6432)?data_in273:10'b0)|
    ((_net_2440)?data_in274:10'b0);
   assign  _add_map_x_128_left = ((_net_6431)?data_in337:10'b0)|
    ((_net_2439)?data_in338:10'b0);
   assign  _add_map_x_128_start = start;
   assign  _add_map_x_128_goal = goal;
   assign  _add_map_x_128_now = ((_net_6428)?10'b0100110001:10'b0)|
    ((_net_2436)?10'b0100110010:10'b0);
   assign  _add_map_x_128_add_exe = (_net_6427|_net_2435);
   assign  _add_map_x_128_p_reset = p_reset;
   assign  _add_map_x_128_m_clock = m_clock;
   assign  _add_map_x_127_moto_org_near = ((_net_6426)?data_in_org304:10'b0)|
    ((_net_2434)?data_in_org303:10'b0);
   assign  _add_map_x_127_moto_org_near1 = ((_net_6425)?data_in_org302:10'b0)|
    ((_net_2433)?data_in_org305:10'b0);
   assign  _add_map_x_127_moto_org_near2 = ((_net_6424)?data_in_org271:10'b0)|
    ((_net_2432)?data_in_org272:10'b0);
   assign  _add_map_x_127_moto_org_near3 = ((_net_6423)?data_in_org335:10'b0)|
    ((_net_2431)?data_in_org336:10'b0);
   assign  _add_map_x_127_moto_org = ((_net_6422)?data_in_org303:10'b0)|
    ((_net_2430)?data_in_org304:10'b0);
   assign  _add_map_x_127_sg_up = ((_net_6421)?sg_in304:2'b0)|
    ((_net_2429)?sg_in303:2'b0);
   assign  _add_map_x_127_sg_down = ((_net_6420)?sg_in271:2'b0)|
    ((_net_2428)?sg_in305:2'b0);
   assign  _add_map_x_127_sg_left = ((_net_6418)?sg_in335:2'b0)|
    ((_net_2426)?sg_in336:2'b0);
   assign  _add_map_x_127_sg_right = ((_net_6419)?sg_in302:2'b0)|
    ((_net_2427)?sg_in272:2'b0);
   assign  _add_map_x_127_wall_t_in = dig_w;
   assign  _add_map_x_127_moto = ((_net_6416)?data_in303:10'b0)|
    ((_net_2424)?data_in304:10'b0);
   assign  _add_map_x_127_up = ((_net_6415)?data_in304:10'b0)|
    ((_net_2423)?data_in303:10'b0);
   assign  _add_map_x_127_right = ((_net_6414)?data_in302:10'b0)|
    ((_net_2422)?data_in305:10'b0);
   assign  _add_map_x_127_down = ((_net_6413)?data_in271:10'b0)|
    ((_net_2421)?data_in272:10'b0);
   assign  _add_map_x_127_left = ((_net_6412)?data_in335:10'b0)|
    ((_net_2420)?data_in336:10'b0);
   assign  _add_map_x_127_start = start;
   assign  _add_map_x_127_goal = goal;
   assign  _add_map_x_127_now = ((_net_6409)?10'b0100101111:10'b0)|
    ((_net_2417)?10'b0100110000:10'b0);
   assign  _add_map_x_127_add_exe = (_net_6408|_net_2416);
   assign  _add_map_x_127_p_reset = p_reset;
   assign  _add_map_x_127_m_clock = m_clock;
   assign  _add_map_x_126_moto_org_near = ((_net_6407)?data_in_org302:10'b0)|
    ((_net_2415)?data_in_org301:10'b0);
   assign  _add_map_x_126_moto_org_near1 = ((_net_6406)?data_in_org300:10'b0)|
    ((_net_2414)?data_in_org303:10'b0);
   assign  _add_map_x_126_moto_org_near2 = ((_net_6405)?data_in_org269:10'b0)|
    ((_net_2413)?data_in_org270:10'b0);
   assign  _add_map_x_126_moto_org_near3 = ((_net_6404)?data_in_org333:10'b0)|
    ((_net_2412)?data_in_org334:10'b0);
   assign  _add_map_x_126_moto_org = ((_net_6403)?data_in_org301:10'b0)|
    ((_net_2411)?data_in_org302:10'b0);
   assign  _add_map_x_126_sg_up = ((_net_6402)?sg_in302:2'b0)|
    ((_net_2410)?sg_in301:2'b0);
   assign  _add_map_x_126_sg_down = ((_net_6401)?sg_in269:2'b0)|
    ((_net_2409)?sg_in303:2'b0);
   assign  _add_map_x_126_sg_left = ((_net_6399)?sg_in333:2'b0)|
    ((_net_2407)?sg_in334:2'b0);
   assign  _add_map_x_126_sg_right = ((_net_6400)?sg_in300:2'b0)|
    ((_net_2408)?sg_in270:2'b0);
   assign  _add_map_x_126_wall_t_in = dig_w;
   assign  _add_map_x_126_moto = ((_net_6397)?data_in301:10'b0)|
    ((_net_2405)?data_in302:10'b0);
   assign  _add_map_x_126_up = ((_net_6396)?data_in302:10'b0)|
    ((_net_2404)?data_in301:10'b0);
   assign  _add_map_x_126_right = ((_net_6395)?data_in300:10'b0)|
    ((_net_2403)?data_in303:10'b0);
   assign  _add_map_x_126_down = ((_net_6394)?data_in269:10'b0)|
    ((_net_2402)?data_in270:10'b0);
   assign  _add_map_x_126_left = ((_net_6393)?data_in333:10'b0)|
    ((_net_2401)?data_in334:10'b0);
   assign  _add_map_x_126_start = start;
   assign  _add_map_x_126_goal = goal;
   assign  _add_map_x_126_now = ((_net_6390)?10'b0100101101:10'b0)|
    ((_net_2398)?10'b0100101110:10'b0);
   assign  _add_map_x_126_add_exe = (_net_6389|_net_2397);
   assign  _add_map_x_126_p_reset = p_reset;
   assign  _add_map_x_126_m_clock = m_clock;
   assign  _add_map_x_125_moto_org_near = ((_net_6388)?data_in_org300:10'b0)|
    ((_net_2396)?data_in_org299:10'b0);
   assign  _add_map_x_125_moto_org_near1 = ((_net_6387)?data_in_org298:10'b0)|
    ((_net_2395)?data_in_org301:10'b0);
   assign  _add_map_x_125_moto_org_near2 = ((_net_6386)?data_in_org267:10'b0)|
    ((_net_2394)?data_in_org268:10'b0);
   assign  _add_map_x_125_moto_org_near3 = ((_net_6385)?data_in_org331:10'b0)|
    ((_net_2393)?data_in_org332:10'b0);
   assign  _add_map_x_125_moto_org = ((_net_6384)?data_in_org299:10'b0)|
    ((_net_2392)?data_in_org300:10'b0);
   assign  _add_map_x_125_sg_up = ((_net_6383)?sg_in300:2'b0)|
    ((_net_2391)?sg_in299:2'b0);
   assign  _add_map_x_125_sg_down = ((_net_6382)?sg_in267:2'b0)|
    ((_net_2390)?sg_in301:2'b0);
   assign  _add_map_x_125_sg_left = ((_net_6380)?sg_in331:2'b0)|
    ((_net_2388)?sg_in332:2'b0);
   assign  _add_map_x_125_sg_right = ((_net_6381)?sg_in298:2'b0)|
    ((_net_2389)?sg_in268:2'b0);
   assign  _add_map_x_125_wall_t_in = dig_w;
   assign  _add_map_x_125_moto = ((_net_6378)?data_in299:10'b0)|
    ((_net_2386)?data_in300:10'b0);
   assign  _add_map_x_125_up = ((_net_6377)?data_in300:10'b0)|
    ((_net_2385)?data_in299:10'b0);
   assign  _add_map_x_125_right = ((_net_6376)?data_in298:10'b0)|
    ((_net_2384)?data_in301:10'b0);
   assign  _add_map_x_125_down = ((_net_6375)?data_in267:10'b0)|
    ((_net_2383)?data_in268:10'b0);
   assign  _add_map_x_125_left = ((_net_6374)?data_in331:10'b0)|
    ((_net_2382)?data_in332:10'b0);
   assign  _add_map_x_125_start = start;
   assign  _add_map_x_125_goal = goal;
   assign  _add_map_x_125_now = ((_net_6371)?10'b0100101011:10'b0)|
    ((_net_2379)?10'b0100101100:10'b0);
   assign  _add_map_x_125_add_exe = (_net_6370|_net_2378);
   assign  _add_map_x_125_p_reset = p_reset;
   assign  _add_map_x_125_m_clock = m_clock;
   assign  _add_map_x_124_moto_org_near = ((_net_6369)?data_in_org298:10'b0)|
    ((_net_2377)?data_in_org297:10'b0);
   assign  _add_map_x_124_moto_org_near1 = ((_net_6368)?data_in_org296:10'b0)|
    ((_net_2376)?data_in_org299:10'b0);
   assign  _add_map_x_124_moto_org_near2 = ((_net_6367)?data_in_org265:10'b0)|
    ((_net_2375)?data_in_org266:10'b0);
   assign  _add_map_x_124_moto_org_near3 = ((_net_6366)?data_in_org329:10'b0)|
    ((_net_2374)?data_in_org330:10'b0);
   assign  _add_map_x_124_moto_org = ((_net_6365)?data_in_org297:10'b0)|
    ((_net_2373)?data_in_org298:10'b0);
   assign  _add_map_x_124_sg_up = ((_net_6364)?sg_in298:2'b0)|
    ((_net_2372)?sg_in297:2'b0);
   assign  _add_map_x_124_sg_down = ((_net_6363)?sg_in265:2'b0)|
    ((_net_2371)?sg_in299:2'b0);
   assign  _add_map_x_124_sg_left = ((_net_6361)?sg_in329:2'b0)|
    ((_net_2369)?sg_in330:2'b0);
   assign  _add_map_x_124_sg_right = ((_net_6362)?sg_in296:2'b0)|
    ((_net_2370)?sg_in266:2'b0);
   assign  _add_map_x_124_wall_t_in = dig_w;
   assign  _add_map_x_124_moto = ((_net_6359)?data_in297:10'b0)|
    ((_net_2367)?data_in298:10'b0);
   assign  _add_map_x_124_up = ((_net_6358)?data_in298:10'b0)|
    ((_net_2366)?data_in297:10'b0);
   assign  _add_map_x_124_right = ((_net_6357)?data_in296:10'b0)|
    ((_net_2365)?data_in299:10'b0);
   assign  _add_map_x_124_down = ((_net_6356)?data_in265:10'b0)|
    ((_net_2364)?data_in266:10'b0);
   assign  _add_map_x_124_left = ((_net_6355)?data_in329:10'b0)|
    ((_net_2363)?data_in330:10'b0);
   assign  _add_map_x_124_start = start;
   assign  _add_map_x_124_goal = goal;
   assign  _add_map_x_124_now = ((_net_6352)?10'b0100101001:10'b0)|
    ((_net_2360)?10'b0100101010:10'b0);
   assign  _add_map_x_124_add_exe = (_net_6351|_net_2359);
   assign  _add_map_x_124_p_reset = p_reset;
   assign  _add_map_x_124_m_clock = m_clock;
   assign  _add_map_x_123_moto_org_near = ((_net_6350)?data_in_org296:10'b0)|
    ((_net_2358)?data_in_org295:10'b0);
   assign  _add_map_x_123_moto_org_near1 = ((_net_6349)?data_in_org294:10'b0)|
    ((_net_2357)?data_in_org297:10'b0);
   assign  _add_map_x_123_moto_org_near2 = ((_net_6348)?data_in_org263:10'b0)|
    ((_net_2356)?data_in_org264:10'b0);
   assign  _add_map_x_123_moto_org_near3 = ((_net_6347)?data_in_org327:10'b0)|
    ((_net_2355)?data_in_org328:10'b0);
   assign  _add_map_x_123_moto_org = ((_net_6346)?data_in_org295:10'b0)|
    ((_net_2354)?data_in_org296:10'b0);
   assign  _add_map_x_123_sg_up = ((_net_6345)?sg_in296:2'b0)|
    ((_net_2353)?sg_in295:2'b0);
   assign  _add_map_x_123_sg_down = ((_net_6344)?sg_in263:2'b0)|
    ((_net_2352)?sg_in297:2'b0);
   assign  _add_map_x_123_sg_left = ((_net_6342)?sg_in327:2'b0)|
    ((_net_2350)?sg_in328:2'b0);
   assign  _add_map_x_123_sg_right = ((_net_6343)?sg_in294:2'b0)|
    ((_net_2351)?sg_in264:2'b0);
   assign  _add_map_x_123_wall_t_in = dig_w;
   assign  _add_map_x_123_moto = ((_net_6340)?data_in295:10'b0)|
    ((_net_2348)?data_in296:10'b0);
   assign  _add_map_x_123_up = ((_net_6339)?data_in296:10'b0)|
    ((_net_2347)?data_in295:10'b0);
   assign  _add_map_x_123_right = ((_net_6338)?data_in294:10'b0)|
    ((_net_2346)?data_in297:10'b0);
   assign  _add_map_x_123_down = ((_net_6337)?data_in263:10'b0)|
    ((_net_2345)?data_in264:10'b0);
   assign  _add_map_x_123_left = ((_net_6336)?data_in327:10'b0)|
    ((_net_2344)?data_in328:10'b0);
   assign  _add_map_x_123_start = start;
   assign  _add_map_x_123_goal = goal;
   assign  _add_map_x_123_now = ((_net_6333)?10'b0100100111:10'b0)|
    ((_net_2341)?10'b0100101000:10'b0);
   assign  _add_map_x_123_add_exe = (_net_6332|_net_2340);
   assign  _add_map_x_123_p_reset = p_reset;
   assign  _add_map_x_123_m_clock = m_clock;
   assign  _add_map_x_122_moto_org_near = ((_net_6331)?data_in_org294:10'b0)|
    ((_net_2339)?data_in_org293:10'b0);
   assign  _add_map_x_122_moto_org_near1 = ((_net_6330)?data_in_org292:10'b0)|
    ((_net_2338)?data_in_org295:10'b0);
   assign  _add_map_x_122_moto_org_near2 = ((_net_6329)?data_in_org261:10'b0)|
    ((_net_2337)?data_in_org262:10'b0);
   assign  _add_map_x_122_moto_org_near3 = ((_net_6328)?data_in_org325:10'b0)|
    ((_net_2336)?data_in_org326:10'b0);
   assign  _add_map_x_122_moto_org = ((_net_6327)?data_in_org293:10'b0)|
    ((_net_2335)?data_in_org294:10'b0);
   assign  _add_map_x_122_sg_up = ((_net_6326)?sg_in294:2'b0)|
    ((_net_2334)?sg_in293:2'b0);
   assign  _add_map_x_122_sg_down = ((_net_6325)?sg_in261:2'b0)|
    ((_net_2333)?sg_in295:2'b0);
   assign  _add_map_x_122_sg_left = ((_net_6323)?sg_in325:2'b0)|
    ((_net_2331)?sg_in326:2'b0);
   assign  _add_map_x_122_sg_right = ((_net_6324)?sg_in292:2'b0)|
    ((_net_2332)?sg_in262:2'b0);
   assign  _add_map_x_122_wall_t_in = dig_w;
   assign  _add_map_x_122_moto = ((_net_6321)?data_in293:10'b0)|
    ((_net_2329)?data_in294:10'b0);
   assign  _add_map_x_122_up = ((_net_6320)?data_in294:10'b0)|
    ((_net_2328)?data_in293:10'b0);
   assign  _add_map_x_122_right = ((_net_6319)?data_in292:10'b0)|
    ((_net_2327)?data_in295:10'b0);
   assign  _add_map_x_122_down = ((_net_6318)?data_in261:10'b0)|
    ((_net_2326)?data_in262:10'b0);
   assign  _add_map_x_122_left = ((_net_6317)?data_in325:10'b0)|
    ((_net_2325)?data_in326:10'b0);
   assign  _add_map_x_122_start = start;
   assign  _add_map_x_122_goal = goal;
   assign  _add_map_x_122_now = ((_net_6314)?10'b0100100101:10'b0)|
    ((_net_2322)?10'b0100100110:10'b0);
   assign  _add_map_x_122_add_exe = (_net_6313|_net_2321);
   assign  _add_map_x_122_p_reset = p_reset;
   assign  _add_map_x_122_m_clock = m_clock;
   assign  _add_map_x_121_moto_org_near = ((_net_6312)?data_in_org292:10'b0)|
    ((_net_2320)?data_in_org291:10'b0);
   assign  _add_map_x_121_moto_org_near1 = ((_net_6311)?data_in_org290:10'b0)|
    ((_net_2319)?data_in_org293:10'b0);
   assign  _add_map_x_121_moto_org_near2 = ((_net_6310)?data_in_org259:10'b0)|
    ((_net_2318)?data_in_org260:10'b0);
   assign  _add_map_x_121_moto_org_near3 = ((_net_6309)?data_in_org323:10'b0)|
    ((_net_2317)?data_in_org324:10'b0);
   assign  _add_map_x_121_moto_org = ((_net_6308)?data_in_org291:10'b0)|
    ((_net_2316)?data_in_org292:10'b0);
   assign  _add_map_x_121_sg_up = ((_net_6307)?sg_in292:2'b0)|
    ((_net_2315)?sg_in291:2'b0);
   assign  _add_map_x_121_sg_down = ((_net_6306)?sg_in259:2'b0)|
    ((_net_2314)?sg_in293:2'b0);
   assign  _add_map_x_121_sg_left = ((_net_6304)?sg_in323:2'b0)|
    ((_net_2312)?sg_in324:2'b0);
   assign  _add_map_x_121_sg_right = ((_net_6305)?sg_in290:2'b0)|
    ((_net_2313)?sg_in260:2'b0);
   assign  _add_map_x_121_wall_t_in = dig_w;
   assign  _add_map_x_121_moto = ((_net_6302)?data_in291:10'b0)|
    ((_net_2310)?data_in292:10'b0);
   assign  _add_map_x_121_up = ((_net_6301)?data_in292:10'b0)|
    ((_net_2309)?data_in291:10'b0);
   assign  _add_map_x_121_right = ((_net_6300)?data_in290:10'b0)|
    ((_net_2308)?data_in293:10'b0);
   assign  _add_map_x_121_down = ((_net_6299)?data_in259:10'b0)|
    ((_net_2307)?data_in260:10'b0);
   assign  _add_map_x_121_left = ((_net_6298)?data_in323:10'b0)|
    ((_net_2306)?data_in324:10'b0);
   assign  _add_map_x_121_start = start;
   assign  _add_map_x_121_goal = goal;
   assign  _add_map_x_121_now = ((_net_6295)?10'b0100100011:10'b0)|
    ((_net_2303)?10'b0100100100:10'b0);
   assign  _add_map_x_121_add_exe = (_net_6294|_net_2302);
   assign  _add_map_x_121_p_reset = p_reset;
   assign  _add_map_x_121_m_clock = m_clock;
   assign  _add_map_x_120_moto_org_near = ((_net_6293)?data_in_org290:10'b0)|
    ((_net_2301)?data_in_org289:10'b0);
   assign  _add_map_x_120_moto_org_near1 = ((_net_6292)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2300)?data_in_org291:10'b0);
   assign  _add_map_x_120_moto_org_near2 = ((_net_6291)?data_in_org257:10'b0)|
    ((_net_2299)?data_in_org258:10'b0);
   assign  _add_map_x_120_moto_org_near3 = ((_net_6290)?data_in_org321:10'b0)|
    ((_net_2298)?data_in_org322:10'b0);
   assign  _add_map_x_120_moto_org = ((_net_6289)?data_in_org289:10'b0)|
    ((_net_2297)?data_in_org290:10'b0);
   assign  _add_map_x_120_sg_up = ((_net_6288)?sg_in290:2'b0)|
    ((_net_2296)?sg_in289:2'b0);
   assign  _add_map_x_120_sg_down = ((_net_6287)?sg_in257:2'b0)|
    ((_net_2295)?sg_in291:2'b0);
   assign  _add_map_x_120_sg_left = ((_net_6285)?sg_in321:2'b0)|
    ((_net_2293)?sg_in322:2'b0);
   assign  _add_map_x_120_sg_right = ((_net_6286)?3'b000:2'b0)|
    ((_net_2294)?sg_in258:2'b0);
   assign  _add_map_x_120_wall_t_in = dig_w;
   assign  _add_map_x_120_moto = ((_net_6283)?data_in289:10'b0)|
    ((_net_2291)?data_in290:10'b0);
   assign  _add_map_x_120_up = ((_net_6282)?data_in290:10'b0)|
    ((_net_2290)?data_in289:10'b0);
   assign  _add_map_x_120_right = ((_net_6281)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2289)?data_in291:10'b0);
   assign  _add_map_x_120_down = ((_net_6280)?data_in257:10'b0)|
    ((_net_2288)?data_in258:10'b0);
   assign  _add_map_x_120_left = ((_net_6279)?data_in321:10'b0)|
    ((_net_2287)?data_in322:10'b0);
   assign  _add_map_x_120_start = start;
   assign  _add_map_x_120_goal = goal;
   assign  _add_map_x_120_now = ((_net_6276)?10'b0100100001:10'b0)|
    ((_net_2284)?10'b0100100010:10'b0);
   assign  _add_map_x_120_add_exe = (_net_6275|_net_2283);
   assign  _add_map_x_120_p_reset = p_reset;
   assign  _add_map_x_120_m_clock = m_clock;
   assign  _add_map_x_119_moto_org_near = ((_net_6274)?data_in_org285:10'b0)|
    ((_net_2282)?data_in_org286:10'b0);
   assign  _add_map_x_119_moto_org_near1 = ((_net_6273)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2281)?data_in_org284:10'b0);
   assign  _add_map_x_119_moto_org_near2 = ((_net_6272)?data_in_org254:10'b0)|
    ((_net_2280)?data_in_org253:10'b0);
   assign  _add_map_x_119_moto_org_near3 = ((_net_6271)?data_in_org318:10'b0)|
    ((_net_2279)?data_in_org317:10'b0);
   assign  _add_map_x_119_moto_org = ((_net_6270)?data_in_org286:10'b0)|
    ((_net_2278)?data_in_org285:10'b0);
   assign  _add_map_x_119_sg_up = ((_net_6269)?sg_in285:2'b0)|
    ((_net_2277)?sg_in286:2'b0);
   assign  _add_map_x_119_sg_down = ((_net_6268)?3'b000:2'b0)|
    ((_net_2276)?sg_in284:2'b0);
   assign  _add_map_x_119_sg_left = ((_net_6266)?sg_in318:2'b0)|
    ((_net_2274)?sg_in317:2'b0);
   assign  _add_map_x_119_sg_right = ((_net_6267)?sg_in254:2'b0)|
    ((_net_2275)?sg_in253:2'b0);
   assign  _add_map_x_119_wall_t_in = dig_w;
   assign  _add_map_x_119_moto = ((_net_6264)?data_in286:10'b0)|
    ((_net_2272)?data_in285:10'b0);
   assign  _add_map_x_119_up = ((_net_6263)?data_in285:10'b0)|
    ((_net_2271)?data_in286:10'b0);
   assign  _add_map_x_119_right = ((_net_6262)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_2270)?data_in284:10'b0);
   assign  _add_map_x_119_down = ((_net_6261)?data_in254:10'b0)|
    ((_net_2269)?data_in253:10'b0);
   assign  _add_map_x_119_left = ((_net_6260)?data_in318:10'b0)|
    ((_net_2268)?data_in317:10'b0);
   assign  _add_map_x_119_start = start;
   assign  _add_map_x_119_goal = goal;
   assign  _add_map_x_119_now = ((_net_6257)?10'b0100011110:10'b0)|
    ((_net_2265)?10'b0100011101:10'b0);
   assign  _add_map_x_119_add_exe = (_net_6256|_net_2264);
   assign  _add_map_x_119_p_reset = p_reset;
   assign  _add_map_x_119_m_clock = m_clock;
   assign  _add_map_x_118_moto_org_near = ((_net_6255)?data_in_org283:10'b0)|
    ((_net_2263)?data_in_org284:10'b0);
   assign  _add_map_x_118_moto_org_near1 = ((_net_6254)?data_in_org285:10'b0)|
    ((_net_2262)?data_in_org282:10'b0);
   assign  _add_map_x_118_moto_org_near2 = ((_net_6253)?data_in_org252:10'b0)|
    ((_net_2261)?data_in_org251:10'b0);
   assign  _add_map_x_118_moto_org_near3 = ((_net_6252)?data_in_org316:10'b0)|
    ((_net_2260)?data_in_org315:10'b0);
   assign  _add_map_x_118_moto_org = ((_net_6251)?data_in_org284:10'b0)|
    ((_net_2259)?data_in_org283:10'b0);
   assign  _add_map_x_118_sg_up = ((_net_6250)?sg_in283:2'b0)|
    ((_net_2258)?sg_in284:2'b0);
   assign  _add_map_x_118_sg_down = ((_net_6249)?sg_in285:2'b0)|
    ((_net_2257)?sg_in282:2'b0);
   assign  _add_map_x_118_sg_left = ((_net_6247)?sg_in316:2'b0)|
    ((_net_2255)?sg_in315:2'b0);
   assign  _add_map_x_118_sg_right = ((_net_6248)?sg_in252:2'b0)|
    ((_net_2256)?sg_in251:2'b0);
   assign  _add_map_x_118_wall_t_in = dig_w;
   assign  _add_map_x_118_moto = ((_net_6245)?data_in284:10'b0)|
    ((_net_2253)?data_in283:10'b0);
   assign  _add_map_x_118_up = ((_net_6244)?data_in283:10'b0)|
    ((_net_2252)?data_in284:10'b0);
   assign  _add_map_x_118_right = ((_net_6243)?data_in285:10'b0)|
    ((_net_2251)?data_in282:10'b0);
   assign  _add_map_x_118_down = ((_net_6242)?data_in252:10'b0)|
    ((_net_2250)?data_in251:10'b0);
   assign  _add_map_x_118_left = ((_net_6241)?data_in316:10'b0)|
    ((_net_2249)?data_in315:10'b0);
   assign  _add_map_x_118_start = start;
   assign  _add_map_x_118_goal = goal;
   assign  _add_map_x_118_now = ((_net_6238)?10'b0100011100:10'b0)|
    ((_net_2246)?10'b0100011011:10'b0);
   assign  _add_map_x_118_add_exe = (_net_6237|_net_2245);
   assign  _add_map_x_118_p_reset = p_reset;
   assign  _add_map_x_118_m_clock = m_clock;
   assign  _add_map_x_117_moto_org_near = ((_net_6236)?data_in_org281:10'b0)|
    ((_net_2244)?data_in_org282:10'b0);
   assign  _add_map_x_117_moto_org_near1 = ((_net_6235)?data_in_org283:10'b0)|
    ((_net_2243)?data_in_org280:10'b0);
   assign  _add_map_x_117_moto_org_near2 = ((_net_6234)?data_in_org250:10'b0)|
    ((_net_2242)?data_in_org249:10'b0);
   assign  _add_map_x_117_moto_org_near3 = ((_net_6233)?data_in_org314:10'b0)|
    ((_net_2241)?data_in_org313:10'b0);
   assign  _add_map_x_117_moto_org = ((_net_6232)?data_in_org282:10'b0)|
    ((_net_2240)?data_in_org281:10'b0);
   assign  _add_map_x_117_sg_up = ((_net_6231)?sg_in281:2'b0)|
    ((_net_2239)?sg_in282:2'b0);
   assign  _add_map_x_117_sg_down = ((_net_6230)?sg_in283:2'b0)|
    ((_net_2238)?sg_in280:2'b0);
   assign  _add_map_x_117_sg_left = ((_net_6228)?sg_in314:2'b0)|
    ((_net_2236)?sg_in313:2'b0);
   assign  _add_map_x_117_sg_right = ((_net_6229)?sg_in250:2'b0)|
    ((_net_2237)?sg_in249:2'b0);
   assign  _add_map_x_117_wall_t_in = dig_w;
   assign  _add_map_x_117_moto = ((_net_6226)?data_in282:10'b0)|
    ((_net_2234)?data_in281:10'b0);
   assign  _add_map_x_117_up = ((_net_6225)?data_in281:10'b0)|
    ((_net_2233)?data_in282:10'b0);
   assign  _add_map_x_117_right = ((_net_6224)?data_in283:10'b0)|
    ((_net_2232)?data_in280:10'b0);
   assign  _add_map_x_117_down = ((_net_6223)?data_in250:10'b0)|
    ((_net_2231)?data_in249:10'b0);
   assign  _add_map_x_117_left = ((_net_6222)?data_in314:10'b0)|
    ((_net_2230)?data_in313:10'b0);
   assign  _add_map_x_117_start = start;
   assign  _add_map_x_117_goal = goal;
   assign  _add_map_x_117_now = ((_net_6219)?10'b0100011010:10'b0)|
    ((_net_2227)?10'b0100011001:10'b0);
   assign  _add_map_x_117_add_exe = (_net_6218|_net_2226);
   assign  _add_map_x_117_p_reset = p_reset;
   assign  _add_map_x_117_m_clock = m_clock;
   assign  _add_map_x_116_moto_org_near = ((_net_6217)?data_in_org279:10'b0)|
    ((_net_2225)?data_in_org280:10'b0);
   assign  _add_map_x_116_moto_org_near1 = ((_net_6216)?data_in_org281:10'b0)|
    ((_net_2224)?data_in_org278:10'b0);
   assign  _add_map_x_116_moto_org_near2 = ((_net_6215)?data_in_org248:10'b0)|
    ((_net_2223)?data_in_org247:10'b0);
   assign  _add_map_x_116_moto_org_near3 = ((_net_6214)?data_in_org312:10'b0)|
    ((_net_2222)?data_in_org311:10'b0);
   assign  _add_map_x_116_moto_org = ((_net_6213)?data_in_org280:10'b0)|
    ((_net_2221)?data_in_org279:10'b0);
   assign  _add_map_x_116_sg_up = ((_net_6212)?sg_in279:2'b0)|
    ((_net_2220)?sg_in280:2'b0);
   assign  _add_map_x_116_sg_down = ((_net_6211)?sg_in281:2'b0)|
    ((_net_2219)?sg_in278:2'b0);
   assign  _add_map_x_116_sg_left = ((_net_6209)?sg_in312:2'b0)|
    ((_net_2217)?sg_in311:2'b0);
   assign  _add_map_x_116_sg_right = ((_net_6210)?sg_in248:2'b0)|
    ((_net_2218)?sg_in247:2'b0);
   assign  _add_map_x_116_wall_t_in = dig_w;
   assign  _add_map_x_116_moto = ((_net_6207)?data_in280:10'b0)|
    ((_net_2215)?data_in279:10'b0);
   assign  _add_map_x_116_up = ((_net_6206)?data_in279:10'b0)|
    ((_net_2214)?data_in280:10'b0);
   assign  _add_map_x_116_right = ((_net_6205)?data_in281:10'b0)|
    ((_net_2213)?data_in278:10'b0);
   assign  _add_map_x_116_down = ((_net_6204)?data_in248:10'b0)|
    ((_net_2212)?data_in247:10'b0);
   assign  _add_map_x_116_left = ((_net_6203)?data_in312:10'b0)|
    ((_net_2211)?data_in311:10'b0);
   assign  _add_map_x_116_start = start;
   assign  _add_map_x_116_goal = goal;
   assign  _add_map_x_116_now = ((_net_6200)?10'b0100011000:10'b0)|
    ((_net_2208)?10'b0100010111:10'b0);
   assign  _add_map_x_116_add_exe = (_net_6199|_net_2207);
   assign  _add_map_x_116_p_reset = p_reset;
   assign  _add_map_x_116_m_clock = m_clock;
   assign  _add_map_x_115_moto_org_near = ((_net_6198)?data_in_org277:10'b0)|
    ((_net_2206)?data_in_org278:10'b0);
   assign  _add_map_x_115_moto_org_near1 = ((_net_6197)?data_in_org279:10'b0)|
    ((_net_2205)?data_in_org276:10'b0);
   assign  _add_map_x_115_moto_org_near2 = ((_net_6196)?data_in_org246:10'b0)|
    ((_net_2204)?data_in_org245:10'b0);
   assign  _add_map_x_115_moto_org_near3 = ((_net_6195)?data_in_org310:10'b0)|
    ((_net_2203)?data_in_org309:10'b0);
   assign  _add_map_x_115_moto_org = ((_net_6194)?data_in_org278:10'b0)|
    ((_net_2202)?data_in_org277:10'b0);
   assign  _add_map_x_115_sg_up = ((_net_6193)?sg_in277:2'b0)|
    ((_net_2201)?sg_in278:2'b0);
   assign  _add_map_x_115_sg_down = ((_net_6192)?sg_in279:2'b0)|
    ((_net_2200)?sg_in276:2'b0);
   assign  _add_map_x_115_sg_left = ((_net_6190)?sg_in310:2'b0)|
    ((_net_2198)?sg_in309:2'b0);
   assign  _add_map_x_115_sg_right = ((_net_6191)?sg_in246:2'b0)|
    ((_net_2199)?sg_in245:2'b0);
   assign  _add_map_x_115_wall_t_in = dig_w;
   assign  _add_map_x_115_moto = ((_net_6188)?data_in278:10'b0)|
    ((_net_2196)?data_in277:10'b0);
   assign  _add_map_x_115_up = ((_net_6187)?data_in277:10'b0)|
    ((_net_2195)?data_in278:10'b0);
   assign  _add_map_x_115_right = ((_net_6186)?data_in279:10'b0)|
    ((_net_2194)?data_in276:10'b0);
   assign  _add_map_x_115_down = ((_net_6185)?data_in246:10'b0)|
    ((_net_2193)?data_in245:10'b0);
   assign  _add_map_x_115_left = ((_net_6184)?data_in310:10'b0)|
    ((_net_2192)?data_in309:10'b0);
   assign  _add_map_x_115_start = start;
   assign  _add_map_x_115_goal = goal;
   assign  _add_map_x_115_now = ((_net_6181)?10'b0100010110:10'b0)|
    ((_net_2189)?10'b0100010101:10'b0);
   assign  _add_map_x_115_add_exe = (_net_6180|_net_2188);
   assign  _add_map_x_115_p_reset = p_reset;
   assign  _add_map_x_115_m_clock = m_clock;
   assign  _add_map_x_114_moto_org_near = ((_net_6179)?data_in_org275:10'b0)|
    ((_net_2187)?data_in_org276:10'b0);
   assign  _add_map_x_114_moto_org_near1 = ((_net_6178)?data_in_org277:10'b0)|
    ((_net_2186)?data_in_org274:10'b0);
   assign  _add_map_x_114_moto_org_near2 = ((_net_6177)?data_in_org244:10'b0)|
    ((_net_2185)?data_in_org243:10'b0);
   assign  _add_map_x_114_moto_org_near3 = ((_net_6176)?data_in_org308:10'b0)|
    ((_net_2184)?data_in_org307:10'b0);
   assign  _add_map_x_114_moto_org = ((_net_6175)?data_in_org276:10'b0)|
    ((_net_2183)?data_in_org275:10'b0);
   assign  _add_map_x_114_sg_up = ((_net_6174)?sg_in275:2'b0)|
    ((_net_2182)?sg_in276:2'b0);
   assign  _add_map_x_114_sg_down = ((_net_6173)?sg_in277:2'b0)|
    ((_net_2181)?sg_in274:2'b0);
   assign  _add_map_x_114_sg_left = ((_net_6171)?sg_in308:2'b0)|
    ((_net_2179)?sg_in307:2'b0);
   assign  _add_map_x_114_sg_right = ((_net_6172)?sg_in244:2'b0)|
    ((_net_2180)?sg_in243:2'b0);
   assign  _add_map_x_114_wall_t_in = dig_w;
   assign  _add_map_x_114_moto = ((_net_6169)?data_in276:10'b0)|
    ((_net_2177)?data_in275:10'b0);
   assign  _add_map_x_114_up = ((_net_6168)?data_in275:10'b0)|
    ((_net_2176)?data_in276:10'b0);
   assign  _add_map_x_114_right = ((_net_6167)?data_in277:10'b0)|
    ((_net_2175)?data_in274:10'b0);
   assign  _add_map_x_114_down = ((_net_6166)?data_in244:10'b0)|
    ((_net_2174)?data_in243:10'b0);
   assign  _add_map_x_114_left = ((_net_6165)?data_in308:10'b0)|
    ((_net_2173)?data_in307:10'b0);
   assign  _add_map_x_114_start = start;
   assign  _add_map_x_114_goal = goal;
   assign  _add_map_x_114_now = ((_net_6162)?10'b0100010100:10'b0)|
    ((_net_2170)?10'b0100010011:10'b0);
   assign  _add_map_x_114_add_exe = (_net_6161|_net_2169);
   assign  _add_map_x_114_p_reset = p_reset;
   assign  _add_map_x_114_m_clock = m_clock;
   assign  _add_map_x_113_moto_org_near = ((_net_6160)?data_in_org273:10'b0)|
    ((_net_2168)?data_in_org274:10'b0);
   assign  _add_map_x_113_moto_org_near1 = ((_net_6159)?data_in_org275:10'b0)|
    ((_net_2167)?data_in_org272:10'b0);
   assign  _add_map_x_113_moto_org_near2 = ((_net_6158)?data_in_org242:10'b0)|
    ((_net_2166)?data_in_org241:10'b0);
   assign  _add_map_x_113_moto_org_near3 = ((_net_6157)?data_in_org306:10'b0)|
    ((_net_2165)?data_in_org305:10'b0);
   assign  _add_map_x_113_moto_org = ((_net_6156)?data_in_org274:10'b0)|
    ((_net_2164)?data_in_org273:10'b0);
   assign  _add_map_x_113_sg_up = ((_net_6155)?sg_in273:2'b0)|
    ((_net_2163)?sg_in274:2'b0);
   assign  _add_map_x_113_sg_down = ((_net_6154)?sg_in275:2'b0)|
    ((_net_2162)?sg_in272:2'b0);
   assign  _add_map_x_113_sg_left = ((_net_6152)?sg_in306:2'b0)|
    ((_net_2160)?sg_in305:2'b0);
   assign  _add_map_x_113_sg_right = ((_net_6153)?sg_in242:2'b0)|
    ((_net_2161)?sg_in241:2'b0);
   assign  _add_map_x_113_wall_t_in = dig_w;
   assign  _add_map_x_113_moto = ((_net_6150)?data_in274:10'b0)|
    ((_net_2158)?data_in273:10'b0);
   assign  _add_map_x_113_up = ((_net_6149)?data_in273:10'b0)|
    ((_net_2157)?data_in274:10'b0);
   assign  _add_map_x_113_right = ((_net_6148)?data_in275:10'b0)|
    ((_net_2156)?data_in272:10'b0);
   assign  _add_map_x_113_down = ((_net_6147)?data_in242:10'b0)|
    ((_net_2155)?data_in241:10'b0);
   assign  _add_map_x_113_left = ((_net_6146)?data_in306:10'b0)|
    ((_net_2154)?data_in305:10'b0);
   assign  _add_map_x_113_start = start;
   assign  _add_map_x_113_goal = goal;
   assign  _add_map_x_113_now = ((_net_6143)?10'b0100010010:10'b0)|
    ((_net_2151)?10'b0100010001:10'b0);
   assign  _add_map_x_113_add_exe = (_net_6142|_net_2150);
   assign  _add_map_x_113_p_reset = p_reset;
   assign  _add_map_x_113_m_clock = m_clock;
   assign  _add_map_x_112_moto_org_near = ((_net_6141)?data_in_org271:10'b0)|
    ((_net_2149)?data_in_org272:10'b0);
   assign  _add_map_x_112_moto_org_near1 = ((_net_6140)?data_in_org273:10'b0)|
    ((_net_2148)?data_in_org270:10'b0);
   assign  _add_map_x_112_moto_org_near2 = ((_net_6139)?data_in_org240:10'b0)|
    ((_net_2147)?data_in_org239:10'b0);
   assign  _add_map_x_112_moto_org_near3 = ((_net_6138)?data_in_org304:10'b0)|
    ((_net_2146)?data_in_org303:10'b0);
   assign  _add_map_x_112_moto_org = ((_net_6137)?data_in_org272:10'b0)|
    ((_net_2145)?data_in_org271:10'b0);
   assign  _add_map_x_112_sg_up = ((_net_6136)?sg_in271:2'b0)|
    ((_net_2144)?sg_in272:2'b0);
   assign  _add_map_x_112_sg_down = ((_net_6135)?sg_in273:2'b0)|
    ((_net_2143)?sg_in270:2'b0);
   assign  _add_map_x_112_sg_left = ((_net_6133)?sg_in304:2'b0)|
    ((_net_2141)?sg_in303:2'b0);
   assign  _add_map_x_112_sg_right = ((_net_6134)?sg_in240:2'b0)|
    ((_net_2142)?sg_in239:2'b0);
   assign  _add_map_x_112_wall_t_in = dig_w;
   assign  _add_map_x_112_moto = ((_net_6131)?data_in272:10'b0)|
    ((_net_2139)?data_in271:10'b0);
   assign  _add_map_x_112_up = ((_net_6130)?data_in271:10'b0)|
    ((_net_2138)?data_in272:10'b0);
   assign  _add_map_x_112_right = ((_net_6129)?data_in273:10'b0)|
    ((_net_2137)?data_in270:10'b0);
   assign  _add_map_x_112_down = ((_net_6128)?data_in240:10'b0)|
    ((_net_2136)?data_in239:10'b0);
   assign  _add_map_x_112_left = ((_net_6127)?data_in304:10'b0)|
    ((_net_2135)?data_in303:10'b0);
   assign  _add_map_x_112_start = start;
   assign  _add_map_x_112_goal = goal;
   assign  _add_map_x_112_now = ((_net_6124)?10'b0100010000:10'b0)|
    ((_net_2132)?10'b0100001111:10'b0);
   assign  _add_map_x_112_add_exe = (_net_6123|_net_2131);
   assign  _add_map_x_112_p_reset = p_reset;
   assign  _add_map_x_112_m_clock = m_clock;
   assign  _add_map_x_111_moto_org_near = ((_net_6122)?data_in_org269:10'b0)|
    ((_net_2130)?data_in_org270:10'b0);
   assign  _add_map_x_111_moto_org_near1 = ((_net_6121)?data_in_org271:10'b0)|
    ((_net_2129)?data_in_org268:10'b0);
   assign  _add_map_x_111_moto_org_near2 = ((_net_6120)?data_in_org238:10'b0)|
    ((_net_2128)?data_in_org237:10'b0);
   assign  _add_map_x_111_moto_org_near3 = ((_net_6119)?data_in_org302:10'b0)|
    ((_net_2127)?data_in_org301:10'b0);
   assign  _add_map_x_111_moto_org = ((_net_6118)?data_in_org270:10'b0)|
    ((_net_2126)?data_in_org269:10'b0);
   assign  _add_map_x_111_sg_up = ((_net_6117)?sg_in269:2'b0)|
    ((_net_2125)?sg_in270:2'b0);
   assign  _add_map_x_111_sg_down = ((_net_6116)?sg_in271:2'b0)|
    ((_net_2124)?sg_in268:2'b0);
   assign  _add_map_x_111_sg_left = ((_net_6114)?sg_in302:2'b0)|
    ((_net_2122)?sg_in301:2'b0);
   assign  _add_map_x_111_sg_right = ((_net_6115)?sg_in238:2'b0)|
    ((_net_2123)?sg_in237:2'b0);
   assign  _add_map_x_111_wall_t_in = dig_w;
   assign  _add_map_x_111_moto = ((_net_6112)?data_in270:10'b0)|
    ((_net_2120)?data_in269:10'b0);
   assign  _add_map_x_111_up = ((_net_6111)?data_in269:10'b0)|
    ((_net_2119)?data_in270:10'b0);
   assign  _add_map_x_111_right = ((_net_6110)?data_in271:10'b0)|
    ((_net_2118)?data_in268:10'b0);
   assign  _add_map_x_111_down = ((_net_6109)?data_in238:10'b0)|
    ((_net_2117)?data_in237:10'b0);
   assign  _add_map_x_111_left = ((_net_6108)?data_in302:10'b0)|
    ((_net_2116)?data_in301:10'b0);
   assign  _add_map_x_111_start = start;
   assign  _add_map_x_111_goal = goal;
   assign  _add_map_x_111_now = ((_net_6105)?10'b0100001110:10'b0)|
    ((_net_2113)?10'b0100001101:10'b0);
   assign  _add_map_x_111_add_exe = (_net_6104|_net_2112);
   assign  _add_map_x_111_p_reset = p_reset;
   assign  _add_map_x_111_m_clock = m_clock;
   assign  _add_map_x_110_moto_org_near = ((_net_6103)?data_in_org267:10'b0)|
    ((_net_2111)?data_in_org268:10'b0);
   assign  _add_map_x_110_moto_org_near1 = ((_net_6102)?data_in_org269:10'b0)|
    ((_net_2110)?data_in_org266:10'b0);
   assign  _add_map_x_110_moto_org_near2 = ((_net_6101)?data_in_org236:10'b0)|
    ((_net_2109)?data_in_org235:10'b0);
   assign  _add_map_x_110_moto_org_near3 = ((_net_6100)?data_in_org300:10'b0)|
    ((_net_2108)?data_in_org299:10'b0);
   assign  _add_map_x_110_moto_org = ((_net_6099)?data_in_org268:10'b0)|
    ((_net_2107)?data_in_org267:10'b0);
   assign  _add_map_x_110_sg_up = ((_net_6098)?sg_in267:2'b0)|
    ((_net_2106)?sg_in268:2'b0);
   assign  _add_map_x_110_sg_down = ((_net_6097)?sg_in269:2'b0)|
    ((_net_2105)?sg_in266:2'b0);
   assign  _add_map_x_110_sg_left = ((_net_6095)?sg_in300:2'b0)|
    ((_net_2103)?sg_in299:2'b0);
   assign  _add_map_x_110_sg_right = ((_net_6096)?sg_in236:2'b0)|
    ((_net_2104)?sg_in235:2'b0);
   assign  _add_map_x_110_wall_t_in = dig_w;
   assign  _add_map_x_110_moto = ((_net_6093)?data_in268:10'b0)|
    ((_net_2101)?data_in267:10'b0);
   assign  _add_map_x_110_up = ((_net_6092)?data_in267:10'b0)|
    ((_net_2100)?data_in268:10'b0);
   assign  _add_map_x_110_right = ((_net_6091)?data_in269:10'b0)|
    ((_net_2099)?data_in266:10'b0);
   assign  _add_map_x_110_down = ((_net_6090)?data_in236:10'b0)|
    ((_net_2098)?data_in235:10'b0);
   assign  _add_map_x_110_left = ((_net_6089)?data_in300:10'b0)|
    ((_net_2097)?data_in299:10'b0);
   assign  _add_map_x_110_start = start;
   assign  _add_map_x_110_goal = goal;
   assign  _add_map_x_110_now = ((_net_6086)?10'b0100001100:10'b0)|
    ((_net_2094)?10'b0100001011:10'b0);
   assign  _add_map_x_110_add_exe = (_net_6085|_net_2093);
   assign  _add_map_x_110_p_reset = p_reset;
   assign  _add_map_x_110_m_clock = m_clock;
   assign  _add_map_x_109_moto_org_near = ((_net_6084)?data_in_org265:10'b0)|
    ((_net_2092)?data_in_org266:10'b0);
   assign  _add_map_x_109_moto_org_near1 = ((_net_6083)?data_in_org267:10'b0)|
    ((_net_2091)?data_in_org264:10'b0);
   assign  _add_map_x_109_moto_org_near2 = ((_net_6082)?data_in_org234:10'b0)|
    ((_net_2090)?data_in_org233:10'b0);
   assign  _add_map_x_109_moto_org_near3 = ((_net_6081)?data_in_org298:10'b0)|
    ((_net_2089)?data_in_org297:10'b0);
   assign  _add_map_x_109_moto_org = ((_net_6080)?data_in_org266:10'b0)|
    ((_net_2088)?data_in_org265:10'b0);
   assign  _add_map_x_109_sg_up = ((_net_6079)?sg_in265:2'b0)|
    ((_net_2087)?sg_in266:2'b0);
   assign  _add_map_x_109_sg_down = ((_net_6078)?sg_in267:2'b0)|
    ((_net_2086)?sg_in264:2'b0);
   assign  _add_map_x_109_sg_left = ((_net_6076)?sg_in298:2'b0)|
    ((_net_2084)?sg_in297:2'b0);
   assign  _add_map_x_109_sg_right = ((_net_6077)?sg_in234:2'b0)|
    ((_net_2085)?sg_in233:2'b0);
   assign  _add_map_x_109_wall_t_in = dig_w;
   assign  _add_map_x_109_moto = ((_net_6074)?data_in266:10'b0)|
    ((_net_2082)?data_in265:10'b0);
   assign  _add_map_x_109_up = ((_net_6073)?data_in265:10'b0)|
    ((_net_2081)?data_in266:10'b0);
   assign  _add_map_x_109_right = ((_net_6072)?data_in267:10'b0)|
    ((_net_2080)?data_in264:10'b0);
   assign  _add_map_x_109_down = ((_net_6071)?data_in234:10'b0)|
    ((_net_2079)?data_in233:10'b0);
   assign  _add_map_x_109_left = ((_net_6070)?data_in298:10'b0)|
    ((_net_2078)?data_in297:10'b0);
   assign  _add_map_x_109_start = start;
   assign  _add_map_x_109_goal = goal;
   assign  _add_map_x_109_now = ((_net_6067)?10'b0100001010:10'b0)|
    ((_net_2075)?10'b0100001001:10'b0);
   assign  _add_map_x_109_add_exe = (_net_6066|_net_2074);
   assign  _add_map_x_109_p_reset = p_reset;
   assign  _add_map_x_109_m_clock = m_clock;
   assign  _add_map_x_108_moto_org_near = ((_net_6065)?data_in_org263:10'b0)|
    ((_net_2073)?data_in_org264:10'b0);
   assign  _add_map_x_108_moto_org_near1 = ((_net_6064)?data_in_org265:10'b0)|
    ((_net_2072)?data_in_org262:10'b0);
   assign  _add_map_x_108_moto_org_near2 = ((_net_6063)?data_in_org232:10'b0)|
    ((_net_2071)?data_in_org231:10'b0);
   assign  _add_map_x_108_moto_org_near3 = ((_net_6062)?data_in_org296:10'b0)|
    ((_net_2070)?data_in_org295:10'b0);
   assign  _add_map_x_108_moto_org = ((_net_6061)?data_in_org264:10'b0)|
    ((_net_2069)?data_in_org263:10'b0);
   assign  _add_map_x_108_sg_up = ((_net_6060)?sg_in263:2'b0)|
    ((_net_2068)?sg_in264:2'b0);
   assign  _add_map_x_108_sg_down = ((_net_6059)?sg_in265:2'b0)|
    ((_net_2067)?sg_in262:2'b0);
   assign  _add_map_x_108_sg_left = ((_net_6057)?sg_in296:2'b0)|
    ((_net_2065)?sg_in295:2'b0);
   assign  _add_map_x_108_sg_right = ((_net_6058)?sg_in232:2'b0)|
    ((_net_2066)?sg_in231:2'b0);
   assign  _add_map_x_108_wall_t_in = dig_w;
   assign  _add_map_x_108_moto = ((_net_6055)?data_in264:10'b0)|
    ((_net_2063)?data_in263:10'b0);
   assign  _add_map_x_108_up = ((_net_6054)?data_in263:10'b0)|
    ((_net_2062)?data_in264:10'b0);
   assign  _add_map_x_108_right = ((_net_6053)?data_in265:10'b0)|
    ((_net_2061)?data_in262:10'b0);
   assign  _add_map_x_108_down = ((_net_6052)?data_in232:10'b0)|
    ((_net_2060)?data_in231:10'b0);
   assign  _add_map_x_108_left = ((_net_6051)?data_in296:10'b0)|
    ((_net_2059)?data_in295:10'b0);
   assign  _add_map_x_108_start = start;
   assign  _add_map_x_108_goal = goal;
   assign  _add_map_x_108_now = ((_net_6048)?10'b0100001000:10'b0)|
    ((_net_2056)?10'b0100000111:10'b0);
   assign  _add_map_x_108_add_exe = (_net_6047|_net_2055);
   assign  _add_map_x_108_p_reset = p_reset;
   assign  _add_map_x_108_m_clock = m_clock;
   assign  _add_map_x_107_moto_org_near = ((_net_6046)?data_in_org261:10'b0)|
    ((_net_2054)?data_in_org262:10'b0);
   assign  _add_map_x_107_moto_org_near1 = ((_net_6045)?data_in_org263:10'b0)|
    ((_net_2053)?data_in_org260:10'b0);
   assign  _add_map_x_107_moto_org_near2 = ((_net_6044)?data_in_org230:10'b0)|
    ((_net_2052)?data_in_org229:10'b0);
   assign  _add_map_x_107_moto_org_near3 = ((_net_6043)?data_in_org294:10'b0)|
    ((_net_2051)?data_in_org293:10'b0);
   assign  _add_map_x_107_moto_org = ((_net_6042)?data_in_org262:10'b0)|
    ((_net_2050)?data_in_org261:10'b0);
   assign  _add_map_x_107_sg_up = ((_net_6041)?sg_in261:2'b0)|
    ((_net_2049)?sg_in262:2'b0);
   assign  _add_map_x_107_sg_down = ((_net_6040)?sg_in263:2'b0)|
    ((_net_2048)?sg_in260:2'b0);
   assign  _add_map_x_107_sg_left = ((_net_6038)?sg_in294:2'b0)|
    ((_net_2046)?sg_in293:2'b0);
   assign  _add_map_x_107_sg_right = ((_net_6039)?sg_in230:2'b0)|
    ((_net_2047)?sg_in229:2'b0);
   assign  _add_map_x_107_wall_t_in = dig_w;
   assign  _add_map_x_107_moto = ((_net_6036)?data_in262:10'b0)|
    ((_net_2044)?data_in261:10'b0);
   assign  _add_map_x_107_up = ((_net_6035)?data_in261:10'b0)|
    ((_net_2043)?data_in262:10'b0);
   assign  _add_map_x_107_right = ((_net_6034)?data_in263:10'b0)|
    ((_net_2042)?data_in260:10'b0);
   assign  _add_map_x_107_down = ((_net_6033)?data_in230:10'b0)|
    ((_net_2041)?data_in229:10'b0);
   assign  _add_map_x_107_left = ((_net_6032)?data_in294:10'b0)|
    ((_net_2040)?data_in293:10'b0);
   assign  _add_map_x_107_start = start;
   assign  _add_map_x_107_goal = goal;
   assign  _add_map_x_107_now = ((_net_6029)?10'b0100000110:10'b0)|
    ((_net_2037)?10'b0100000101:10'b0);
   assign  _add_map_x_107_add_exe = (_net_6028|_net_2036);
   assign  _add_map_x_107_p_reset = p_reset;
   assign  _add_map_x_107_m_clock = m_clock;
   assign  _add_map_x_106_moto_org_near = ((_net_6027)?data_in_org259:10'b0)|
    ((_net_2035)?data_in_org260:10'b0);
   assign  _add_map_x_106_moto_org_near1 = ((_net_6026)?data_in_org261:10'b0)|
    ((_net_2034)?data_in_org258:10'b0);
   assign  _add_map_x_106_moto_org_near2 = ((_net_6025)?data_in_org228:10'b0)|
    ((_net_2033)?data_in_org227:10'b0);
   assign  _add_map_x_106_moto_org_near3 = ((_net_6024)?data_in_org292:10'b0)|
    ((_net_2032)?data_in_org291:10'b0);
   assign  _add_map_x_106_moto_org = ((_net_6023)?data_in_org260:10'b0)|
    ((_net_2031)?data_in_org259:10'b0);
   assign  _add_map_x_106_sg_up = ((_net_6022)?sg_in259:2'b0)|
    ((_net_2030)?sg_in260:2'b0);
   assign  _add_map_x_106_sg_down = ((_net_6021)?sg_in261:2'b0)|
    ((_net_2029)?sg_in258:2'b0);
   assign  _add_map_x_106_sg_left = ((_net_6019)?sg_in292:2'b0)|
    ((_net_2027)?sg_in291:2'b0);
   assign  _add_map_x_106_sg_right = ((_net_6020)?sg_in228:2'b0)|
    ((_net_2028)?sg_in227:2'b0);
   assign  _add_map_x_106_wall_t_in = dig_w;
   assign  _add_map_x_106_moto = ((_net_6017)?data_in260:10'b0)|
    ((_net_2025)?data_in259:10'b0);
   assign  _add_map_x_106_up = ((_net_6016)?data_in259:10'b0)|
    ((_net_2024)?data_in260:10'b0);
   assign  _add_map_x_106_right = ((_net_6015)?data_in261:10'b0)|
    ((_net_2023)?data_in258:10'b0);
   assign  _add_map_x_106_down = ((_net_6014)?data_in228:10'b0)|
    ((_net_2022)?data_in227:10'b0);
   assign  _add_map_x_106_left = ((_net_6013)?data_in292:10'b0)|
    ((_net_2021)?data_in291:10'b0);
   assign  _add_map_x_106_start = start;
   assign  _add_map_x_106_goal = goal;
   assign  _add_map_x_106_now = ((_net_6010)?10'b0100000100:10'b0)|
    ((_net_2018)?10'b0100000011:10'b0);
   assign  _add_map_x_106_add_exe = (_net_6009|_net_2017);
   assign  _add_map_x_106_p_reset = p_reset;
   assign  _add_map_x_106_m_clock = m_clock;
   assign  _add_map_x_105_moto_org_near = ((_net_6008)?data_in_org257:10'b0)|
    ((_net_2016)?data_in_org258:10'b0);
   assign  _add_map_x_105_moto_org_near1 = ((_net_6007)?data_in_org259:10'b0)|
    ((_net_2015)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_105_moto_org_near2 = ((_net_6006)?data_in_org226:10'b0)|
    ((_net_2014)?data_in_org225:10'b0);
   assign  _add_map_x_105_moto_org_near3 = ((_net_6005)?data_in_org290:10'b0)|
    ((_net_2013)?data_in_org289:10'b0);
   assign  _add_map_x_105_moto_org = ((_net_6004)?data_in_org258:10'b0)|
    ((_net_2012)?data_in_org257:10'b0);
   assign  _add_map_x_105_sg_up = ((_net_6003)?sg_in257:2'b0)|
    ((_net_2011)?sg_in258:2'b0);
   assign  _add_map_x_105_sg_down = ((_net_6002)?sg_in259:2'b0)|
    ((_net_2010)?3'b000:2'b0);
   assign  _add_map_x_105_sg_left = ((_net_6000)?sg_in290:2'b0)|
    ((_net_2008)?sg_in289:2'b0);
   assign  _add_map_x_105_sg_right = ((_net_6001)?sg_in226:2'b0)|
    ((_net_2009)?sg_in225:2'b0);
   assign  _add_map_x_105_wall_t_in = dig_w;
   assign  _add_map_x_105_moto = ((_net_5998)?data_in258:10'b0)|
    ((_net_2006)?data_in257:10'b0);
   assign  _add_map_x_105_up = ((_net_5997)?data_in257:10'b0)|
    ((_net_2005)?data_in258:10'b0);
   assign  _add_map_x_105_right = ((_net_5996)?data_in259:10'b0)|
    ((_net_2004)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_105_down = ((_net_5995)?data_in226:10'b0)|
    ((_net_2003)?data_in225:10'b0);
   assign  _add_map_x_105_left = ((_net_5994)?data_in290:10'b0)|
    ((_net_2002)?data_in289:10'b0);
   assign  _add_map_x_105_start = start;
   assign  _add_map_x_105_goal = goal;
   assign  _add_map_x_105_now = ((_net_5991)?10'b0100000010:10'b0)|
    ((_net_1999)?10'b0100000001:10'b0);
   assign  _add_map_x_105_add_exe = (_net_5990|_net_1998);
   assign  _add_map_x_105_p_reset = p_reset;
   assign  _add_map_x_105_m_clock = m_clock;
   assign  _add_map_x_104_moto_org_near = ((_net_5989)?data_in_org254:10'b0)|
    ((_net_1997)?data_in_org253:10'b0);
   assign  _add_map_x_104_moto_org_near1 = ((_net_5988)?data_in_org252:10'b0)|
    ((_net_1996)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_104_moto_org_near2 = ((_net_5987)?data_in_org221:10'b0)|
    ((_net_1995)?data_in_org222:10'b0);
   assign  _add_map_x_104_moto_org_near3 = ((_net_5986)?data_in_org285:10'b0)|
    ((_net_1994)?data_in_org286:10'b0);
   assign  _add_map_x_104_moto_org = ((_net_5985)?data_in_org253:10'b0)|
    ((_net_1993)?data_in_org254:10'b0);
   assign  _add_map_x_104_sg_up = ((_net_5984)?sg_in254:2'b0)|
    ((_net_1992)?sg_in253:2'b0);
   assign  _add_map_x_104_sg_down = ((_net_5983)?sg_in221:2'b0)|
    ((_net_1991)?3'b000:2'b0);
   assign  _add_map_x_104_sg_left = ((_net_5981)?sg_in285:2'b0)|
    ((_net_1989)?sg_in286:2'b0);
   assign  _add_map_x_104_sg_right = ((_net_5982)?sg_in252:2'b0)|
    ((_net_1990)?sg_in222:2'b0);
   assign  _add_map_x_104_wall_t_in = dig_w;
   assign  _add_map_x_104_moto = ((_net_5979)?data_in253:10'b0)|
    ((_net_1987)?data_in254:10'b0);
   assign  _add_map_x_104_up = ((_net_5978)?data_in254:10'b0)|
    ((_net_1986)?data_in253:10'b0);
   assign  _add_map_x_104_right = ((_net_5977)?data_in252:10'b0)|
    ((_net_1985)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_104_down = ((_net_5976)?data_in221:10'b0)|
    ((_net_1984)?data_in222:10'b0);
   assign  _add_map_x_104_left = ((_net_5975)?data_in285:10'b0)|
    ((_net_1983)?data_in286:10'b0);
   assign  _add_map_x_104_start = start;
   assign  _add_map_x_104_goal = goal;
   assign  _add_map_x_104_now = ((_net_5972)?10'b0011111101:10'b0)|
    ((_net_1980)?10'b0011111110:10'b0);
   assign  _add_map_x_104_add_exe = (_net_5971|_net_1979);
   assign  _add_map_x_104_p_reset = p_reset;
   assign  _add_map_x_104_m_clock = m_clock;
   assign  _add_map_x_103_moto_org_near = ((_net_5970)?data_in_org252:10'b0)|
    ((_net_1978)?data_in_org251:10'b0);
   assign  _add_map_x_103_moto_org_near1 = ((_net_5969)?data_in_org250:10'b0)|
    ((_net_1977)?data_in_org253:10'b0);
   assign  _add_map_x_103_moto_org_near2 = ((_net_5968)?data_in_org219:10'b0)|
    ((_net_1976)?data_in_org220:10'b0);
   assign  _add_map_x_103_moto_org_near3 = ((_net_5967)?data_in_org283:10'b0)|
    ((_net_1975)?data_in_org284:10'b0);
   assign  _add_map_x_103_moto_org = ((_net_5966)?data_in_org251:10'b0)|
    ((_net_1974)?data_in_org252:10'b0);
   assign  _add_map_x_103_sg_up = ((_net_5965)?sg_in252:2'b0)|
    ((_net_1973)?sg_in251:2'b0);
   assign  _add_map_x_103_sg_down = ((_net_5964)?sg_in219:2'b0)|
    ((_net_1972)?sg_in253:2'b0);
   assign  _add_map_x_103_sg_left = ((_net_5962)?sg_in283:2'b0)|
    ((_net_1970)?sg_in284:2'b0);
   assign  _add_map_x_103_sg_right = ((_net_5963)?sg_in250:2'b0)|
    ((_net_1971)?sg_in220:2'b0);
   assign  _add_map_x_103_wall_t_in = dig_w;
   assign  _add_map_x_103_moto = ((_net_5960)?data_in251:10'b0)|
    ((_net_1968)?data_in252:10'b0);
   assign  _add_map_x_103_up = ((_net_5959)?data_in252:10'b0)|
    ((_net_1967)?data_in251:10'b0);
   assign  _add_map_x_103_right = ((_net_5958)?data_in250:10'b0)|
    ((_net_1966)?data_in253:10'b0);
   assign  _add_map_x_103_down = ((_net_5957)?data_in219:10'b0)|
    ((_net_1965)?data_in220:10'b0);
   assign  _add_map_x_103_left = ((_net_5956)?data_in283:10'b0)|
    ((_net_1964)?data_in284:10'b0);
   assign  _add_map_x_103_start = start;
   assign  _add_map_x_103_goal = goal;
   assign  _add_map_x_103_now = ((_net_5953)?10'b0011111011:10'b0)|
    ((_net_1961)?10'b0011111100:10'b0);
   assign  _add_map_x_103_add_exe = (_net_5952|_net_1960);
   assign  _add_map_x_103_p_reset = p_reset;
   assign  _add_map_x_103_m_clock = m_clock;
   assign  _add_map_x_102_moto_org_near = ((_net_5951)?data_in_org250:10'b0)|
    ((_net_1959)?data_in_org249:10'b0);
   assign  _add_map_x_102_moto_org_near1 = ((_net_5950)?data_in_org248:10'b0)|
    ((_net_1958)?data_in_org251:10'b0);
   assign  _add_map_x_102_moto_org_near2 = ((_net_5949)?data_in_org217:10'b0)|
    ((_net_1957)?data_in_org218:10'b0);
   assign  _add_map_x_102_moto_org_near3 = ((_net_5948)?data_in_org281:10'b0)|
    ((_net_1956)?data_in_org282:10'b0);
   assign  _add_map_x_102_moto_org = ((_net_5947)?data_in_org249:10'b0)|
    ((_net_1955)?data_in_org250:10'b0);
   assign  _add_map_x_102_sg_up = ((_net_5946)?sg_in250:2'b0)|
    ((_net_1954)?sg_in249:2'b0);
   assign  _add_map_x_102_sg_down = ((_net_5945)?sg_in217:2'b0)|
    ((_net_1953)?sg_in251:2'b0);
   assign  _add_map_x_102_sg_left = ((_net_5943)?sg_in281:2'b0)|
    ((_net_1951)?sg_in282:2'b0);
   assign  _add_map_x_102_sg_right = ((_net_5944)?sg_in248:2'b0)|
    ((_net_1952)?sg_in218:2'b0);
   assign  _add_map_x_102_wall_t_in = dig_w;
   assign  _add_map_x_102_moto = ((_net_5941)?data_in249:10'b0)|
    ((_net_1949)?data_in250:10'b0);
   assign  _add_map_x_102_up = ((_net_5940)?data_in250:10'b0)|
    ((_net_1948)?data_in249:10'b0);
   assign  _add_map_x_102_right = ((_net_5939)?data_in248:10'b0)|
    ((_net_1947)?data_in251:10'b0);
   assign  _add_map_x_102_down = ((_net_5938)?data_in217:10'b0)|
    ((_net_1946)?data_in218:10'b0);
   assign  _add_map_x_102_left = ((_net_5937)?data_in281:10'b0)|
    ((_net_1945)?data_in282:10'b0);
   assign  _add_map_x_102_start = start;
   assign  _add_map_x_102_goal = goal;
   assign  _add_map_x_102_now = ((_net_5934)?10'b0011111001:10'b0)|
    ((_net_1942)?10'b0011111010:10'b0);
   assign  _add_map_x_102_add_exe = (_net_5933|_net_1941);
   assign  _add_map_x_102_p_reset = p_reset;
   assign  _add_map_x_102_m_clock = m_clock;
   assign  _add_map_x_101_moto_org_near = ((_net_5932)?data_in_org248:10'b0)|
    ((_net_1940)?data_in_org247:10'b0);
   assign  _add_map_x_101_moto_org_near1 = ((_net_5931)?data_in_org246:10'b0)|
    ((_net_1939)?data_in_org249:10'b0);
   assign  _add_map_x_101_moto_org_near2 = ((_net_5930)?data_in_org215:10'b0)|
    ((_net_1938)?data_in_org216:10'b0);
   assign  _add_map_x_101_moto_org_near3 = ((_net_5929)?data_in_org279:10'b0)|
    ((_net_1937)?data_in_org280:10'b0);
   assign  _add_map_x_101_moto_org = ((_net_5928)?data_in_org247:10'b0)|
    ((_net_1936)?data_in_org248:10'b0);
   assign  _add_map_x_101_sg_up = ((_net_5927)?sg_in248:2'b0)|
    ((_net_1935)?sg_in247:2'b0);
   assign  _add_map_x_101_sg_down = ((_net_5926)?sg_in215:2'b0)|
    ((_net_1934)?sg_in249:2'b0);
   assign  _add_map_x_101_sg_left = ((_net_5924)?sg_in279:2'b0)|
    ((_net_1932)?sg_in280:2'b0);
   assign  _add_map_x_101_sg_right = ((_net_5925)?sg_in246:2'b0)|
    ((_net_1933)?sg_in216:2'b0);
   assign  _add_map_x_101_wall_t_in = dig_w;
   assign  _add_map_x_101_moto = ((_net_5922)?data_in247:10'b0)|
    ((_net_1930)?data_in248:10'b0);
   assign  _add_map_x_101_up = ((_net_5921)?data_in248:10'b0)|
    ((_net_1929)?data_in247:10'b0);
   assign  _add_map_x_101_right = ((_net_5920)?data_in246:10'b0)|
    ((_net_1928)?data_in249:10'b0);
   assign  _add_map_x_101_down = ((_net_5919)?data_in215:10'b0)|
    ((_net_1927)?data_in216:10'b0);
   assign  _add_map_x_101_left = ((_net_5918)?data_in279:10'b0)|
    ((_net_1926)?data_in280:10'b0);
   assign  _add_map_x_101_start = start;
   assign  _add_map_x_101_goal = goal;
   assign  _add_map_x_101_now = ((_net_5915)?10'b0011110111:10'b0)|
    ((_net_1923)?10'b0011111000:10'b0);
   assign  _add_map_x_101_add_exe = (_net_5914|_net_1922);
   assign  _add_map_x_101_p_reset = p_reset;
   assign  _add_map_x_101_m_clock = m_clock;
   assign  _add_map_x_100_moto_org_near = ((_net_5913)?data_in_org246:10'b0)|
    ((_net_1921)?data_in_org245:10'b0);
   assign  _add_map_x_100_moto_org_near1 = ((_net_5912)?data_in_org244:10'b0)|
    ((_net_1920)?data_in_org247:10'b0);
   assign  _add_map_x_100_moto_org_near2 = ((_net_5911)?data_in_org213:10'b0)|
    ((_net_1919)?data_in_org214:10'b0);
   assign  _add_map_x_100_moto_org_near3 = ((_net_5910)?data_in_org277:10'b0)|
    ((_net_1918)?data_in_org278:10'b0);
   assign  _add_map_x_100_moto_org = ((_net_5909)?data_in_org245:10'b0)|
    ((_net_1917)?data_in_org246:10'b0);
   assign  _add_map_x_100_sg_up = ((_net_5908)?sg_in246:2'b0)|
    ((_net_1916)?sg_in245:2'b0);
   assign  _add_map_x_100_sg_down = ((_net_5907)?sg_in213:2'b0)|
    ((_net_1915)?sg_in247:2'b0);
   assign  _add_map_x_100_sg_left = ((_net_5905)?sg_in277:2'b0)|
    ((_net_1913)?sg_in278:2'b0);
   assign  _add_map_x_100_sg_right = ((_net_5906)?sg_in244:2'b0)|
    ((_net_1914)?sg_in214:2'b0);
   assign  _add_map_x_100_wall_t_in = dig_w;
   assign  _add_map_x_100_moto = ((_net_5903)?data_in245:10'b0)|
    ((_net_1911)?data_in246:10'b0);
   assign  _add_map_x_100_up = ((_net_5902)?data_in246:10'b0)|
    ((_net_1910)?data_in245:10'b0);
   assign  _add_map_x_100_right = ((_net_5901)?data_in244:10'b0)|
    ((_net_1909)?data_in247:10'b0);
   assign  _add_map_x_100_down = ((_net_5900)?data_in213:10'b0)|
    ((_net_1908)?data_in214:10'b0);
   assign  _add_map_x_100_left = ((_net_5899)?data_in277:10'b0)|
    ((_net_1907)?data_in278:10'b0);
   assign  _add_map_x_100_start = start;
   assign  _add_map_x_100_goal = goal;
   assign  _add_map_x_100_now = ((_net_5896)?10'b0011110101:10'b0)|
    ((_net_1904)?10'b0011110110:10'b0);
   assign  _add_map_x_100_add_exe = (_net_5895|_net_1903);
   assign  _add_map_x_100_p_reset = p_reset;
   assign  _add_map_x_100_m_clock = m_clock;
   assign  _add_map_x_99_moto_org_near = ((_net_5894)?data_in_org244:10'b0)|
    ((_net_1902)?data_in_org243:10'b0);
   assign  _add_map_x_99_moto_org_near1 = ((_net_5893)?data_in_org242:10'b0)|
    ((_net_1901)?data_in_org245:10'b0);
   assign  _add_map_x_99_moto_org_near2 = ((_net_5892)?data_in_org211:10'b0)|
    ((_net_1900)?data_in_org212:10'b0);
   assign  _add_map_x_99_moto_org_near3 = ((_net_5891)?data_in_org275:10'b0)|
    ((_net_1899)?data_in_org276:10'b0);
   assign  _add_map_x_99_moto_org = ((_net_5890)?data_in_org243:10'b0)|
    ((_net_1898)?data_in_org244:10'b0);
   assign  _add_map_x_99_sg_up = ((_net_5889)?sg_in244:2'b0)|
    ((_net_1897)?sg_in243:2'b0);
   assign  _add_map_x_99_sg_down = ((_net_5888)?sg_in211:2'b0)|
    ((_net_1896)?sg_in245:2'b0);
   assign  _add_map_x_99_sg_left = ((_net_5886)?sg_in275:2'b0)|
    ((_net_1894)?sg_in276:2'b0);
   assign  _add_map_x_99_sg_right = ((_net_5887)?sg_in242:2'b0)|
    ((_net_1895)?sg_in212:2'b0);
   assign  _add_map_x_99_wall_t_in = dig_w;
   assign  _add_map_x_99_moto = ((_net_5884)?data_in243:10'b0)|
    ((_net_1892)?data_in244:10'b0);
   assign  _add_map_x_99_up = ((_net_5883)?data_in244:10'b0)|
    ((_net_1891)?data_in243:10'b0);
   assign  _add_map_x_99_right = ((_net_5882)?data_in242:10'b0)|
    ((_net_1890)?data_in245:10'b0);
   assign  _add_map_x_99_down = ((_net_5881)?data_in211:10'b0)|
    ((_net_1889)?data_in212:10'b0);
   assign  _add_map_x_99_left = ((_net_5880)?data_in275:10'b0)|
    ((_net_1888)?data_in276:10'b0);
   assign  _add_map_x_99_start = start;
   assign  _add_map_x_99_goal = goal;
   assign  _add_map_x_99_now = ((_net_5877)?10'b0011110011:10'b0)|
    ((_net_1885)?10'b0011110100:10'b0);
   assign  _add_map_x_99_add_exe = (_net_5876|_net_1884);
   assign  _add_map_x_99_p_reset = p_reset;
   assign  _add_map_x_99_m_clock = m_clock;
   assign  _add_map_x_98_moto_org_near = ((_net_5875)?data_in_org242:10'b0)|
    ((_net_1883)?data_in_org241:10'b0);
   assign  _add_map_x_98_moto_org_near1 = ((_net_5874)?data_in_org240:10'b0)|
    ((_net_1882)?data_in_org243:10'b0);
   assign  _add_map_x_98_moto_org_near2 = ((_net_5873)?data_in_org209:10'b0)|
    ((_net_1881)?data_in_org210:10'b0);
   assign  _add_map_x_98_moto_org_near3 = ((_net_5872)?data_in_org273:10'b0)|
    ((_net_1880)?data_in_org274:10'b0);
   assign  _add_map_x_98_moto_org = ((_net_5871)?data_in_org241:10'b0)|
    ((_net_1879)?data_in_org242:10'b0);
   assign  _add_map_x_98_sg_up = ((_net_5870)?sg_in242:2'b0)|
    ((_net_1878)?sg_in241:2'b0);
   assign  _add_map_x_98_sg_down = ((_net_5869)?sg_in209:2'b0)|
    ((_net_1877)?sg_in243:2'b0);
   assign  _add_map_x_98_sg_left = ((_net_5867)?sg_in273:2'b0)|
    ((_net_1875)?sg_in274:2'b0);
   assign  _add_map_x_98_sg_right = ((_net_5868)?sg_in240:2'b0)|
    ((_net_1876)?sg_in210:2'b0);
   assign  _add_map_x_98_wall_t_in = dig_w;
   assign  _add_map_x_98_moto = ((_net_5865)?data_in241:10'b0)|
    ((_net_1873)?data_in242:10'b0);
   assign  _add_map_x_98_up = ((_net_5864)?data_in242:10'b0)|
    ((_net_1872)?data_in241:10'b0);
   assign  _add_map_x_98_right = ((_net_5863)?data_in240:10'b0)|
    ((_net_1871)?data_in243:10'b0);
   assign  _add_map_x_98_down = ((_net_5862)?data_in209:10'b0)|
    ((_net_1870)?data_in210:10'b0);
   assign  _add_map_x_98_left = ((_net_5861)?data_in273:10'b0)|
    ((_net_1869)?data_in274:10'b0);
   assign  _add_map_x_98_start = start;
   assign  _add_map_x_98_goal = goal;
   assign  _add_map_x_98_now = ((_net_5858)?10'b0011110001:10'b0)|
    ((_net_1866)?10'b0011110010:10'b0);
   assign  _add_map_x_98_add_exe = (_net_5857|_net_1865);
   assign  _add_map_x_98_p_reset = p_reset;
   assign  _add_map_x_98_m_clock = m_clock;
   assign  _add_map_x_97_moto_org_near = ((_net_5856)?data_in_org240:10'b0)|
    ((_net_1864)?data_in_org239:10'b0);
   assign  _add_map_x_97_moto_org_near1 = ((_net_5855)?data_in_org238:10'b0)|
    ((_net_1863)?data_in_org241:10'b0);
   assign  _add_map_x_97_moto_org_near2 = ((_net_5854)?data_in_org207:10'b0)|
    ((_net_1862)?data_in_org208:10'b0);
   assign  _add_map_x_97_moto_org_near3 = ((_net_5853)?data_in_org271:10'b0)|
    ((_net_1861)?data_in_org272:10'b0);
   assign  _add_map_x_97_moto_org = ((_net_5852)?data_in_org239:10'b0)|
    ((_net_1860)?data_in_org240:10'b0);
   assign  _add_map_x_97_sg_up = ((_net_5851)?sg_in240:2'b0)|
    ((_net_1859)?sg_in239:2'b0);
   assign  _add_map_x_97_sg_down = ((_net_5850)?sg_in207:2'b0)|
    ((_net_1858)?sg_in241:2'b0);
   assign  _add_map_x_97_sg_left = ((_net_5848)?sg_in271:2'b0)|
    ((_net_1856)?sg_in272:2'b0);
   assign  _add_map_x_97_sg_right = ((_net_5849)?sg_in238:2'b0)|
    ((_net_1857)?sg_in208:2'b0);
   assign  _add_map_x_97_wall_t_in = dig_w;
   assign  _add_map_x_97_moto = ((_net_5846)?data_in239:10'b0)|
    ((_net_1854)?data_in240:10'b0);
   assign  _add_map_x_97_up = ((_net_5845)?data_in240:10'b0)|
    ((_net_1853)?data_in239:10'b0);
   assign  _add_map_x_97_right = ((_net_5844)?data_in238:10'b0)|
    ((_net_1852)?data_in241:10'b0);
   assign  _add_map_x_97_down = ((_net_5843)?data_in207:10'b0)|
    ((_net_1851)?data_in208:10'b0);
   assign  _add_map_x_97_left = ((_net_5842)?data_in271:10'b0)|
    ((_net_1850)?data_in272:10'b0);
   assign  _add_map_x_97_start = start;
   assign  _add_map_x_97_goal = goal;
   assign  _add_map_x_97_now = ((_net_5839)?10'b0011101111:10'b0)|
    ((_net_1847)?10'b0011110000:10'b0);
   assign  _add_map_x_97_add_exe = (_net_5838|_net_1846);
   assign  _add_map_x_97_p_reset = p_reset;
   assign  _add_map_x_97_m_clock = m_clock;
   assign  _add_map_x_96_moto_org_near = ((_net_5837)?data_in_org238:10'b0)|
    ((_net_1845)?data_in_org237:10'b0);
   assign  _add_map_x_96_moto_org_near1 = ((_net_5836)?data_in_org236:10'b0)|
    ((_net_1844)?data_in_org239:10'b0);
   assign  _add_map_x_96_moto_org_near2 = ((_net_5835)?data_in_org205:10'b0)|
    ((_net_1843)?data_in_org206:10'b0);
   assign  _add_map_x_96_moto_org_near3 = ((_net_5834)?data_in_org269:10'b0)|
    ((_net_1842)?data_in_org270:10'b0);
   assign  _add_map_x_96_moto_org = ((_net_5833)?data_in_org237:10'b0)|
    ((_net_1841)?data_in_org238:10'b0);
   assign  _add_map_x_96_sg_up = ((_net_5832)?sg_in238:2'b0)|
    ((_net_1840)?sg_in237:2'b0);
   assign  _add_map_x_96_sg_down = ((_net_5831)?sg_in205:2'b0)|
    ((_net_1839)?sg_in239:2'b0);
   assign  _add_map_x_96_sg_left = ((_net_5829)?sg_in269:2'b0)|
    ((_net_1837)?sg_in270:2'b0);
   assign  _add_map_x_96_sg_right = ((_net_5830)?sg_in236:2'b0)|
    ((_net_1838)?sg_in206:2'b0);
   assign  _add_map_x_96_wall_t_in = dig_w;
   assign  _add_map_x_96_moto = ((_net_5827)?data_in237:10'b0)|
    ((_net_1835)?data_in238:10'b0);
   assign  _add_map_x_96_up = ((_net_5826)?data_in238:10'b0)|
    ((_net_1834)?data_in237:10'b0);
   assign  _add_map_x_96_right = ((_net_5825)?data_in236:10'b0)|
    ((_net_1833)?data_in239:10'b0);
   assign  _add_map_x_96_down = ((_net_5824)?data_in205:10'b0)|
    ((_net_1832)?data_in206:10'b0);
   assign  _add_map_x_96_left = ((_net_5823)?data_in269:10'b0)|
    ((_net_1831)?data_in270:10'b0);
   assign  _add_map_x_96_start = start;
   assign  _add_map_x_96_goal = goal;
   assign  _add_map_x_96_now = ((_net_5820)?10'b0011101101:10'b0)|
    ((_net_1828)?10'b0011101110:10'b0);
   assign  _add_map_x_96_add_exe = (_net_5819|_net_1827);
   assign  _add_map_x_96_p_reset = p_reset;
   assign  _add_map_x_96_m_clock = m_clock;
   assign  _add_map_x_95_moto_org_near = ((_net_5818)?data_in_org236:10'b0)|
    ((_net_1826)?data_in_org235:10'b0);
   assign  _add_map_x_95_moto_org_near1 = ((_net_5817)?data_in_org234:10'b0)|
    ((_net_1825)?data_in_org237:10'b0);
   assign  _add_map_x_95_moto_org_near2 = ((_net_5816)?data_in_org203:10'b0)|
    ((_net_1824)?data_in_org204:10'b0);
   assign  _add_map_x_95_moto_org_near3 = ((_net_5815)?data_in_org267:10'b0)|
    ((_net_1823)?data_in_org268:10'b0);
   assign  _add_map_x_95_moto_org = ((_net_5814)?data_in_org235:10'b0)|
    ((_net_1822)?data_in_org236:10'b0);
   assign  _add_map_x_95_sg_up = ((_net_5813)?sg_in236:2'b0)|
    ((_net_1821)?sg_in235:2'b0);
   assign  _add_map_x_95_sg_down = ((_net_5812)?sg_in203:2'b0)|
    ((_net_1820)?sg_in237:2'b0);
   assign  _add_map_x_95_sg_left = ((_net_5810)?sg_in267:2'b0)|
    ((_net_1818)?sg_in268:2'b0);
   assign  _add_map_x_95_sg_right = ((_net_5811)?sg_in234:2'b0)|
    ((_net_1819)?sg_in204:2'b0);
   assign  _add_map_x_95_wall_t_in = dig_w;
   assign  _add_map_x_95_moto = ((_net_5808)?data_in235:10'b0)|
    ((_net_1816)?data_in236:10'b0);
   assign  _add_map_x_95_up = ((_net_5807)?data_in236:10'b0)|
    ((_net_1815)?data_in235:10'b0);
   assign  _add_map_x_95_right = ((_net_5806)?data_in234:10'b0)|
    ((_net_1814)?data_in237:10'b0);
   assign  _add_map_x_95_down = ((_net_5805)?data_in203:10'b0)|
    ((_net_1813)?data_in204:10'b0);
   assign  _add_map_x_95_left = ((_net_5804)?data_in267:10'b0)|
    ((_net_1812)?data_in268:10'b0);
   assign  _add_map_x_95_start = start;
   assign  _add_map_x_95_goal = goal;
   assign  _add_map_x_95_now = ((_net_5801)?10'b0011101011:10'b0)|
    ((_net_1809)?10'b0011101100:10'b0);
   assign  _add_map_x_95_add_exe = (_net_5800|_net_1808);
   assign  _add_map_x_95_p_reset = p_reset;
   assign  _add_map_x_95_m_clock = m_clock;
   assign  _add_map_x_94_moto_org_near = ((_net_5799)?data_in_org234:10'b0)|
    ((_net_1807)?data_in_org233:10'b0);
   assign  _add_map_x_94_moto_org_near1 = ((_net_5798)?data_in_org232:10'b0)|
    ((_net_1806)?data_in_org235:10'b0);
   assign  _add_map_x_94_moto_org_near2 = ((_net_5797)?data_in_org201:10'b0)|
    ((_net_1805)?data_in_org202:10'b0);
   assign  _add_map_x_94_moto_org_near3 = ((_net_5796)?data_in_org265:10'b0)|
    ((_net_1804)?data_in_org266:10'b0);
   assign  _add_map_x_94_moto_org = ((_net_5795)?data_in_org233:10'b0)|
    ((_net_1803)?data_in_org234:10'b0);
   assign  _add_map_x_94_sg_up = ((_net_5794)?sg_in234:2'b0)|
    ((_net_1802)?sg_in233:2'b0);
   assign  _add_map_x_94_sg_down = ((_net_5793)?sg_in201:2'b0)|
    ((_net_1801)?sg_in235:2'b0);
   assign  _add_map_x_94_sg_left = ((_net_5791)?sg_in265:2'b0)|
    ((_net_1799)?sg_in266:2'b0);
   assign  _add_map_x_94_sg_right = ((_net_5792)?sg_in232:2'b0)|
    ((_net_1800)?sg_in202:2'b0);
   assign  _add_map_x_94_wall_t_in = dig_w;
   assign  _add_map_x_94_moto = ((_net_5789)?data_in233:10'b0)|
    ((_net_1797)?data_in234:10'b0);
   assign  _add_map_x_94_up = ((_net_5788)?data_in234:10'b0)|
    ((_net_1796)?data_in233:10'b0);
   assign  _add_map_x_94_right = ((_net_5787)?data_in232:10'b0)|
    ((_net_1795)?data_in235:10'b0);
   assign  _add_map_x_94_down = ((_net_5786)?data_in201:10'b0)|
    ((_net_1794)?data_in202:10'b0);
   assign  _add_map_x_94_left = ((_net_5785)?data_in265:10'b0)|
    ((_net_1793)?data_in266:10'b0);
   assign  _add_map_x_94_start = start;
   assign  _add_map_x_94_goal = goal;
   assign  _add_map_x_94_now = ((_net_5782)?10'b0011101001:10'b0)|
    ((_net_1790)?10'b0011101010:10'b0);
   assign  _add_map_x_94_add_exe = (_net_5781|_net_1789);
   assign  _add_map_x_94_p_reset = p_reset;
   assign  _add_map_x_94_m_clock = m_clock;
   assign  _add_map_x_93_moto_org_near = ((_net_5780)?data_in_org232:10'b0)|
    ((_net_1788)?data_in_org231:10'b0);
   assign  _add_map_x_93_moto_org_near1 = ((_net_5779)?data_in_org230:10'b0)|
    ((_net_1787)?data_in_org233:10'b0);
   assign  _add_map_x_93_moto_org_near2 = ((_net_5778)?data_in_org199:10'b0)|
    ((_net_1786)?data_in_org200:10'b0);
   assign  _add_map_x_93_moto_org_near3 = ((_net_5777)?data_in_org263:10'b0)|
    ((_net_1785)?data_in_org264:10'b0);
   assign  _add_map_x_93_moto_org = ((_net_5776)?data_in_org231:10'b0)|
    ((_net_1784)?data_in_org232:10'b0);
   assign  _add_map_x_93_sg_up = ((_net_5775)?sg_in232:2'b0)|
    ((_net_1783)?sg_in231:2'b0);
   assign  _add_map_x_93_sg_down = ((_net_5774)?sg_in199:2'b0)|
    ((_net_1782)?sg_in233:2'b0);
   assign  _add_map_x_93_sg_left = ((_net_5772)?sg_in263:2'b0)|
    ((_net_1780)?sg_in264:2'b0);
   assign  _add_map_x_93_sg_right = ((_net_5773)?sg_in230:2'b0)|
    ((_net_1781)?sg_in200:2'b0);
   assign  _add_map_x_93_wall_t_in = dig_w;
   assign  _add_map_x_93_moto = ((_net_5770)?data_in231:10'b0)|
    ((_net_1778)?data_in232:10'b0);
   assign  _add_map_x_93_up = ((_net_5769)?data_in232:10'b0)|
    ((_net_1777)?data_in231:10'b0);
   assign  _add_map_x_93_right = ((_net_5768)?data_in230:10'b0)|
    ((_net_1776)?data_in233:10'b0);
   assign  _add_map_x_93_down = ((_net_5767)?data_in199:10'b0)|
    ((_net_1775)?data_in200:10'b0);
   assign  _add_map_x_93_left = ((_net_5766)?data_in263:10'b0)|
    ((_net_1774)?data_in264:10'b0);
   assign  _add_map_x_93_start = start;
   assign  _add_map_x_93_goal = goal;
   assign  _add_map_x_93_now = ((_net_5763)?10'b0011100111:10'b0)|
    ((_net_1771)?10'b0011101000:10'b0);
   assign  _add_map_x_93_add_exe = (_net_5762|_net_1770);
   assign  _add_map_x_93_p_reset = p_reset;
   assign  _add_map_x_93_m_clock = m_clock;
   assign  _add_map_x_92_moto_org_near = ((_net_5761)?data_in_org230:10'b0)|
    ((_net_1769)?data_in_org229:10'b0);
   assign  _add_map_x_92_moto_org_near1 = ((_net_5760)?data_in_org228:10'b0)|
    ((_net_1768)?data_in_org231:10'b0);
   assign  _add_map_x_92_moto_org_near2 = ((_net_5759)?data_in_org197:10'b0)|
    ((_net_1767)?data_in_org198:10'b0);
   assign  _add_map_x_92_moto_org_near3 = ((_net_5758)?data_in_org261:10'b0)|
    ((_net_1766)?data_in_org262:10'b0);
   assign  _add_map_x_92_moto_org = ((_net_5757)?data_in_org229:10'b0)|
    ((_net_1765)?data_in_org230:10'b0);
   assign  _add_map_x_92_sg_up = ((_net_5756)?sg_in230:2'b0)|
    ((_net_1764)?sg_in229:2'b0);
   assign  _add_map_x_92_sg_down = ((_net_5755)?sg_in197:2'b0)|
    ((_net_1763)?sg_in231:2'b0);
   assign  _add_map_x_92_sg_left = ((_net_5753)?sg_in261:2'b0)|
    ((_net_1761)?sg_in262:2'b0);
   assign  _add_map_x_92_sg_right = ((_net_5754)?sg_in228:2'b0)|
    ((_net_1762)?sg_in198:2'b0);
   assign  _add_map_x_92_wall_t_in = dig_w;
   assign  _add_map_x_92_moto = ((_net_5751)?data_in229:10'b0)|
    ((_net_1759)?data_in230:10'b0);
   assign  _add_map_x_92_up = ((_net_5750)?data_in230:10'b0)|
    ((_net_1758)?data_in229:10'b0);
   assign  _add_map_x_92_right = ((_net_5749)?data_in228:10'b0)|
    ((_net_1757)?data_in231:10'b0);
   assign  _add_map_x_92_down = ((_net_5748)?data_in197:10'b0)|
    ((_net_1756)?data_in198:10'b0);
   assign  _add_map_x_92_left = ((_net_5747)?data_in261:10'b0)|
    ((_net_1755)?data_in262:10'b0);
   assign  _add_map_x_92_start = start;
   assign  _add_map_x_92_goal = goal;
   assign  _add_map_x_92_now = ((_net_5744)?10'b0011100101:10'b0)|
    ((_net_1752)?10'b0011100110:10'b0);
   assign  _add_map_x_92_add_exe = (_net_5743|_net_1751);
   assign  _add_map_x_92_p_reset = p_reset;
   assign  _add_map_x_92_m_clock = m_clock;
   assign  _add_map_x_91_moto_org_near = ((_net_5742)?data_in_org228:10'b0)|
    ((_net_1750)?data_in_org227:10'b0);
   assign  _add_map_x_91_moto_org_near1 = ((_net_5741)?data_in_org226:10'b0)|
    ((_net_1749)?data_in_org229:10'b0);
   assign  _add_map_x_91_moto_org_near2 = ((_net_5740)?data_in_org195:10'b0)|
    ((_net_1748)?data_in_org196:10'b0);
   assign  _add_map_x_91_moto_org_near3 = ((_net_5739)?data_in_org259:10'b0)|
    ((_net_1747)?data_in_org260:10'b0);
   assign  _add_map_x_91_moto_org = ((_net_5738)?data_in_org227:10'b0)|
    ((_net_1746)?data_in_org228:10'b0);
   assign  _add_map_x_91_sg_up = ((_net_5737)?sg_in228:2'b0)|
    ((_net_1745)?sg_in227:2'b0);
   assign  _add_map_x_91_sg_down = ((_net_5736)?sg_in195:2'b0)|
    ((_net_1744)?sg_in229:2'b0);
   assign  _add_map_x_91_sg_left = ((_net_5734)?sg_in259:2'b0)|
    ((_net_1742)?sg_in260:2'b0);
   assign  _add_map_x_91_sg_right = ((_net_5735)?sg_in226:2'b0)|
    ((_net_1743)?sg_in196:2'b0);
   assign  _add_map_x_91_wall_t_in = dig_w;
   assign  _add_map_x_91_moto = ((_net_5732)?data_in227:10'b0)|
    ((_net_1740)?data_in228:10'b0);
   assign  _add_map_x_91_up = ((_net_5731)?data_in228:10'b0)|
    ((_net_1739)?data_in227:10'b0);
   assign  _add_map_x_91_right = ((_net_5730)?data_in226:10'b0)|
    ((_net_1738)?data_in229:10'b0);
   assign  _add_map_x_91_down = ((_net_5729)?data_in195:10'b0)|
    ((_net_1737)?data_in196:10'b0);
   assign  _add_map_x_91_left = ((_net_5728)?data_in259:10'b0)|
    ((_net_1736)?data_in260:10'b0);
   assign  _add_map_x_91_start = start;
   assign  _add_map_x_91_goal = goal;
   assign  _add_map_x_91_now = ((_net_5725)?10'b0011100011:10'b0)|
    ((_net_1733)?10'b0011100100:10'b0);
   assign  _add_map_x_91_add_exe = (_net_5724|_net_1732);
   assign  _add_map_x_91_p_reset = p_reset;
   assign  _add_map_x_91_m_clock = m_clock;
   assign  _add_map_x_90_moto_org_near = ((_net_5723)?data_in_org226:10'b0)|
    ((_net_1731)?data_in_org225:10'b0);
   assign  _add_map_x_90_moto_org_near1 = ((_net_5722)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1730)?data_in_org227:10'b0);
   assign  _add_map_x_90_moto_org_near2 = ((_net_5721)?data_in_org193:10'b0)|
    ((_net_1729)?data_in_org194:10'b0);
   assign  _add_map_x_90_moto_org_near3 = ((_net_5720)?data_in_org257:10'b0)|
    ((_net_1728)?data_in_org258:10'b0);
   assign  _add_map_x_90_moto_org = ((_net_5719)?data_in_org225:10'b0)|
    ((_net_1727)?data_in_org226:10'b0);
   assign  _add_map_x_90_sg_up = ((_net_5718)?sg_in226:2'b0)|
    ((_net_1726)?sg_in225:2'b0);
   assign  _add_map_x_90_sg_down = ((_net_5717)?sg_in193:2'b0)|
    ((_net_1725)?sg_in227:2'b0);
   assign  _add_map_x_90_sg_left = ((_net_5715)?sg_in257:2'b0)|
    ((_net_1723)?sg_in258:2'b0);
   assign  _add_map_x_90_sg_right = ((_net_5716)?3'b000:2'b0)|
    ((_net_1724)?sg_in194:2'b0);
   assign  _add_map_x_90_wall_t_in = dig_w;
   assign  _add_map_x_90_moto = ((_net_5713)?data_in225:10'b0)|
    ((_net_1721)?data_in226:10'b0);
   assign  _add_map_x_90_up = ((_net_5712)?data_in226:10'b0)|
    ((_net_1720)?data_in225:10'b0);
   assign  _add_map_x_90_right = ((_net_5711)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1719)?data_in227:10'b0);
   assign  _add_map_x_90_down = ((_net_5710)?data_in193:10'b0)|
    ((_net_1718)?data_in194:10'b0);
   assign  _add_map_x_90_left = ((_net_5709)?data_in257:10'b0)|
    ((_net_1717)?data_in258:10'b0);
   assign  _add_map_x_90_start = start;
   assign  _add_map_x_90_goal = goal;
   assign  _add_map_x_90_now = ((_net_5706)?10'b0011100001:10'b0)|
    ((_net_1714)?10'b0011100010:10'b0);
   assign  _add_map_x_90_add_exe = (_net_5705|_net_1713);
   assign  _add_map_x_90_p_reset = p_reset;
   assign  _add_map_x_90_m_clock = m_clock;
   assign  _add_map_x_89_moto_org_near = ((_net_5704)?data_in_org221:10'b0)|
    ((_net_1712)?data_in_org222:10'b0);
   assign  _add_map_x_89_moto_org_near1 = ((_net_5703)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1711)?data_in_org220:10'b0);
   assign  _add_map_x_89_moto_org_near2 = ((_net_5702)?data_in_org190:10'b0)|
    ((_net_1710)?data_in_org189:10'b0);
   assign  _add_map_x_89_moto_org_near3 = ((_net_5701)?data_in_org254:10'b0)|
    ((_net_1709)?data_in_org253:10'b0);
   assign  _add_map_x_89_moto_org = ((_net_5700)?data_in_org222:10'b0)|
    ((_net_1708)?data_in_org221:10'b0);
   assign  _add_map_x_89_sg_up = ((_net_5699)?sg_in221:2'b0)|
    ((_net_1707)?sg_in222:2'b0);
   assign  _add_map_x_89_sg_down = ((_net_5698)?3'b000:2'b0)|
    ((_net_1706)?sg_in220:2'b0);
   assign  _add_map_x_89_sg_left = ((_net_5696)?sg_in254:2'b0)|
    ((_net_1704)?sg_in253:2'b0);
   assign  _add_map_x_89_sg_right = ((_net_5697)?sg_in190:2'b0)|
    ((_net_1705)?sg_in189:2'b0);
   assign  _add_map_x_89_wall_t_in = dig_w;
   assign  _add_map_x_89_moto = ((_net_5694)?data_in222:10'b0)|
    ((_net_1702)?data_in221:10'b0);
   assign  _add_map_x_89_up = ((_net_5693)?data_in221:10'b0)|
    ((_net_1701)?data_in222:10'b0);
   assign  _add_map_x_89_right = ((_net_5692)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1700)?data_in220:10'b0);
   assign  _add_map_x_89_down = ((_net_5691)?data_in190:10'b0)|
    ((_net_1699)?data_in189:10'b0);
   assign  _add_map_x_89_left = ((_net_5690)?data_in254:10'b0)|
    ((_net_1698)?data_in253:10'b0);
   assign  _add_map_x_89_start = start;
   assign  _add_map_x_89_goal = goal;
   assign  _add_map_x_89_now = ((_net_5687)?10'b0011011110:10'b0)|
    ((_net_1695)?10'b0011011101:10'b0);
   assign  _add_map_x_89_add_exe = (_net_5686|_net_1694);
   assign  _add_map_x_89_p_reset = p_reset;
   assign  _add_map_x_89_m_clock = m_clock;
   assign  _add_map_x_88_moto_org_near = ((_net_5685)?data_in_org219:10'b0)|
    ((_net_1693)?data_in_org220:10'b0);
   assign  _add_map_x_88_moto_org_near1 = ((_net_5684)?data_in_org221:10'b0)|
    ((_net_1692)?data_in_org218:10'b0);
   assign  _add_map_x_88_moto_org_near2 = ((_net_5683)?data_in_org188:10'b0)|
    ((_net_1691)?data_in_org187:10'b0);
   assign  _add_map_x_88_moto_org_near3 = ((_net_5682)?data_in_org252:10'b0)|
    ((_net_1690)?data_in_org251:10'b0);
   assign  _add_map_x_88_moto_org = ((_net_5681)?data_in_org220:10'b0)|
    ((_net_1689)?data_in_org219:10'b0);
   assign  _add_map_x_88_sg_up = ((_net_5680)?sg_in219:2'b0)|
    ((_net_1688)?sg_in220:2'b0);
   assign  _add_map_x_88_sg_down = ((_net_5679)?sg_in221:2'b0)|
    ((_net_1687)?sg_in218:2'b0);
   assign  _add_map_x_88_sg_left = ((_net_5677)?sg_in252:2'b0)|
    ((_net_1685)?sg_in251:2'b0);
   assign  _add_map_x_88_sg_right = ((_net_5678)?sg_in188:2'b0)|
    ((_net_1686)?sg_in187:2'b0);
   assign  _add_map_x_88_wall_t_in = dig_w;
   assign  _add_map_x_88_moto = ((_net_5675)?data_in220:10'b0)|
    ((_net_1683)?data_in219:10'b0);
   assign  _add_map_x_88_up = ((_net_5674)?data_in219:10'b0)|
    ((_net_1682)?data_in220:10'b0);
   assign  _add_map_x_88_right = ((_net_5673)?data_in221:10'b0)|
    ((_net_1681)?data_in218:10'b0);
   assign  _add_map_x_88_down = ((_net_5672)?data_in188:10'b0)|
    ((_net_1680)?data_in187:10'b0);
   assign  _add_map_x_88_left = ((_net_5671)?data_in252:10'b0)|
    ((_net_1679)?data_in251:10'b0);
   assign  _add_map_x_88_start = start;
   assign  _add_map_x_88_goal = goal;
   assign  _add_map_x_88_now = ((_net_5668)?10'b0011011100:10'b0)|
    ((_net_1676)?10'b0011011011:10'b0);
   assign  _add_map_x_88_add_exe = (_net_5667|_net_1675);
   assign  _add_map_x_88_p_reset = p_reset;
   assign  _add_map_x_88_m_clock = m_clock;
   assign  _add_map_x_87_moto_org_near = ((_net_5666)?data_in_org217:10'b0)|
    ((_net_1674)?data_in_org218:10'b0);
   assign  _add_map_x_87_moto_org_near1 = ((_net_5665)?data_in_org219:10'b0)|
    ((_net_1673)?data_in_org216:10'b0);
   assign  _add_map_x_87_moto_org_near2 = ((_net_5664)?data_in_org186:10'b0)|
    ((_net_1672)?data_in_org185:10'b0);
   assign  _add_map_x_87_moto_org_near3 = ((_net_5663)?data_in_org250:10'b0)|
    ((_net_1671)?data_in_org249:10'b0);
   assign  _add_map_x_87_moto_org = ((_net_5662)?data_in_org218:10'b0)|
    ((_net_1670)?data_in_org217:10'b0);
   assign  _add_map_x_87_sg_up = ((_net_5661)?sg_in217:2'b0)|
    ((_net_1669)?sg_in218:2'b0);
   assign  _add_map_x_87_sg_down = ((_net_5660)?sg_in219:2'b0)|
    ((_net_1668)?sg_in216:2'b0);
   assign  _add_map_x_87_sg_left = ((_net_5658)?sg_in250:2'b0)|
    ((_net_1666)?sg_in249:2'b0);
   assign  _add_map_x_87_sg_right = ((_net_5659)?sg_in186:2'b0)|
    ((_net_1667)?sg_in185:2'b0);
   assign  _add_map_x_87_wall_t_in = dig_w;
   assign  _add_map_x_87_moto = ((_net_5656)?data_in218:10'b0)|
    ((_net_1664)?data_in217:10'b0);
   assign  _add_map_x_87_up = ((_net_5655)?data_in217:10'b0)|
    ((_net_1663)?data_in218:10'b0);
   assign  _add_map_x_87_right = ((_net_5654)?data_in219:10'b0)|
    ((_net_1662)?data_in216:10'b0);
   assign  _add_map_x_87_down = ((_net_5653)?data_in186:10'b0)|
    ((_net_1661)?data_in185:10'b0);
   assign  _add_map_x_87_left = ((_net_5652)?data_in250:10'b0)|
    ((_net_1660)?data_in249:10'b0);
   assign  _add_map_x_87_start = start;
   assign  _add_map_x_87_goal = goal;
   assign  _add_map_x_87_now = ((_net_5649)?10'b0011011010:10'b0)|
    ((_net_1657)?10'b0011011001:10'b0);
   assign  _add_map_x_87_add_exe = (_net_5648|_net_1656);
   assign  _add_map_x_87_p_reset = p_reset;
   assign  _add_map_x_87_m_clock = m_clock;
   assign  _add_map_x_86_moto_org_near = ((_net_5647)?data_in_org215:10'b0)|
    ((_net_1655)?data_in_org216:10'b0);
   assign  _add_map_x_86_moto_org_near1 = ((_net_5646)?data_in_org217:10'b0)|
    ((_net_1654)?data_in_org214:10'b0);
   assign  _add_map_x_86_moto_org_near2 = ((_net_5645)?data_in_org184:10'b0)|
    ((_net_1653)?data_in_org183:10'b0);
   assign  _add_map_x_86_moto_org_near3 = ((_net_5644)?data_in_org248:10'b0)|
    ((_net_1652)?data_in_org247:10'b0);
   assign  _add_map_x_86_moto_org = ((_net_5643)?data_in_org216:10'b0)|
    ((_net_1651)?data_in_org215:10'b0);
   assign  _add_map_x_86_sg_up = ((_net_5642)?sg_in215:2'b0)|
    ((_net_1650)?sg_in216:2'b0);
   assign  _add_map_x_86_sg_down = ((_net_5641)?sg_in217:2'b0)|
    ((_net_1649)?sg_in214:2'b0);
   assign  _add_map_x_86_sg_left = ((_net_5639)?sg_in248:2'b0)|
    ((_net_1647)?sg_in247:2'b0);
   assign  _add_map_x_86_sg_right = ((_net_5640)?sg_in184:2'b0)|
    ((_net_1648)?sg_in183:2'b0);
   assign  _add_map_x_86_wall_t_in = dig_w;
   assign  _add_map_x_86_moto = ((_net_5637)?data_in216:10'b0)|
    ((_net_1645)?data_in215:10'b0);
   assign  _add_map_x_86_up = ((_net_5636)?data_in215:10'b0)|
    ((_net_1644)?data_in216:10'b0);
   assign  _add_map_x_86_right = ((_net_5635)?data_in217:10'b0)|
    ((_net_1643)?data_in214:10'b0);
   assign  _add_map_x_86_down = ((_net_5634)?data_in184:10'b0)|
    ((_net_1642)?data_in183:10'b0);
   assign  _add_map_x_86_left = ((_net_5633)?data_in248:10'b0)|
    ((_net_1641)?data_in247:10'b0);
   assign  _add_map_x_86_start = start;
   assign  _add_map_x_86_goal = goal;
   assign  _add_map_x_86_now = ((_net_5630)?10'b0011011000:10'b0)|
    ((_net_1638)?10'b0011010111:10'b0);
   assign  _add_map_x_86_add_exe = (_net_5629|_net_1637);
   assign  _add_map_x_86_p_reset = p_reset;
   assign  _add_map_x_86_m_clock = m_clock;
   assign  _add_map_x_85_moto_org_near = ((_net_5628)?data_in_org213:10'b0)|
    ((_net_1636)?data_in_org214:10'b0);
   assign  _add_map_x_85_moto_org_near1 = ((_net_5627)?data_in_org215:10'b0)|
    ((_net_1635)?data_in_org212:10'b0);
   assign  _add_map_x_85_moto_org_near2 = ((_net_5626)?data_in_org182:10'b0)|
    ((_net_1634)?data_in_org181:10'b0);
   assign  _add_map_x_85_moto_org_near3 = ((_net_5625)?data_in_org246:10'b0)|
    ((_net_1633)?data_in_org245:10'b0);
   assign  _add_map_x_85_moto_org = ((_net_5624)?data_in_org214:10'b0)|
    ((_net_1632)?data_in_org213:10'b0);
   assign  _add_map_x_85_sg_up = ((_net_5623)?sg_in213:2'b0)|
    ((_net_1631)?sg_in214:2'b0);
   assign  _add_map_x_85_sg_down = ((_net_5622)?sg_in215:2'b0)|
    ((_net_1630)?sg_in212:2'b0);
   assign  _add_map_x_85_sg_left = ((_net_5620)?sg_in246:2'b0)|
    ((_net_1628)?sg_in245:2'b0);
   assign  _add_map_x_85_sg_right = ((_net_5621)?sg_in182:2'b0)|
    ((_net_1629)?sg_in181:2'b0);
   assign  _add_map_x_85_wall_t_in = dig_w;
   assign  _add_map_x_85_moto = ((_net_5618)?data_in214:10'b0)|
    ((_net_1626)?data_in213:10'b0);
   assign  _add_map_x_85_up = ((_net_5617)?data_in213:10'b0)|
    ((_net_1625)?data_in214:10'b0);
   assign  _add_map_x_85_right = ((_net_5616)?data_in215:10'b0)|
    ((_net_1624)?data_in212:10'b0);
   assign  _add_map_x_85_down = ((_net_5615)?data_in182:10'b0)|
    ((_net_1623)?data_in181:10'b0);
   assign  _add_map_x_85_left = ((_net_5614)?data_in246:10'b0)|
    ((_net_1622)?data_in245:10'b0);
   assign  _add_map_x_85_start = start;
   assign  _add_map_x_85_goal = goal;
   assign  _add_map_x_85_now = ((_net_5611)?10'b0011010110:10'b0)|
    ((_net_1619)?10'b0011010101:10'b0);
   assign  _add_map_x_85_add_exe = (_net_5610|_net_1618);
   assign  _add_map_x_85_p_reset = p_reset;
   assign  _add_map_x_85_m_clock = m_clock;
   assign  _add_map_x_84_moto_org_near = ((_net_5609)?data_in_org211:10'b0)|
    ((_net_1617)?data_in_org212:10'b0);
   assign  _add_map_x_84_moto_org_near1 = ((_net_5608)?data_in_org213:10'b0)|
    ((_net_1616)?data_in_org210:10'b0);
   assign  _add_map_x_84_moto_org_near2 = ((_net_5607)?data_in_org180:10'b0)|
    ((_net_1615)?data_in_org179:10'b0);
   assign  _add_map_x_84_moto_org_near3 = ((_net_5606)?data_in_org244:10'b0)|
    ((_net_1614)?data_in_org243:10'b0);
   assign  _add_map_x_84_moto_org = ((_net_5605)?data_in_org212:10'b0)|
    ((_net_1613)?data_in_org211:10'b0);
   assign  _add_map_x_84_sg_up = ((_net_5604)?sg_in211:2'b0)|
    ((_net_1612)?sg_in212:2'b0);
   assign  _add_map_x_84_sg_down = ((_net_5603)?sg_in213:2'b0)|
    ((_net_1611)?sg_in210:2'b0);
   assign  _add_map_x_84_sg_left = ((_net_5601)?sg_in244:2'b0)|
    ((_net_1609)?sg_in243:2'b0);
   assign  _add_map_x_84_sg_right = ((_net_5602)?sg_in180:2'b0)|
    ((_net_1610)?sg_in179:2'b0);
   assign  _add_map_x_84_wall_t_in = dig_w;
   assign  _add_map_x_84_moto = ((_net_5599)?data_in212:10'b0)|
    ((_net_1607)?data_in211:10'b0);
   assign  _add_map_x_84_up = ((_net_5598)?data_in211:10'b0)|
    ((_net_1606)?data_in212:10'b0);
   assign  _add_map_x_84_right = ((_net_5597)?data_in213:10'b0)|
    ((_net_1605)?data_in210:10'b0);
   assign  _add_map_x_84_down = ((_net_5596)?data_in180:10'b0)|
    ((_net_1604)?data_in179:10'b0);
   assign  _add_map_x_84_left = ((_net_5595)?data_in244:10'b0)|
    ((_net_1603)?data_in243:10'b0);
   assign  _add_map_x_84_start = start;
   assign  _add_map_x_84_goal = goal;
   assign  _add_map_x_84_now = ((_net_5592)?10'b0011010100:10'b0)|
    ((_net_1600)?10'b0011010011:10'b0);
   assign  _add_map_x_84_add_exe = (_net_5591|_net_1599);
   assign  _add_map_x_84_p_reset = p_reset;
   assign  _add_map_x_84_m_clock = m_clock;
   assign  _add_map_x_83_moto_org_near = ((_net_5590)?data_in_org209:10'b0)|
    ((_net_1598)?data_in_org210:10'b0);
   assign  _add_map_x_83_moto_org_near1 = ((_net_5589)?data_in_org211:10'b0)|
    ((_net_1597)?data_in_org208:10'b0);
   assign  _add_map_x_83_moto_org_near2 = ((_net_5588)?data_in_org178:10'b0)|
    ((_net_1596)?data_in_org177:10'b0);
   assign  _add_map_x_83_moto_org_near3 = ((_net_5587)?data_in_org242:10'b0)|
    ((_net_1595)?data_in_org241:10'b0);
   assign  _add_map_x_83_moto_org = ((_net_5586)?data_in_org210:10'b0)|
    ((_net_1594)?data_in_org209:10'b0);
   assign  _add_map_x_83_sg_up = ((_net_5585)?sg_in209:2'b0)|
    ((_net_1593)?sg_in210:2'b0);
   assign  _add_map_x_83_sg_down = ((_net_5584)?sg_in211:2'b0)|
    ((_net_1592)?sg_in208:2'b0);
   assign  _add_map_x_83_sg_left = ((_net_5582)?sg_in242:2'b0)|
    ((_net_1590)?sg_in241:2'b0);
   assign  _add_map_x_83_sg_right = ((_net_5583)?sg_in178:2'b0)|
    ((_net_1591)?sg_in177:2'b0);
   assign  _add_map_x_83_wall_t_in = dig_w;
   assign  _add_map_x_83_moto = ((_net_5580)?data_in210:10'b0)|
    ((_net_1588)?data_in209:10'b0);
   assign  _add_map_x_83_up = ((_net_5579)?data_in209:10'b0)|
    ((_net_1587)?data_in210:10'b0);
   assign  _add_map_x_83_right = ((_net_5578)?data_in211:10'b0)|
    ((_net_1586)?data_in208:10'b0);
   assign  _add_map_x_83_down = ((_net_5577)?data_in178:10'b0)|
    ((_net_1585)?data_in177:10'b0);
   assign  _add_map_x_83_left = ((_net_5576)?data_in242:10'b0)|
    ((_net_1584)?data_in241:10'b0);
   assign  _add_map_x_83_start = start;
   assign  _add_map_x_83_goal = goal;
   assign  _add_map_x_83_now = ((_net_5573)?10'b0011010010:10'b0)|
    ((_net_1581)?10'b0011010001:10'b0);
   assign  _add_map_x_83_add_exe = (_net_5572|_net_1580);
   assign  _add_map_x_83_p_reset = p_reset;
   assign  _add_map_x_83_m_clock = m_clock;
   assign  _add_map_x_82_moto_org_near = ((_net_5571)?data_in_org207:10'b0)|
    ((_net_1579)?data_in_org208:10'b0);
   assign  _add_map_x_82_moto_org_near1 = ((_net_5570)?data_in_org209:10'b0)|
    ((_net_1578)?data_in_org206:10'b0);
   assign  _add_map_x_82_moto_org_near2 = ((_net_5569)?data_in_org176:10'b0)|
    ((_net_1577)?data_in_org175:10'b0);
   assign  _add_map_x_82_moto_org_near3 = ((_net_5568)?data_in_org240:10'b0)|
    ((_net_1576)?data_in_org239:10'b0);
   assign  _add_map_x_82_moto_org = ((_net_5567)?data_in_org208:10'b0)|
    ((_net_1575)?data_in_org207:10'b0);
   assign  _add_map_x_82_sg_up = ((_net_5566)?sg_in207:2'b0)|
    ((_net_1574)?sg_in208:2'b0);
   assign  _add_map_x_82_sg_down = ((_net_5565)?sg_in209:2'b0)|
    ((_net_1573)?sg_in206:2'b0);
   assign  _add_map_x_82_sg_left = ((_net_5563)?sg_in240:2'b0)|
    ((_net_1571)?sg_in239:2'b0);
   assign  _add_map_x_82_sg_right = ((_net_5564)?sg_in176:2'b0)|
    ((_net_1572)?sg_in175:2'b0);
   assign  _add_map_x_82_wall_t_in = dig_w;
   assign  _add_map_x_82_moto = ((_net_5561)?data_in208:10'b0)|
    ((_net_1569)?data_in207:10'b0);
   assign  _add_map_x_82_up = ((_net_5560)?data_in207:10'b0)|
    ((_net_1568)?data_in208:10'b0);
   assign  _add_map_x_82_right = ((_net_5559)?data_in209:10'b0)|
    ((_net_1567)?data_in206:10'b0);
   assign  _add_map_x_82_down = ((_net_5558)?data_in176:10'b0)|
    ((_net_1566)?data_in175:10'b0);
   assign  _add_map_x_82_left = ((_net_5557)?data_in240:10'b0)|
    ((_net_1565)?data_in239:10'b0);
   assign  _add_map_x_82_start = start;
   assign  _add_map_x_82_goal = goal;
   assign  _add_map_x_82_now = ((_net_5554)?10'b0011010000:10'b0)|
    ((_net_1562)?10'b0011001111:10'b0);
   assign  _add_map_x_82_add_exe = (_net_5553|_net_1561);
   assign  _add_map_x_82_p_reset = p_reset;
   assign  _add_map_x_82_m_clock = m_clock;
   assign  _add_map_x_81_moto_org_near = ((_net_5552)?data_in_org205:10'b0)|
    ((_net_1560)?data_in_org206:10'b0);
   assign  _add_map_x_81_moto_org_near1 = ((_net_5551)?data_in_org207:10'b0)|
    ((_net_1559)?data_in_org204:10'b0);
   assign  _add_map_x_81_moto_org_near2 = ((_net_5550)?data_in_org174:10'b0)|
    ((_net_1558)?data_in_org173:10'b0);
   assign  _add_map_x_81_moto_org_near3 = ((_net_5549)?data_in_org238:10'b0)|
    ((_net_1557)?data_in_org237:10'b0);
   assign  _add_map_x_81_moto_org = ((_net_5548)?data_in_org206:10'b0)|
    ((_net_1556)?data_in_org205:10'b0);
   assign  _add_map_x_81_sg_up = ((_net_5547)?sg_in205:2'b0)|
    ((_net_1555)?sg_in206:2'b0);
   assign  _add_map_x_81_sg_down = ((_net_5546)?sg_in207:2'b0)|
    ((_net_1554)?sg_in204:2'b0);
   assign  _add_map_x_81_sg_left = ((_net_5544)?sg_in238:2'b0)|
    ((_net_1552)?sg_in237:2'b0);
   assign  _add_map_x_81_sg_right = ((_net_5545)?sg_in174:2'b0)|
    ((_net_1553)?sg_in173:2'b0);
   assign  _add_map_x_81_wall_t_in = dig_w;
   assign  _add_map_x_81_moto = ((_net_5542)?data_in206:10'b0)|
    ((_net_1550)?data_in205:10'b0);
   assign  _add_map_x_81_up = ((_net_5541)?data_in205:10'b0)|
    ((_net_1549)?data_in206:10'b0);
   assign  _add_map_x_81_right = ((_net_5540)?data_in207:10'b0)|
    ((_net_1548)?data_in204:10'b0);
   assign  _add_map_x_81_down = ((_net_5539)?data_in174:10'b0)|
    ((_net_1547)?data_in173:10'b0);
   assign  _add_map_x_81_left = ((_net_5538)?data_in238:10'b0)|
    ((_net_1546)?data_in237:10'b0);
   assign  _add_map_x_81_start = start;
   assign  _add_map_x_81_goal = goal;
   assign  _add_map_x_81_now = ((_net_5535)?10'b0011001110:10'b0)|
    ((_net_1543)?10'b0011001101:10'b0);
   assign  _add_map_x_81_add_exe = (_net_5534|_net_1542);
   assign  _add_map_x_81_p_reset = p_reset;
   assign  _add_map_x_81_m_clock = m_clock;
   assign  _add_map_x_80_moto_org_near = ((_net_5533)?data_in_org203:10'b0)|
    ((_net_1541)?data_in_org204:10'b0);
   assign  _add_map_x_80_moto_org_near1 = ((_net_5532)?data_in_org205:10'b0)|
    ((_net_1540)?data_in_org202:10'b0);
   assign  _add_map_x_80_moto_org_near2 = ((_net_5531)?data_in_org172:10'b0)|
    ((_net_1539)?data_in_org171:10'b0);
   assign  _add_map_x_80_moto_org_near3 = ((_net_5530)?data_in_org236:10'b0)|
    ((_net_1538)?data_in_org235:10'b0);
   assign  _add_map_x_80_moto_org = ((_net_5529)?data_in_org204:10'b0)|
    ((_net_1537)?data_in_org203:10'b0);
   assign  _add_map_x_80_sg_up = ((_net_5528)?sg_in203:2'b0)|
    ((_net_1536)?sg_in204:2'b0);
   assign  _add_map_x_80_sg_down = ((_net_5527)?sg_in205:2'b0)|
    ((_net_1535)?sg_in202:2'b0);
   assign  _add_map_x_80_sg_left = ((_net_5525)?sg_in236:2'b0)|
    ((_net_1533)?sg_in235:2'b0);
   assign  _add_map_x_80_sg_right = ((_net_5526)?sg_in172:2'b0)|
    ((_net_1534)?sg_in171:2'b0);
   assign  _add_map_x_80_wall_t_in = dig_w;
   assign  _add_map_x_80_moto = ((_net_5523)?data_in204:10'b0)|
    ((_net_1531)?data_in203:10'b0);
   assign  _add_map_x_80_up = ((_net_5522)?data_in203:10'b0)|
    ((_net_1530)?data_in204:10'b0);
   assign  _add_map_x_80_right = ((_net_5521)?data_in205:10'b0)|
    ((_net_1529)?data_in202:10'b0);
   assign  _add_map_x_80_down = ((_net_5520)?data_in172:10'b0)|
    ((_net_1528)?data_in171:10'b0);
   assign  _add_map_x_80_left = ((_net_5519)?data_in236:10'b0)|
    ((_net_1527)?data_in235:10'b0);
   assign  _add_map_x_80_start = start;
   assign  _add_map_x_80_goal = goal;
   assign  _add_map_x_80_now = ((_net_5516)?10'b0011001100:10'b0)|
    ((_net_1524)?10'b0011001011:10'b0);
   assign  _add_map_x_80_add_exe = (_net_5515|_net_1523);
   assign  _add_map_x_80_p_reset = p_reset;
   assign  _add_map_x_80_m_clock = m_clock;
   assign  _add_map_x_79_moto_org_near = ((_net_5514)?data_in_org201:10'b0)|
    ((_net_1522)?data_in_org202:10'b0);
   assign  _add_map_x_79_moto_org_near1 = ((_net_5513)?data_in_org203:10'b0)|
    ((_net_1521)?data_in_org200:10'b0);
   assign  _add_map_x_79_moto_org_near2 = ((_net_5512)?data_in_org170:10'b0)|
    ((_net_1520)?data_in_org169:10'b0);
   assign  _add_map_x_79_moto_org_near3 = ((_net_5511)?data_in_org234:10'b0)|
    ((_net_1519)?data_in_org233:10'b0);
   assign  _add_map_x_79_moto_org = ((_net_5510)?data_in_org202:10'b0)|
    ((_net_1518)?data_in_org201:10'b0);
   assign  _add_map_x_79_sg_up = ((_net_5509)?sg_in201:2'b0)|
    ((_net_1517)?sg_in202:2'b0);
   assign  _add_map_x_79_sg_down = ((_net_5508)?sg_in203:2'b0)|
    ((_net_1516)?sg_in200:2'b0);
   assign  _add_map_x_79_sg_left = ((_net_5506)?sg_in234:2'b0)|
    ((_net_1514)?sg_in233:2'b0);
   assign  _add_map_x_79_sg_right = ((_net_5507)?sg_in170:2'b0)|
    ((_net_1515)?sg_in169:2'b0);
   assign  _add_map_x_79_wall_t_in = dig_w;
   assign  _add_map_x_79_moto = ((_net_5504)?data_in202:10'b0)|
    ((_net_1512)?data_in201:10'b0);
   assign  _add_map_x_79_up = ((_net_5503)?data_in201:10'b0)|
    ((_net_1511)?data_in202:10'b0);
   assign  _add_map_x_79_right = ((_net_5502)?data_in203:10'b0)|
    ((_net_1510)?data_in200:10'b0);
   assign  _add_map_x_79_down = ((_net_5501)?data_in170:10'b0)|
    ((_net_1509)?data_in169:10'b0);
   assign  _add_map_x_79_left = ((_net_5500)?data_in234:10'b0)|
    ((_net_1508)?data_in233:10'b0);
   assign  _add_map_x_79_start = start;
   assign  _add_map_x_79_goal = goal;
   assign  _add_map_x_79_now = ((_net_5497)?10'b0011001010:10'b0)|
    ((_net_1505)?10'b0011001001:10'b0);
   assign  _add_map_x_79_add_exe = (_net_5496|_net_1504);
   assign  _add_map_x_79_p_reset = p_reset;
   assign  _add_map_x_79_m_clock = m_clock;
   assign  _add_map_x_78_moto_org_near = ((_net_5495)?data_in_org199:10'b0)|
    ((_net_1503)?data_in_org200:10'b0);
   assign  _add_map_x_78_moto_org_near1 = ((_net_5494)?data_in_org201:10'b0)|
    ((_net_1502)?data_in_org198:10'b0);
   assign  _add_map_x_78_moto_org_near2 = ((_net_5493)?data_in_org168:10'b0)|
    ((_net_1501)?data_in_org167:10'b0);
   assign  _add_map_x_78_moto_org_near3 = ((_net_5492)?data_in_org232:10'b0)|
    ((_net_1500)?data_in_org231:10'b0);
   assign  _add_map_x_78_moto_org = ((_net_5491)?data_in_org200:10'b0)|
    ((_net_1499)?data_in_org199:10'b0);
   assign  _add_map_x_78_sg_up = ((_net_5490)?sg_in199:2'b0)|
    ((_net_1498)?sg_in200:2'b0);
   assign  _add_map_x_78_sg_down = ((_net_5489)?sg_in201:2'b0)|
    ((_net_1497)?sg_in198:2'b0);
   assign  _add_map_x_78_sg_left = ((_net_5487)?sg_in232:2'b0)|
    ((_net_1495)?sg_in231:2'b0);
   assign  _add_map_x_78_sg_right = ((_net_5488)?sg_in168:2'b0)|
    ((_net_1496)?sg_in167:2'b0);
   assign  _add_map_x_78_wall_t_in = dig_w;
   assign  _add_map_x_78_moto = ((_net_5485)?data_in200:10'b0)|
    ((_net_1493)?data_in199:10'b0);
   assign  _add_map_x_78_up = ((_net_5484)?data_in199:10'b0)|
    ((_net_1492)?data_in200:10'b0);
   assign  _add_map_x_78_right = ((_net_5483)?data_in201:10'b0)|
    ((_net_1491)?data_in198:10'b0);
   assign  _add_map_x_78_down = ((_net_5482)?data_in168:10'b0)|
    ((_net_1490)?data_in167:10'b0);
   assign  _add_map_x_78_left = ((_net_5481)?data_in232:10'b0)|
    ((_net_1489)?data_in231:10'b0);
   assign  _add_map_x_78_start = start;
   assign  _add_map_x_78_goal = goal;
   assign  _add_map_x_78_now = ((_net_5478)?10'b0011001000:10'b0)|
    ((_net_1486)?10'b0011000111:10'b0);
   assign  _add_map_x_78_add_exe = (_net_5477|_net_1485);
   assign  _add_map_x_78_p_reset = p_reset;
   assign  _add_map_x_78_m_clock = m_clock;
   assign  _add_map_x_77_moto_org_near = ((_net_5476)?data_in_org197:10'b0)|
    ((_net_1484)?data_in_org198:10'b0);
   assign  _add_map_x_77_moto_org_near1 = ((_net_5475)?data_in_org199:10'b0)|
    ((_net_1483)?data_in_org196:10'b0);
   assign  _add_map_x_77_moto_org_near2 = ((_net_5474)?data_in_org166:10'b0)|
    ((_net_1482)?data_in_org165:10'b0);
   assign  _add_map_x_77_moto_org_near3 = ((_net_5473)?data_in_org230:10'b0)|
    ((_net_1481)?data_in_org229:10'b0);
   assign  _add_map_x_77_moto_org = ((_net_5472)?data_in_org198:10'b0)|
    ((_net_1480)?data_in_org197:10'b0);
   assign  _add_map_x_77_sg_up = ((_net_5471)?sg_in197:2'b0)|
    ((_net_1479)?sg_in198:2'b0);
   assign  _add_map_x_77_sg_down = ((_net_5470)?sg_in199:2'b0)|
    ((_net_1478)?sg_in196:2'b0);
   assign  _add_map_x_77_sg_left = ((_net_5468)?sg_in230:2'b0)|
    ((_net_1476)?sg_in229:2'b0);
   assign  _add_map_x_77_sg_right = ((_net_5469)?sg_in166:2'b0)|
    ((_net_1477)?sg_in165:2'b0);
   assign  _add_map_x_77_wall_t_in = dig_w;
   assign  _add_map_x_77_moto = ((_net_5466)?data_in198:10'b0)|
    ((_net_1474)?data_in197:10'b0);
   assign  _add_map_x_77_up = ((_net_5465)?data_in197:10'b0)|
    ((_net_1473)?data_in198:10'b0);
   assign  _add_map_x_77_right = ((_net_5464)?data_in199:10'b0)|
    ((_net_1472)?data_in196:10'b0);
   assign  _add_map_x_77_down = ((_net_5463)?data_in166:10'b0)|
    ((_net_1471)?data_in165:10'b0);
   assign  _add_map_x_77_left = ((_net_5462)?data_in230:10'b0)|
    ((_net_1470)?data_in229:10'b0);
   assign  _add_map_x_77_start = start;
   assign  _add_map_x_77_goal = goal;
   assign  _add_map_x_77_now = ((_net_5459)?10'b0011000110:10'b0)|
    ((_net_1467)?10'b0011000101:10'b0);
   assign  _add_map_x_77_add_exe = (_net_5458|_net_1466);
   assign  _add_map_x_77_p_reset = p_reset;
   assign  _add_map_x_77_m_clock = m_clock;
   assign  _add_map_x_76_moto_org_near = ((_net_5457)?data_in_org195:10'b0)|
    ((_net_1465)?data_in_org196:10'b0);
   assign  _add_map_x_76_moto_org_near1 = ((_net_5456)?data_in_org197:10'b0)|
    ((_net_1464)?data_in_org194:10'b0);
   assign  _add_map_x_76_moto_org_near2 = ((_net_5455)?data_in_org164:10'b0)|
    ((_net_1463)?data_in_org163:10'b0);
   assign  _add_map_x_76_moto_org_near3 = ((_net_5454)?data_in_org228:10'b0)|
    ((_net_1462)?data_in_org227:10'b0);
   assign  _add_map_x_76_moto_org = ((_net_5453)?data_in_org196:10'b0)|
    ((_net_1461)?data_in_org195:10'b0);
   assign  _add_map_x_76_sg_up = ((_net_5452)?sg_in195:2'b0)|
    ((_net_1460)?sg_in196:2'b0);
   assign  _add_map_x_76_sg_down = ((_net_5451)?sg_in197:2'b0)|
    ((_net_1459)?sg_in194:2'b0);
   assign  _add_map_x_76_sg_left = ((_net_5449)?sg_in228:2'b0)|
    ((_net_1457)?sg_in227:2'b0);
   assign  _add_map_x_76_sg_right = ((_net_5450)?sg_in164:2'b0)|
    ((_net_1458)?sg_in163:2'b0);
   assign  _add_map_x_76_wall_t_in = dig_w;
   assign  _add_map_x_76_moto = ((_net_5447)?data_in196:10'b0)|
    ((_net_1455)?data_in195:10'b0);
   assign  _add_map_x_76_up = ((_net_5446)?data_in195:10'b0)|
    ((_net_1454)?data_in196:10'b0);
   assign  _add_map_x_76_right = ((_net_5445)?data_in197:10'b0)|
    ((_net_1453)?data_in194:10'b0);
   assign  _add_map_x_76_down = ((_net_5444)?data_in164:10'b0)|
    ((_net_1452)?data_in163:10'b0);
   assign  _add_map_x_76_left = ((_net_5443)?data_in228:10'b0)|
    ((_net_1451)?data_in227:10'b0);
   assign  _add_map_x_76_start = start;
   assign  _add_map_x_76_goal = goal;
   assign  _add_map_x_76_now = ((_net_5440)?10'b0011000100:10'b0)|
    ((_net_1448)?10'b0011000011:10'b0);
   assign  _add_map_x_76_add_exe = (_net_5439|_net_1447);
   assign  _add_map_x_76_p_reset = p_reset;
   assign  _add_map_x_76_m_clock = m_clock;
   assign  _add_map_x_75_moto_org_near = ((_net_5438)?data_in_org193:10'b0)|
    ((_net_1446)?data_in_org194:10'b0);
   assign  _add_map_x_75_moto_org_near1 = ((_net_5437)?data_in_org195:10'b0)|
    ((_net_1445)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_75_moto_org_near2 = ((_net_5436)?data_in_org162:10'b0)|
    ((_net_1444)?data_in_org161:10'b0);
   assign  _add_map_x_75_moto_org_near3 = ((_net_5435)?data_in_org226:10'b0)|
    ((_net_1443)?data_in_org225:10'b0);
   assign  _add_map_x_75_moto_org = ((_net_5434)?data_in_org194:10'b0)|
    ((_net_1442)?data_in_org193:10'b0);
   assign  _add_map_x_75_sg_up = ((_net_5433)?sg_in193:2'b0)|
    ((_net_1441)?sg_in194:2'b0);
   assign  _add_map_x_75_sg_down = ((_net_5432)?sg_in195:2'b0)|
    ((_net_1440)?3'b000:2'b0);
   assign  _add_map_x_75_sg_left = ((_net_5430)?sg_in226:2'b0)|
    ((_net_1438)?sg_in225:2'b0);
   assign  _add_map_x_75_sg_right = ((_net_5431)?sg_in162:2'b0)|
    ((_net_1439)?sg_in161:2'b0);
   assign  _add_map_x_75_wall_t_in = dig_w;
   assign  _add_map_x_75_moto = ((_net_5428)?data_in194:10'b0)|
    ((_net_1436)?data_in193:10'b0);
   assign  _add_map_x_75_up = ((_net_5427)?data_in193:10'b0)|
    ((_net_1435)?data_in194:10'b0);
   assign  _add_map_x_75_right = ((_net_5426)?data_in195:10'b0)|
    ((_net_1434)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_75_down = ((_net_5425)?data_in162:10'b0)|
    ((_net_1433)?data_in161:10'b0);
   assign  _add_map_x_75_left = ((_net_5424)?data_in226:10'b0)|
    ((_net_1432)?data_in225:10'b0);
   assign  _add_map_x_75_start = start;
   assign  _add_map_x_75_goal = goal;
   assign  _add_map_x_75_now = ((_net_5421)?10'b0011000010:10'b0)|
    ((_net_1429)?10'b0011000001:10'b0);
   assign  _add_map_x_75_add_exe = (_net_5420|_net_1428);
   assign  _add_map_x_75_p_reset = p_reset;
   assign  _add_map_x_75_m_clock = m_clock;
   assign  _add_map_x_74_moto_org_near = ((_net_5419)?data_in_org190:10'b0)|
    ((_net_1427)?data_in_org189:10'b0);
   assign  _add_map_x_74_moto_org_near1 = ((_net_5418)?data_in_org188:10'b0)|
    ((_net_1426)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_74_moto_org_near2 = ((_net_5417)?data_in_org157:10'b0)|
    ((_net_1425)?data_in_org158:10'b0);
   assign  _add_map_x_74_moto_org_near3 = ((_net_5416)?data_in_org221:10'b0)|
    ((_net_1424)?data_in_org222:10'b0);
   assign  _add_map_x_74_moto_org = ((_net_5415)?data_in_org189:10'b0)|
    ((_net_1423)?data_in_org190:10'b0);
   assign  _add_map_x_74_sg_up = ((_net_5414)?sg_in190:2'b0)|
    ((_net_1422)?sg_in189:2'b0);
   assign  _add_map_x_74_sg_down = ((_net_5413)?sg_in157:2'b0)|
    ((_net_1421)?3'b000:2'b0);
   assign  _add_map_x_74_sg_left = ((_net_5411)?sg_in221:2'b0)|
    ((_net_1419)?sg_in222:2'b0);
   assign  _add_map_x_74_sg_right = ((_net_5412)?sg_in188:2'b0)|
    ((_net_1420)?sg_in158:2'b0);
   assign  _add_map_x_74_wall_t_in = dig_w;
   assign  _add_map_x_74_moto = ((_net_5409)?data_in189:10'b0)|
    ((_net_1417)?data_in190:10'b0);
   assign  _add_map_x_74_up = ((_net_5408)?data_in190:10'b0)|
    ((_net_1416)?data_in189:10'b0);
   assign  _add_map_x_74_right = ((_net_5407)?data_in188:10'b0)|
    ((_net_1415)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_74_down = ((_net_5406)?data_in157:10'b0)|
    ((_net_1414)?data_in158:10'b0);
   assign  _add_map_x_74_left = ((_net_5405)?data_in221:10'b0)|
    ((_net_1413)?data_in222:10'b0);
   assign  _add_map_x_74_start = start;
   assign  _add_map_x_74_goal = goal;
   assign  _add_map_x_74_now = ((_net_5402)?10'b0010111101:10'b0)|
    ((_net_1410)?10'b0010111110:10'b0);
   assign  _add_map_x_74_add_exe = (_net_5401|_net_1409);
   assign  _add_map_x_74_p_reset = p_reset;
   assign  _add_map_x_74_m_clock = m_clock;
   assign  _add_map_x_73_moto_org_near = ((_net_5400)?data_in_org188:10'b0)|
    ((_net_1408)?data_in_org187:10'b0);
   assign  _add_map_x_73_moto_org_near1 = ((_net_5399)?data_in_org186:10'b0)|
    ((_net_1407)?data_in_org189:10'b0);
   assign  _add_map_x_73_moto_org_near2 = ((_net_5398)?data_in_org155:10'b0)|
    ((_net_1406)?data_in_org156:10'b0);
   assign  _add_map_x_73_moto_org_near3 = ((_net_5397)?data_in_org219:10'b0)|
    ((_net_1405)?data_in_org220:10'b0);
   assign  _add_map_x_73_moto_org = ((_net_5396)?data_in_org187:10'b0)|
    ((_net_1404)?data_in_org188:10'b0);
   assign  _add_map_x_73_sg_up = ((_net_5395)?sg_in188:2'b0)|
    ((_net_1403)?sg_in187:2'b0);
   assign  _add_map_x_73_sg_down = ((_net_5394)?sg_in155:2'b0)|
    ((_net_1402)?sg_in189:2'b0);
   assign  _add_map_x_73_sg_left = ((_net_5392)?sg_in219:2'b0)|
    ((_net_1400)?sg_in220:2'b0);
   assign  _add_map_x_73_sg_right = ((_net_5393)?sg_in186:2'b0)|
    ((_net_1401)?sg_in156:2'b0);
   assign  _add_map_x_73_wall_t_in = dig_w;
   assign  _add_map_x_73_moto = ((_net_5390)?data_in187:10'b0)|
    ((_net_1398)?data_in188:10'b0);
   assign  _add_map_x_73_up = ((_net_5389)?data_in188:10'b0)|
    ((_net_1397)?data_in187:10'b0);
   assign  _add_map_x_73_right = ((_net_5388)?data_in186:10'b0)|
    ((_net_1396)?data_in189:10'b0);
   assign  _add_map_x_73_down = ((_net_5387)?data_in155:10'b0)|
    ((_net_1395)?data_in156:10'b0);
   assign  _add_map_x_73_left = ((_net_5386)?data_in219:10'b0)|
    ((_net_1394)?data_in220:10'b0);
   assign  _add_map_x_73_start = start;
   assign  _add_map_x_73_goal = goal;
   assign  _add_map_x_73_now = ((_net_5383)?10'b0010111011:10'b0)|
    ((_net_1391)?10'b0010111100:10'b0);
   assign  _add_map_x_73_add_exe = (_net_5382|_net_1390);
   assign  _add_map_x_73_p_reset = p_reset;
   assign  _add_map_x_73_m_clock = m_clock;
   assign  _add_map_x_72_moto_org_near = ((_net_5381)?data_in_org186:10'b0)|
    ((_net_1389)?data_in_org185:10'b0);
   assign  _add_map_x_72_moto_org_near1 = ((_net_5380)?data_in_org184:10'b0)|
    ((_net_1388)?data_in_org187:10'b0);
   assign  _add_map_x_72_moto_org_near2 = ((_net_5379)?data_in_org153:10'b0)|
    ((_net_1387)?data_in_org154:10'b0);
   assign  _add_map_x_72_moto_org_near3 = ((_net_5378)?data_in_org217:10'b0)|
    ((_net_1386)?data_in_org218:10'b0);
   assign  _add_map_x_72_moto_org = ((_net_5377)?data_in_org185:10'b0)|
    ((_net_1385)?data_in_org186:10'b0);
   assign  _add_map_x_72_sg_up = ((_net_5376)?sg_in186:2'b0)|
    ((_net_1384)?sg_in185:2'b0);
   assign  _add_map_x_72_sg_down = ((_net_5375)?sg_in153:2'b0)|
    ((_net_1383)?sg_in187:2'b0);
   assign  _add_map_x_72_sg_left = ((_net_5373)?sg_in217:2'b0)|
    ((_net_1381)?sg_in218:2'b0);
   assign  _add_map_x_72_sg_right = ((_net_5374)?sg_in184:2'b0)|
    ((_net_1382)?sg_in154:2'b0);
   assign  _add_map_x_72_wall_t_in = dig_w;
   assign  _add_map_x_72_moto = ((_net_5371)?data_in185:10'b0)|
    ((_net_1379)?data_in186:10'b0);
   assign  _add_map_x_72_up = ((_net_5370)?data_in186:10'b0)|
    ((_net_1378)?data_in185:10'b0);
   assign  _add_map_x_72_right = ((_net_5369)?data_in184:10'b0)|
    ((_net_1377)?data_in187:10'b0);
   assign  _add_map_x_72_down = ((_net_5368)?data_in153:10'b0)|
    ((_net_1376)?data_in154:10'b0);
   assign  _add_map_x_72_left = ((_net_5367)?data_in217:10'b0)|
    ((_net_1375)?data_in218:10'b0);
   assign  _add_map_x_72_start = start;
   assign  _add_map_x_72_goal = goal;
   assign  _add_map_x_72_now = ((_net_5364)?10'b0010111001:10'b0)|
    ((_net_1372)?10'b0010111010:10'b0);
   assign  _add_map_x_72_add_exe = (_net_5363|_net_1371);
   assign  _add_map_x_72_p_reset = p_reset;
   assign  _add_map_x_72_m_clock = m_clock;
   assign  _add_map_x_71_moto_org_near = ((_net_5362)?data_in_org184:10'b0)|
    ((_net_1370)?data_in_org183:10'b0);
   assign  _add_map_x_71_moto_org_near1 = ((_net_5361)?data_in_org182:10'b0)|
    ((_net_1369)?data_in_org185:10'b0);
   assign  _add_map_x_71_moto_org_near2 = ((_net_5360)?data_in_org151:10'b0)|
    ((_net_1368)?data_in_org152:10'b0);
   assign  _add_map_x_71_moto_org_near3 = ((_net_5359)?data_in_org215:10'b0)|
    ((_net_1367)?data_in_org216:10'b0);
   assign  _add_map_x_71_moto_org = ((_net_5358)?data_in_org183:10'b0)|
    ((_net_1366)?data_in_org184:10'b0);
   assign  _add_map_x_71_sg_up = ((_net_5357)?sg_in184:2'b0)|
    ((_net_1365)?sg_in183:2'b0);
   assign  _add_map_x_71_sg_down = ((_net_5356)?sg_in151:2'b0)|
    ((_net_1364)?sg_in185:2'b0);
   assign  _add_map_x_71_sg_left = ((_net_5354)?sg_in215:2'b0)|
    ((_net_1362)?sg_in216:2'b0);
   assign  _add_map_x_71_sg_right = ((_net_5355)?sg_in182:2'b0)|
    ((_net_1363)?sg_in152:2'b0);
   assign  _add_map_x_71_wall_t_in = dig_w;
   assign  _add_map_x_71_moto = ((_net_5352)?data_in183:10'b0)|
    ((_net_1360)?data_in184:10'b0);
   assign  _add_map_x_71_up = ((_net_5351)?data_in184:10'b0)|
    ((_net_1359)?data_in183:10'b0);
   assign  _add_map_x_71_right = ((_net_5350)?data_in182:10'b0)|
    ((_net_1358)?data_in185:10'b0);
   assign  _add_map_x_71_down = ((_net_5349)?data_in151:10'b0)|
    ((_net_1357)?data_in152:10'b0);
   assign  _add_map_x_71_left = ((_net_5348)?data_in215:10'b0)|
    ((_net_1356)?data_in216:10'b0);
   assign  _add_map_x_71_start = start;
   assign  _add_map_x_71_goal = goal;
   assign  _add_map_x_71_now = ((_net_5345)?10'b0010110111:10'b0)|
    ((_net_1353)?10'b0010111000:10'b0);
   assign  _add_map_x_71_add_exe = (_net_5344|_net_1352);
   assign  _add_map_x_71_p_reset = p_reset;
   assign  _add_map_x_71_m_clock = m_clock;
   assign  _add_map_x_70_moto_org_near = ((_net_5343)?data_in_org182:10'b0)|
    ((_net_1351)?data_in_org181:10'b0);
   assign  _add_map_x_70_moto_org_near1 = ((_net_5342)?data_in_org180:10'b0)|
    ((_net_1350)?data_in_org183:10'b0);
   assign  _add_map_x_70_moto_org_near2 = ((_net_5341)?data_in_org149:10'b0)|
    ((_net_1349)?data_in_org150:10'b0);
   assign  _add_map_x_70_moto_org_near3 = ((_net_5340)?data_in_org213:10'b0)|
    ((_net_1348)?data_in_org214:10'b0);
   assign  _add_map_x_70_moto_org = ((_net_5339)?data_in_org181:10'b0)|
    ((_net_1347)?data_in_org182:10'b0);
   assign  _add_map_x_70_sg_up = ((_net_5338)?sg_in182:2'b0)|
    ((_net_1346)?sg_in181:2'b0);
   assign  _add_map_x_70_sg_down = ((_net_5337)?sg_in149:2'b0)|
    ((_net_1345)?sg_in183:2'b0);
   assign  _add_map_x_70_sg_left = ((_net_5335)?sg_in213:2'b0)|
    ((_net_1343)?sg_in214:2'b0);
   assign  _add_map_x_70_sg_right = ((_net_5336)?sg_in180:2'b0)|
    ((_net_1344)?sg_in150:2'b0);
   assign  _add_map_x_70_wall_t_in = dig_w;
   assign  _add_map_x_70_moto = ((_net_5333)?data_in181:10'b0)|
    ((_net_1341)?data_in182:10'b0);
   assign  _add_map_x_70_up = ((_net_5332)?data_in182:10'b0)|
    ((_net_1340)?data_in181:10'b0);
   assign  _add_map_x_70_right = ((_net_5331)?data_in180:10'b0)|
    ((_net_1339)?data_in183:10'b0);
   assign  _add_map_x_70_down = ((_net_5330)?data_in149:10'b0)|
    ((_net_1338)?data_in150:10'b0);
   assign  _add_map_x_70_left = ((_net_5329)?data_in213:10'b0)|
    ((_net_1337)?data_in214:10'b0);
   assign  _add_map_x_70_start = start;
   assign  _add_map_x_70_goal = goal;
   assign  _add_map_x_70_now = ((_net_5326)?10'b0010110101:10'b0)|
    ((_net_1334)?10'b0010110110:10'b0);
   assign  _add_map_x_70_add_exe = (_net_5325|_net_1333);
   assign  _add_map_x_70_p_reset = p_reset;
   assign  _add_map_x_70_m_clock = m_clock;
   assign  _add_map_x_69_moto_org_near = ((_net_5324)?data_in_org180:10'b0)|
    ((_net_1332)?data_in_org179:10'b0);
   assign  _add_map_x_69_moto_org_near1 = ((_net_5323)?data_in_org178:10'b0)|
    ((_net_1331)?data_in_org181:10'b0);
   assign  _add_map_x_69_moto_org_near2 = ((_net_5322)?data_in_org147:10'b0)|
    ((_net_1330)?data_in_org148:10'b0);
   assign  _add_map_x_69_moto_org_near3 = ((_net_5321)?data_in_org211:10'b0)|
    ((_net_1329)?data_in_org212:10'b0);
   assign  _add_map_x_69_moto_org = ((_net_5320)?data_in_org179:10'b0)|
    ((_net_1328)?data_in_org180:10'b0);
   assign  _add_map_x_69_sg_up = ((_net_5319)?sg_in180:2'b0)|
    ((_net_1327)?sg_in179:2'b0);
   assign  _add_map_x_69_sg_down = ((_net_5318)?sg_in147:2'b0)|
    ((_net_1326)?sg_in181:2'b0);
   assign  _add_map_x_69_sg_left = ((_net_5316)?sg_in211:2'b0)|
    ((_net_1324)?sg_in212:2'b0);
   assign  _add_map_x_69_sg_right = ((_net_5317)?sg_in178:2'b0)|
    ((_net_1325)?sg_in148:2'b0);
   assign  _add_map_x_69_wall_t_in = dig_w;
   assign  _add_map_x_69_moto = ((_net_5314)?data_in179:10'b0)|
    ((_net_1322)?data_in180:10'b0);
   assign  _add_map_x_69_up = ((_net_5313)?data_in180:10'b0)|
    ((_net_1321)?data_in179:10'b0);
   assign  _add_map_x_69_right = ((_net_5312)?data_in178:10'b0)|
    ((_net_1320)?data_in181:10'b0);
   assign  _add_map_x_69_down = ((_net_5311)?data_in147:10'b0)|
    ((_net_1319)?data_in148:10'b0);
   assign  _add_map_x_69_left = ((_net_5310)?data_in211:10'b0)|
    ((_net_1318)?data_in212:10'b0);
   assign  _add_map_x_69_start = start;
   assign  _add_map_x_69_goal = goal;
   assign  _add_map_x_69_now = ((_net_5307)?10'b0010110011:10'b0)|
    ((_net_1315)?10'b0010110100:10'b0);
   assign  _add_map_x_69_add_exe = (_net_5306|_net_1314);
   assign  _add_map_x_69_p_reset = p_reset;
   assign  _add_map_x_69_m_clock = m_clock;
   assign  _add_map_x_68_moto_org_near = ((_net_5305)?data_in_org178:10'b0)|
    ((_net_1313)?data_in_org177:10'b0);
   assign  _add_map_x_68_moto_org_near1 = ((_net_5304)?data_in_org176:10'b0)|
    ((_net_1312)?data_in_org179:10'b0);
   assign  _add_map_x_68_moto_org_near2 = ((_net_5303)?data_in_org145:10'b0)|
    ((_net_1311)?data_in_org146:10'b0);
   assign  _add_map_x_68_moto_org_near3 = ((_net_5302)?data_in_org209:10'b0)|
    ((_net_1310)?data_in_org210:10'b0);
   assign  _add_map_x_68_moto_org = ((_net_5301)?data_in_org177:10'b0)|
    ((_net_1309)?data_in_org178:10'b0);
   assign  _add_map_x_68_sg_up = ((_net_5300)?sg_in178:2'b0)|
    ((_net_1308)?sg_in177:2'b0);
   assign  _add_map_x_68_sg_down = ((_net_5299)?sg_in145:2'b0)|
    ((_net_1307)?sg_in179:2'b0);
   assign  _add_map_x_68_sg_left = ((_net_5297)?sg_in209:2'b0)|
    ((_net_1305)?sg_in210:2'b0);
   assign  _add_map_x_68_sg_right = ((_net_5298)?sg_in176:2'b0)|
    ((_net_1306)?sg_in146:2'b0);
   assign  _add_map_x_68_wall_t_in = dig_w;
   assign  _add_map_x_68_moto = ((_net_5295)?data_in177:10'b0)|
    ((_net_1303)?data_in178:10'b0);
   assign  _add_map_x_68_up = ((_net_5294)?data_in178:10'b0)|
    ((_net_1302)?data_in177:10'b0);
   assign  _add_map_x_68_right = ((_net_5293)?data_in176:10'b0)|
    ((_net_1301)?data_in179:10'b0);
   assign  _add_map_x_68_down = ((_net_5292)?data_in145:10'b0)|
    ((_net_1300)?data_in146:10'b0);
   assign  _add_map_x_68_left = ((_net_5291)?data_in209:10'b0)|
    ((_net_1299)?data_in210:10'b0);
   assign  _add_map_x_68_start = start;
   assign  _add_map_x_68_goal = goal;
   assign  _add_map_x_68_now = ((_net_5288)?10'b0010110001:10'b0)|
    ((_net_1296)?10'b0010110010:10'b0);
   assign  _add_map_x_68_add_exe = (_net_5287|_net_1295);
   assign  _add_map_x_68_p_reset = p_reset;
   assign  _add_map_x_68_m_clock = m_clock;
   assign  _add_map_x_67_moto_org_near = ((_net_5286)?data_in_org176:10'b0)|
    ((_net_1294)?data_in_org175:10'b0);
   assign  _add_map_x_67_moto_org_near1 = ((_net_5285)?data_in_org174:10'b0)|
    ((_net_1293)?data_in_org177:10'b0);
   assign  _add_map_x_67_moto_org_near2 = ((_net_5284)?data_in_org143:10'b0)|
    ((_net_1292)?data_in_org144:10'b0);
   assign  _add_map_x_67_moto_org_near3 = ((_net_5283)?data_in_org207:10'b0)|
    ((_net_1291)?data_in_org208:10'b0);
   assign  _add_map_x_67_moto_org = ((_net_5282)?data_in_org175:10'b0)|
    ((_net_1290)?data_in_org176:10'b0);
   assign  _add_map_x_67_sg_up = ((_net_5281)?sg_in176:2'b0)|
    ((_net_1289)?sg_in175:2'b0);
   assign  _add_map_x_67_sg_down = ((_net_5280)?sg_in143:2'b0)|
    ((_net_1288)?sg_in177:2'b0);
   assign  _add_map_x_67_sg_left = ((_net_5278)?sg_in207:2'b0)|
    ((_net_1286)?sg_in208:2'b0);
   assign  _add_map_x_67_sg_right = ((_net_5279)?sg_in174:2'b0)|
    ((_net_1287)?sg_in144:2'b0);
   assign  _add_map_x_67_wall_t_in = dig_w;
   assign  _add_map_x_67_moto = ((_net_5276)?data_in175:10'b0)|
    ((_net_1284)?data_in176:10'b0);
   assign  _add_map_x_67_up = ((_net_5275)?data_in176:10'b0)|
    ((_net_1283)?data_in175:10'b0);
   assign  _add_map_x_67_right = ((_net_5274)?data_in174:10'b0)|
    ((_net_1282)?data_in177:10'b0);
   assign  _add_map_x_67_down = ((_net_5273)?data_in143:10'b0)|
    ((_net_1281)?data_in144:10'b0);
   assign  _add_map_x_67_left = ((_net_5272)?data_in207:10'b0)|
    ((_net_1280)?data_in208:10'b0);
   assign  _add_map_x_67_start = start;
   assign  _add_map_x_67_goal = goal;
   assign  _add_map_x_67_now = ((_net_5269)?10'b0010101111:10'b0)|
    ((_net_1277)?10'b0010110000:10'b0);
   assign  _add_map_x_67_add_exe = (_net_5268|_net_1276);
   assign  _add_map_x_67_p_reset = p_reset;
   assign  _add_map_x_67_m_clock = m_clock;
   assign  _add_map_x_66_moto_org_near = ((_net_5267)?data_in_org174:10'b0)|
    ((_net_1275)?data_in_org173:10'b0);
   assign  _add_map_x_66_moto_org_near1 = ((_net_5266)?data_in_org172:10'b0)|
    ((_net_1274)?data_in_org175:10'b0);
   assign  _add_map_x_66_moto_org_near2 = ((_net_5265)?data_in_org141:10'b0)|
    ((_net_1273)?data_in_org142:10'b0);
   assign  _add_map_x_66_moto_org_near3 = ((_net_5264)?data_in_org205:10'b0)|
    ((_net_1272)?data_in_org206:10'b0);
   assign  _add_map_x_66_moto_org = ((_net_5263)?data_in_org173:10'b0)|
    ((_net_1271)?data_in_org174:10'b0);
   assign  _add_map_x_66_sg_up = ((_net_5262)?sg_in174:2'b0)|
    ((_net_1270)?sg_in173:2'b0);
   assign  _add_map_x_66_sg_down = ((_net_5261)?sg_in141:2'b0)|
    ((_net_1269)?sg_in175:2'b0);
   assign  _add_map_x_66_sg_left = ((_net_5259)?sg_in205:2'b0)|
    ((_net_1267)?sg_in206:2'b0);
   assign  _add_map_x_66_sg_right = ((_net_5260)?sg_in172:2'b0)|
    ((_net_1268)?sg_in142:2'b0);
   assign  _add_map_x_66_wall_t_in = dig_w;
   assign  _add_map_x_66_moto = ((_net_5257)?data_in173:10'b0)|
    ((_net_1265)?data_in174:10'b0);
   assign  _add_map_x_66_up = ((_net_5256)?data_in174:10'b0)|
    ((_net_1264)?data_in173:10'b0);
   assign  _add_map_x_66_right = ((_net_5255)?data_in172:10'b0)|
    ((_net_1263)?data_in175:10'b0);
   assign  _add_map_x_66_down = ((_net_5254)?data_in141:10'b0)|
    ((_net_1262)?data_in142:10'b0);
   assign  _add_map_x_66_left = ((_net_5253)?data_in205:10'b0)|
    ((_net_1261)?data_in206:10'b0);
   assign  _add_map_x_66_start = start;
   assign  _add_map_x_66_goal = goal;
   assign  _add_map_x_66_now = ((_net_5250)?10'b0010101101:10'b0)|
    ((_net_1258)?10'b0010101110:10'b0);
   assign  _add_map_x_66_add_exe = (_net_5249|_net_1257);
   assign  _add_map_x_66_p_reset = p_reset;
   assign  _add_map_x_66_m_clock = m_clock;
   assign  _add_map_x_65_moto_org_near = ((_net_5248)?data_in_org172:10'b0)|
    ((_net_1256)?data_in_org171:10'b0);
   assign  _add_map_x_65_moto_org_near1 = ((_net_5247)?data_in_org170:10'b0)|
    ((_net_1255)?data_in_org173:10'b0);
   assign  _add_map_x_65_moto_org_near2 = ((_net_5246)?data_in_org139:10'b0)|
    ((_net_1254)?data_in_org140:10'b0);
   assign  _add_map_x_65_moto_org_near3 = ((_net_5245)?data_in_org203:10'b0)|
    ((_net_1253)?data_in_org204:10'b0);
   assign  _add_map_x_65_moto_org = ((_net_5244)?data_in_org171:10'b0)|
    ((_net_1252)?data_in_org172:10'b0);
   assign  _add_map_x_65_sg_up = ((_net_5243)?sg_in172:2'b0)|
    ((_net_1251)?sg_in171:2'b0);
   assign  _add_map_x_65_sg_down = ((_net_5242)?sg_in139:2'b0)|
    ((_net_1250)?sg_in173:2'b0);
   assign  _add_map_x_65_sg_left = ((_net_5240)?sg_in203:2'b0)|
    ((_net_1248)?sg_in204:2'b0);
   assign  _add_map_x_65_sg_right = ((_net_5241)?sg_in170:2'b0)|
    ((_net_1249)?sg_in140:2'b0);
   assign  _add_map_x_65_wall_t_in = dig_w;
   assign  _add_map_x_65_moto = ((_net_5238)?data_in171:10'b0)|
    ((_net_1246)?data_in172:10'b0);
   assign  _add_map_x_65_up = ((_net_5237)?data_in172:10'b0)|
    ((_net_1245)?data_in171:10'b0);
   assign  _add_map_x_65_right = ((_net_5236)?data_in170:10'b0)|
    ((_net_1244)?data_in173:10'b0);
   assign  _add_map_x_65_down = ((_net_5235)?data_in139:10'b0)|
    ((_net_1243)?data_in140:10'b0);
   assign  _add_map_x_65_left = ((_net_5234)?data_in203:10'b0)|
    ((_net_1242)?data_in204:10'b0);
   assign  _add_map_x_65_start = start;
   assign  _add_map_x_65_goal = goal;
   assign  _add_map_x_65_now = ((_net_5231)?10'b0010101011:10'b0)|
    ((_net_1239)?10'b0010101100:10'b0);
   assign  _add_map_x_65_add_exe = (_net_5230|_net_1238);
   assign  _add_map_x_65_p_reset = p_reset;
   assign  _add_map_x_65_m_clock = m_clock;
   assign  _add_map_x_64_moto_org_near = ((_net_5229)?data_in_org170:10'b0)|
    ((_net_1237)?data_in_org169:10'b0);
   assign  _add_map_x_64_moto_org_near1 = ((_net_5228)?data_in_org168:10'b0)|
    ((_net_1236)?data_in_org171:10'b0);
   assign  _add_map_x_64_moto_org_near2 = ((_net_5227)?data_in_org137:10'b0)|
    ((_net_1235)?data_in_org138:10'b0);
   assign  _add_map_x_64_moto_org_near3 = ((_net_5226)?data_in_org201:10'b0)|
    ((_net_1234)?data_in_org202:10'b0);
   assign  _add_map_x_64_moto_org = ((_net_5225)?data_in_org169:10'b0)|
    ((_net_1233)?data_in_org170:10'b0);
   assign  _add_map_x_64_sg_up = ((_net_5224)?sg_in170:2'b0)|
    ((_net_1232)?sg_in169:2'b0);
   assign  _add_map_x_64_sg_down = ((_net_5223)?sg_in137:2'b0)|
    ((_net_1231)?sg_in171:2'b0);
   assign  _add_map_x_64_sg_left = ((_net_5221)?sg_in201:2'b0)|
    ((_net_1229)?sg_in202:2'b0);
   assign  _add_map_x_64_sg_right = ((_net_5222)?sg_in168:2'b0)|
    ((_net_1230)?sg_in138:2'b0);
   assign  _add_map_x_64_wall_t_in = dig_w;
   assign  _add_map_x_64_moto = ((_net_5219)?data_in169:10'b0)|
    ((_net_1227)?data_in170:10'b0);
   assign  _add_map_x_64_up = ((_net_5218)?data_in170:10'b0)|
    ((_net_1226)?data_in169:10'b0);
   assign  _add_map_x_64_right = ((_net_5217)?data_in168:10'b0)|
    ((_net_1225)?data_in171:10'b0);
   assign  _add_map_x_64_down = ((_net_5216)?data_in137:10'b0)|
    ((_net_1224)?data_in138:10'b0);
   assign  _add_map_x_64_left = ((_net_5215)?data_in201:10'b0)|
    ((_net_1223)?data_in202:10'b0);
   assign  _add_map_x_64_start = start;
   assign  _add_map_x_64_goal = goal;
   assign  _add_map_x_64_now = ((_net_5212)?10'b0010101001:10'b0)|
    ((_net_1220)?10'b0010101010:10'b0);
   assign  _add_map_x_64_add_exe = (_net_5211|_net_1219);
   assign  _add_map_x_64_p_reset = p_reset;
   assign  _add_map_x_64_m_clock = m_clock;
   assign  _add_map_x_63_moto_org_near = ((_net_5210)?data_in_org168:10'b0)|
    ((_net_1218)?data_in_org167:10'b0);
   assign  _add_map_x_63_moto_org_near1 = ((_net_5209)?data_in_org166:10'b0)|
    ((_net_1217)?data_in_org169:10'b0);
   assign  _add_map_x_63_moto_org_near2 = ((_net_5208)?data_in_org135:10'b0)|
    ((_net_1216)?data_in_org136:10'b0);
   assign  _add_map_x_63_moto_org_near3 = ((_net_5207)?data_in_org199:10'b0)|
    ((_net_1215)?data_in_org200:10'b0);
   assign  _add_map_x_63_moto_org = ((_net_5206)?data_in_org167:10'b0)|
    ((_net_1214)?data_in_org168:10'b0);
   assign  _add_map_x_63_sg_up = ((_net_5205)?sg_in168:2'b0)|
    ((_net_1213)?sg_in167:2'b0);
   assign  _add_map_x_63_sg_down = ((_net_5204)?sg_in135:2'b0)|
    ((_net_1212)?sg_in169:2'b0);
   assign  _add_map_x_63_sg_left = ((_net_5202)?sg_in199:2'b0)|
    ((_net_1210)?sg_in200:2'b0);
   assign  _add_map_x_63_sg_right = ((_net_5203)?sg_in166:2'b0)|
    ((_net_1211)?sg_in136:2'b0);
   assign  _add_map_x_63_wall_t_in = dig_w;
   assign  _add_map_x_63_moto = ((_net_5200)?data_in167:10'b0)|
    ((_net_1208)?data_in168:10'b0);
   assign  _add_map_x_63_up = ((_net_5199)?data_in168:10'b0)|
    ((_net_1207)?data_in167:10'b0);
   assign  _add_map_x_63_right = ((_net_5198)?data_in166:10'b0)|
    ((_net_1206)?data_in169:10'b0);
   assign  _add_map_x_63_down = ((_net_5197)?data_in135:10'b0)|
    ((_net_1205)?data_in136:10'b0);
   assign  _add_map_x_63_left = ((_net_5196)?data_in199:10'b0)|
    ((_net_1204)?data_in200:10'b0);
   assign  _add_map_x_63_start = start;
   assign  _add_map_x_63_goal = goal;
   assign  _add_map_x_63_now = ((_net_5193)?10'b0010100111:10'b0)|
    ((_net_1201)?10'b0010101000:10'b0);
   assign  _add_map_x_63_add_exe = (_net_5192|_net_1200);
   assign  _add_map_x_63_p_reset = p_reset;
   assign  _add_map_x_63_m_clock = m_clock;
   assign  _add_map_x_62_moto_org_near = ((_net_5191)?data_in_org166:10'b0)|
    ((_net_1199)?data_in_org165:10'b0);
   assign  _add_map_x_62_moto_org_near1 = ((_net_5190)?data_in_org164:10'b0)|
    ((_net_1198)?data_in_org167:10'b0);
   assign  _add_map_x_62_moto_org_near2 = ((_net_5189)?data_in_org133:10'b0)|
    ((_net_1197)?data_in_org134:10'b0);
   assign  _add_map_x_62_moto_org_near3 = ((_net_5188)?data_in_org197:10'b0)|
    ((_net_1196)?data_in_org198:10'b0);
   assign  _add_map_x_62_moto_org = ((_net_5187)?data_in_org165:10'b0)|
    ((_net_1195)?data_in_org166:10'b0);
   assign  _add_map_x_62_sg_up = ((_net_5186)?sg_in166:2'b0)|
    ((_net_1194)?sg_in165:2'b0);
   assign  _add_map_x_62_sg_down = ((_net_5185)?sg_in133:2'b0)|
    ((_net_1193)?sg_in167:2'b0);
   assign  _add_map_x_62_sg_left = ((_net_5183)?sg_in197:2'b0)|
    ((_net_1191)?sg_in198:2'b0);
   assign  _add_map_x_62_sg_right = ((_net_5184)?sg_in164:2'b0)|
    ((_net_1192)?sg_in134:2'b0);
   assign  _add_map_x_62_wall_t_in = dig_w;
   assign  _add_map_x_62_moto = ((_net_5181)?data_in165:10'b0)|
    ((_net_1189)?data_in166:10'b0);
   assign  _add_map_x_62_up = ((_net_5180)?data_in166:10'b0)|
    ((_net_1188)?data_in165:10'b0);
   assign  _add_map_x_62_right = ((_net_5179)?data_in164:10'b0)|
    ((_net_1187)?data_in167:10'b0);
   assign  _add_map_x_62_down = ((_net_5178)?data_in133:10'b0)|
    ((_net_1186)?data_in134:10'b0);
   assign  _add_map_x_62_left = ((_net_5177)?data_in197:10'b0)|
    ((_net_1185)?data_in198:10'b0);
   assign  _add_map_x_62_start = start;
   assign  _add_map_x_62_goal = goal;
   assign  _add_map_x_62_now = ((_net_5174)?10'b0010100101:10'b0)|
    ((_net_1182)?10'b0010100110:10'b0);
   assign  _add_map_x_62_add_exe = (_net_5173|_net_1181);
   assign  _add_map_x_62_p_reset = p_reset;
   assign  _add_map_x_62_m_clock = m_clock;
   assign  _add_map_x_61_moto_org_near = ((_net_5172)?data_in_org164:10'b0)|
    ((_net_1180)?data_in_org163:10'b0);
   assign  _add_map_x_61_moto_org_near1 = ((_net_5171)?data_in_org162:10'b0)|
    ((_net_1179)?data_in_org165:10'b0);
   assign  _add_map_x_61_moto_org_near2 = ((_net_5170)?data_in_org131:10'b0)|
    ((_net_1178)?data_in_org132:10'b0);
   assign  _add_map_x_61_moto_org_near3 = ((_net_5169)?data_in_org195:10'b0)|
    ((_net_1177)?data_in_org196:10'b0);
   assign  _add_map_x_61_moto_org = ((_net_5168)?data_in_org163:10'b0)|
    ((_net_1176)?data_in_org164:10'b0);
   assign  _add_map_x_61_sg_up = ((_net_5167)?sg_in164:2'b0)|
    ((_net_1175)?sg_in163:2'b0);
   assign  _add_map_x_61_sg_down = ((_net_5166)?sg_in131:2'b0)|
    ((_net_1174)?sg_in165:2'b0);
   assign  _add_map_x_61_sg_left = ((_net_5164)?sg_in195:2'b0)|
    ((_net_1172)?sg_in196:2'b0);
   assign  _add_map_x_61_sg_right = ((_net_5165)?sg_in162:2'b0)|
    ((_net_1173)?sg_in132:2'b0);
   assign  _add_map_x_61_wall_t_in = dig_w;
   assign  _add_map_x_61_moto = ((_net_5162)?data_in163:10'b0)|
    ((_net_1170)?data_in164:10'b0);
   assign  _add_map_x_61_up = ((_net_5161)?data_in164:10'b0)|
    ((_net_1169)?data_in163:10'b0);
   assign  _add_map_x_61_right = ((_net_5160)?data_in162:10'b0)|
    ((_net_1168)?data_in165:10'b0);
   assign  _add_map_x_61_down = ((_net_5159)?data_in131:10'b0)|
    ((_net_1167)?data_in132:10'b0);
   assign  _add_map_x_61_left = ((_net_5158)?data_in195:10'b0)|
    ((_net_1166)?data_in196:10'b0);
   assign  _add_map_x_61_start = start;
   assign  _add_map_x_61_goal = goal;
   assign  _add_map_x_61_now = ((_net_5155)?10'b0010100011:10'b0)|
    ((_net_1163)?10'b0010100100:10'b0);
   assign  _add_map_x_61_add_exe = (_net_5154|_net_1162);
   assign  _add_map_x_61_p_reset = p_reset;
   assign  _add_map_x_61_m_clock = m_clock;
   assign  _add_map_x_60_moto_org_near = ((_net_5153)?data_in_org162:10'b0)|
    ((_net_1161)?data_in_org161:10'b0);
   assign  _add_map_x_60_moto_org_near1 = ((_net_5152)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1160)?data_in_org163:10'b0);
   assign  _add_map_x_60_moto_org_near2 = ((_net_5151)?data_in_org129:10'b0)|
    ((_net_1159)?data_in_org130:10'b0);
   assign  _add_map_x_60_moto_org_near3 = ((_net_5150)?data_in_org193:10'b0)|
    ((_net_1158)?data_in_org194:10'b0);
   assign  _add_map_x_60_moto_org = ((_net_5149)?data_in_org161:10'b0)|
    ((_net_1157)?data_in_org162:10'b0);
   assign  _add_map_x_60_sg_up = ((_net_5148)?sg_in162:2'b0)|
    ((_net_1156)?sg_in161:2'b0);
   assign  _add_map_x_60_sg_down = ((_net_5147)?sg_in129:2'b0)|
    ((_net_1155)?sg_in163:2'b0);
   assign  _add_map_x_60_sg_left = ((_net_5145)?sg_in193:2'b0)|
    ((_net_1153)?sg_in194:2'b0);
   assign  _add_map_x_60_sg_right = ((_net_5146)?3'b000:2'b0)|
    ((_net_1154)?sg_in130:2'b0);
   assign  _add_map_x_60_wall_t_in = dig_w;
   assign  _add_map_x_60_moto = ((_net_5143)?data_in161:10'b0)|
    ((_net_1151)?data_in162:10'b0);
   assign  _add_map_x_60_up = ((_net_5142)?data_in162:10'b0)|
    ((_net_1150)?data_in161:10'b0);
   assign  _add_map_x_60_right = ((_net_5141)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1149)?data_in163:10'b0);
   assign  _add_map_x_60_down = ((_net_5140)?data_in129:10'b0)|
    ((_net_1148)?data_in130:10'b0);
   assign  _add_map_x_60_left = ((_net_5139)?data_in193:10'b0)|
    ((_net_1147)?data_in194:10'b0);
   assign  _add_map_x_60_start = start;
   assign  _add_map_x_60_goal = goal;
   assign  _add_map_x_60_now = ((_net_5136)?10'b0010100001:10'b0)|
    ((_net_1144)?10'b0010100010:10'b0);
   assign  _add_map_x_60_add_exe = (_net_5135|_net_1143);
   assign  _add_map_x_60_p_reset = p_reset;
   assign  _add_map_x_60_m_clock = m_clock;
   assign  _add_map_x_59_moto_org_near = ((_net_5134)?data_in_org157:10'b0)|
    ((_net_1142)?data_in_org158:10'b0);
   assign  _add_map_x_59_moto_org_near1 = ((_net_5133)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1141)?data_in_org156:10'b0);
   assign  _add_map_x_59_moto_org_near2 = ((_net_5132)?data_in_org126:10'b0)|
    ((_net_1140)?data_in_org125:10'b0);
   assign  _add_map_x_59_moto_org_near3 = ((_net_5131)?data_in_org190:10'b0)|
    ((_net_1139)?data_in_org189:10'b0);
   assign  _add_map_x_59_moto_org = ((_net_5130)?data_in_org158:10'b0)|
    ((_net_1138)?data_in_org157:10'b0);
   assign  _add_map_x_59_sg_up = ((_net_5129)?sg_in157:2'b0)|
    ((_net_1137)?sg_in158:2'b0);
   assign  _add_map_x_59_sg_down = ((_net_5128)?3'b000:2'b0)|
    ((_net_1136)?sg_in156:2'b0);
   assign  _add_map_x_59_sg_left = ((_net_5126)?sg_in190:2'b0)|
    ((_net_1134)?sg_in189:2'b0);
   assign  _add_map_x_59_sg_right = ((_net_5127)?sg_in126:2'b0)|
    ((_net_1135)?sg_in125:2'b0);
   assign  _add_map_x_59_wall_t_in = dig_w;
   assign  _add_map_x_59_moto = ((_net_5124)?data_in158:10'b0)|
    ((_net_1132)?data_in157:10'b0);
   assign  _add_map_x_59_up = ((_net_5123)?data_in157:10'b0)|
    ((_net_1131)?data_in158:10'b0);
   assign  _add_map_x_59_right = ((_net_5122)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_1130)?data_in156:10'b0);
   assign  _add_map_x_59_down = ((_net_5121)?data_in126:10'b0)|
    ((_net_1129)?data_in125:10'b0);
   assign  _add_map_x_59_left = ((_net_5120)?data_in190:10'b0)|
    ((_net_1128)?data_in189:10'b0);
   assign  _add_map_x_59_start = start;
   assign  _add_map_x_59_goal = goal;
   assign  _add_map_x_59_now = ((_net_5117)?10'b0010011110:10'b0)|
    ((_net_1125)?10'b0010011101:10'b0);
   assign  _add_map_x_59_add_exe = (_net_5116|_net_1124);
   assign  _add_map_x_59_p_reset = p_reset;
   assign  _add_map_x_59_m_clock = m_clock;
   assign  _add_map_x_58_moto_org_near = ((_net_5115)?data_in_org155:10'b0)|
    ((_net_1123)?data_in_org156:10'b0);
   assign  _add_map_x_58_moto_org_near1 = ((_net_5114)?data_in_org157:10'b0)|
    ((_net_1122)?data_in_org154:10'b0);
   assign  _add_map_x_58_moto_org_near2 = ((_net_5113)?data_in_org124:10'b0)|
    ((_net_1121)?data_in_org123:10'b0);
   assign  _add_map_x_58_moto_org_near3 = ((_net_5112)?data_in_org188:10'b0)|
    ((_net_1120)?data_in_org187:10'b0);
   assign  _add_map_x_58_moto_org = ((_net_5111)?data_in_org156:10'b0)|
    ((_net_1119)?data_in_org155:10'b0);
   assign  _add_map_x_58_sg_up = ((_net_5110)?sg_in155:2'b0)|
    ((_net_1118)?sg_in156:2'b0);
   assign  _add_map_x_58_sg_down = ((_net_5109)?sg_in157:2'b0)|
    ((_net_1117)?sg_in154:2'b0);
   assign  _add_map_x_58_sg_left = ((_net_5107)?sg_in188:2'b0)|
    ((_net_1115)?sg_in187:2'b0);
   assign  _add_map_x_58_sg_right = ((_net_5108)?sg_in124:2'b0)|
    ((_net_1116)?sg_in123:2'b0);
   assign  _add_map_x_58_wall_t_in = dig_w;
   assign  _add_map_x_58_moto = ((_net_5105)?data_in156:10'b0)|
    ((_net_1113)?data_in155:10'b0);
   assign  _add_map_x_58_up = ((_net_5104)?data_in155:10'b0)|
    ((_net_1112)?data_in156:10'b0);
   assign  _add_map_x_58_right = ((_net_5103)?data_in157:10'b0)|
    ((_net_1111)?data_in154:10'b0);
   assign  _add_map_x_58_down = ((_net_5102)?data_in124:10'b0)|
    ((_net_1110)?data_in123:10'b0);
   assign  _add_map_x_58_left = ((_net_5101)?data_in188:10'b0)|
    ((_net_1109)?data_in187:10'b0);
   assign  _add_map_x_58_start = start;
   assign  _add_map_x_58_goal = goal;
   assign  _add_map_x_58_now = ((_net_5098)?10'b0010011100:10'b0)|
    ((_net_1106)?10'b0010011011:10'b0);
   assign  _add_map_x_58_add_exe = (_net_5097|_net_1105);
   assign  _add_map_x_58_p_reset = p_reset;
   assign  _add_map_x_58_m_clock = m_clock;
   assign  _add_map_x_57_moto_org_near = ((_net_5096)?data_in_org153:10'b0)|
    ((_net_1104)?data_in_org154:10'b0);
   assign  _add_map_x_57_moto_org_near1 = ((_net_5095)?data_in_org155:10'b0)|
    ((_net_1103)?data_in_org152:10'b0);
   assign  _add_map_x_57_moto_org_near2 = ((_net_5094)?data_in_org122:10'b0)|
    ((_net_1102)?data_in_org121:10'b0);
   assign  _add_map_x_57_moto_org_near3 = ((_net_5093)?data_in_org186:10'b0)|
    ((_net_1101)?data_in_org185:10'b0);
   assign  _add_map_x_57_moto_org = ((_net_5092)?data_in_org154:10'b0)|
    ((_net_1100)?data_in_org153:10'b0);
   assign  _add_map_x_57_sg_up = ((_net_5091)?sg_in153:2'b0)|
    ((_net_1099)?sg_in154:2'b0);
   assign  _add_map_x_57_sg_down = ((_net_5090)?sg_in155:2'b0)|
    ((_net_1098)?sg_in152:2'b0);
   assign  _add_map_x_57_sg_left = ((_net_5088)?sg_in186:2'b0)|
    ((_net_1096)?sg_in185:2'b0);
   assign  _add_map_x_57_sg_right = ((_net_5089)?sg_in122:2'b0)|
    ((_net_1097)?sg_in121:2'b0);
   assign  _add_map_x_57_wall_t_in = dig_w;
   assign  _add_map_x_57_moto = ((_net_5086)?data_in154:10'b0)|
    ((_net_1094)?data_in153:10'b0);
   assign  _add_map_x_57_up = ((_net_5085)?data_in153:10'b0)|
    ((_net_1093)?data_in154:10'b0);
   assign  _add_map_x_57_right = ((_net_5084)?data_in155:10'b0)|
    ((_net_1092)?data_in152:10'b0);
   assign  _add_map_x_57_down = ((_net_5083)?data_in122:10'b0)|
    ((_net_1091)?data_in121:10'b0);
   assign  _add_map_x_57_left = ((_net_5082)?data_in186:10'b0)|
    ((_net_1090)?data_in185:10'b0);
   assign  _add_map_x_57_start = start;
   assign  _add_map_x_57_goal = goal;
   assign  _add_map_x_57_now = ((_net_5079)?10'b0010011010:10'b0)|
    ((_net_1087)?10'b0010011001:10'b0);
   assign  _add_map_x_57_add_exe = (_net_5078|_net_1086);
   assign  _add_map_x_57_p_reset = p_reset;
   assign  _add_map_x_57_m_clock = m_clock;
   assign  _add_map_x_56_moto_org_near = ((_net_5077)?data_in_org151:10'b0)|
    ((_net_1085)?data_in_org152:10'b0);
   assign  _add_map_x_56_moto_org_near1 = ((_net_5076)?data_in_org153:10'b0)|
    ((_net_1084)?data_in_org150:10'b0);
   assign  _add_map_x_56_moto_org_near2 = ((_net_5075)?data_in_org120:10'b0)|
    ((_net_1083)?data_in_org119:10'b0);
   assign  _add_map_x_56_moto_org_near3 = ((_net_5074)?data_in_org184:10'b0)|
    ((_net_1082)?data_in_org183:10'b0);
   assign  _add_map_x_56_moto_org = ((_net_5073)?data_in_org152:10'b0)|
    ((_net_1081)?data_in_org151:10'b0);
   assign  _add_map_x_56_sg_up = ((_net_5072)?sg_in151:2'b0)|
    ((_net_1080)?sg_in152:2'b0);
   assign  _add_map_x_56_sg_down = ((_net_5071)?sg_in153:2'b0)|
    ((_net_1079)?sg_in150:2'b0);
   assign  _add_map_x_56_sg_left = ((_net_5069)?sg_in184:2'b0)|
    ((_net_1077)?sg_in183:2'b0);
   assign  _add_map_x_56_sg_right = ((_net_5070)?sg_in120:2'b0)|
    ((_net_1078)?sg_in119:2'b0);
   assign  _add_map_x_56_wall_t_in = dig_w;
   assign  _add_map_x_56_moto = ((_net_5067)?data_in152:10'b0)|
    ((_net_1075)?data_in151:10'b0);
   assign  _add_map_x_56_up = ((_net_5066)?data_in151:10'b0)|
    ((_net_1074)?data_in152:10'b0);
   assign  _add_map_x_56_right = ((_net_5065)?data_in153:10'b0)|
    ((_net_1073)?data_in150:10'b0);
   assign  _add_map_x_56_down = ((_net_5064)?data_in120:10'b0)|
    ((_net_1072)?data_in119:10'b0);
   assign  _add_map_x_56_left = ((_net_5063)?data_in184:10'b0)|
    ((_net_1071)?data_in183:10'b0);
   assign  _add_map_x_56_start = start;
   assign  _add_map_x_56_goal = goal;
   assign  _add_map_x_56_now = ((_net_5060)?10'b0010011000:10'b0)|
    ((_net_1068)?10'b0010010111:10'b0);
   assign  _add_map_x_56_add_exe = (_net_5059|_net_1067);
   assign  _add_map_x_56_p_reset = p_reset;
   assign  _add_map_x_56_m_clock = m_clock;
   assign  _add_map_x_55_moto_org_near = ((_net_5058)?data_in_org149:10'b0)|
    ((_net_1066)?data_in_org150:10'b0);
   assign  _add_map_x_55_moto_org_near1 = ((_net_5057)?data_in_org151:10'b0)|
    ((_net_1065)?data_in_org148:10'b0);
   assign  _add_map_x_55_moto_org_near2 = ((_net_5056)?data_in_org118:10'b0)|
    ((_net_1064)?data_in_org117:10'b0);
   assign  _add_map_x_55_moto_org_near3 = ((_net_5055)?data_in_org182:10'b0)|
    ((_net_1063)?data_in_org181:10'b0);
   assign  _add_map_x_55_moto_org = ((_net_5054)?data_in_org150:10'b0)|
    ((_net_1062)?data_in_org149:10'b0);
   assign  _add_map_x_55_sg_up = ((_net_5053)?sg_in149:2'b0)|
    ((_net_1061)?sg_in150:2'b0);
   assign  _add_map_x_55_sg_down = ((_net_5052)?sg_in151:2'b0)|
    ((_net_1060)?sg_in148:2'b0);
   assign  _add_map_x_55_sg_left = ((_net_5050)?sg_in182:2'b0)|
    ((_net_1058)?sg_in181:2'b0);
   assign  _add_map_x_55_sg_right = ((_net_5051)?sg_in118:2'b0)|
    ((_net_1059)?sg_in117:2'b0);
   assign  _add_map_x_55_wall_t_in = dig_w;
   assign  _add_map_x_55_moto = ((_net_5048)?data_in150:10'b0)|
    ((_net_1056)?data_in149:10'b0);
   assign  _add_map_x_55_up = ((_net_5047)?data_in149:10'b0)|
    ((_net_1055)?data_in150:10'b0);
   assign  _add_map_x_55_right = ((_net_5046)?data_in151:10'b0)|
    ((_net_1054)?data_in148:10'b0);
   assign  _add_map_x_55_down = ((_net_5045)?data_in118:10'b0)|
    ((_net_1053)?data_in117:10'b0);
   assign  _add_map_x_55_left = ((_net_5044)?data_in182:10'b0)|
    ((_net_1052)?data_in181:10'b0);
   assign  _add_map_x_55_start = start;
   assign  _add_map_x_55_goal = goal;
   assign  _add_map_x_55_now = ((_net_5041)?10'b0010010110:10'b0)|
    ((_net_1049)?10'b0010010101:10'b0);
   assign  _add_map_x_55_add_exe = (_net_5040|_net_1048);
   assign  _add_map_x_55_p_reset = p_reset;
   assign  _add_map_x_55_m_clock = m_clock;
   assign  _add_map_x_54_moto_org_near = ((_net_5039)?data_in_org147:10'b0)|
    ((_net_1047)?data_in_org148:10'b0);
   assign  _add_map_x_54_moto_org_near1 = ((_net_5038)?data_in_org149:10'b0)|
    ((_net_1046)?data_in_org146:10'b0);
   assign  _add_map_x_54_moto_org_near2 = ((_net_5037)?data_in_org116:10'b0)|
    ((_net_1045)?data_in_org115:10'b0);
   assign  _add_map_x_54_moto_org_near3 = ((_net_5036)?data_in_org180:10'b0)|
    ((_net_1044)?data_in_org179:10'b0);
   assign  _add_map_x_54_moto_org = ((_net_5035)?data_in_org148:10'b0)|
    ((_net_1043)?data_in_org147:10'b0);
   assign  _add_map_x_54_sg_up = ((_net_5034)?sg_in147:2'b0)|
    ((_net_1042)?sg_in148:2'b0);
   assign  _add_map_x_54_sg_down = ((_net_5033)?sg_in149:2'b0)|
    ((_net_1041)?sg_in146:2'b0);
   assign  _add_map_x_54_sg_left = ((_net_5031)?sg_in180:2'b0)|
    ((_net_1039)?sg_in179:2'b0);
   assign  _add_map_x_54_sg_right = ((_net_5032)?sg_in116:2'b0)|
    ((_net_1040)?sg_in115:2'b0);
   assign  _add_map_x_54_wall_t_in = dig_w;
   assign  _add_map_x_54_moto = ((_net_5029)?data_in148:10'b0)|
    ((_net_1037)?data_in147:10'b0);
   assign  _add_map_x_54_up = ((_net_5028)?data_in147:10'b0)|
    ((_net_1036)?data_in148:10'b0);
   assign  _add_map_x_54_right = ((_net_5027)?data_in149:10'b0)|
    ((_net_1035)?data_in146:10'b0);
   assign  _add_map_x_54_down = ((_net_5026)?data_in116:10'b0)|
    ((_net_1034)?data_in115:10'b0);
   assign  _add_map_x_54_left = ((_net_5025)?data_in180:10'b0)|
    ((_net_1033)?data_in179:10'b0);
   assign  _add_map_x_54_start = start;
   assign  _add_map_x_54_goal = goal;
   assign  _add_map_x_54_now = ((_net_5022)?10'b0010010100:10'b0)|
    ((_net_1030)?10'b0010010011:10'b0);
   assign  _add_map_x_54_add_exe = (_net_5021|_net_1029);
   assign  _add_map_x_54_p_reset = p_reset;
   assign  _add_map_x_54_m_clock = m_clock;
   assign  _add_map_x_53_moto_org_near = ((_net_5020)?data_in_org145:10'b0)|
    ((_net_1028)?data_in_org146:10'b0);
   assign  _add_map_x_53_moto_org_near1 = ((_net_5019)?data_in_org147:10'b0)|
    ((_net_1027)?data_in_org144:10'b0);
   assign  _add_map_x_53_moto_org_near2 = ((_net_5018)?data_in_org114:10'b0)|
    ((_net_1026)?data_in_org113:10'b0);
   assign  _add_map_x_53_moto_org_near3 = ((_net_5017)?data_in_org178:10'b0)|
    ((_net_1025)?data_in_org177:10'b0);
   assign  _add_map_x_53_moto_org = ((_net_5016)?data_in_org146:10'b0)|
    ((_net_1024)?data_in_org145:10'b0);
   assign  _add_map_x_53_sg_up = ((_net_5015)?sg_in145:2'b0)|
    ((_net_1023)?sg_in146:2'b0);
   assign  _add_map_x_53_sg_down = ((_net_5014)?sg_in147:2'b0)|
    ((_net_1022)?sg_in144:2'b0);
   assign  _add_map_x_53_sg_left = ((_net_5012)?sg_in178:2'b0)|
    ((_net_1020)?sg_in177:2'b0);
   assign  _add_map_x_53_sg_right = ((_net_5013)?sg_in114:2'b0)|
    ((_net_1021)?sg_in113:2'b0);
   assign  _add_map_x_53_wall_t_in = dig_w;
   assign  _add_map_x_53_moto = ((_net_5010)?data_in146:10'b0)|
    ((_net_1018)?data_in145:10'b0);
   assign  _add_map_x_53_up = ((_net_5009)?data_in145:10'b0)|
    ((_net_1017)?data_in146:10'b0);
   assign  _add_map_x_53_right = ((_net_5008)?data_in147:10'b0)|
    ((_net_1016)?data_in144:10'b0);
   assign  _add_map_x_53_down = ((_net_5007)?data_in114:10'b0)|
    ((_net_1015)?data_in113:10'b0);
   assign  _add_map_x_53_left = ((_net_5006)?data_in178:10'b0)|
    ((_net_1014)?data_in177:10'b0);
   assign  _add_map_x_53_start = start;
   assign  _add_map_x_53_goal = goal;
   assign  _add_map_x_53_now = ((_net_5003)?10'b0010010010:10'b0)|
    ((_net_1011)?10'b0010010001:10'b0);
   assign  _add_map_x_53_add_exe = (_net_5002|_net_1010);
   assign  _add_map_x_53_p_reset = p_reset;
   assign  _add_map_x_53_m_clock = m_clock;
   assign  _add_map_x_52_moto_org_near = ((_net_5001)?data_in_org143:10'b0)|
    ((_net_1009)?data_in_org144:10'b0);
   assign  _add_map_x_52_moto_org_near1 = ((_net_5000)?data_in_org145:10'b0)|
    ((_net_1008)?data_in_org142:10'b0);
   assign  _add_map_x_52_moto_org_near2 = ((_net_4999)?data_in_org112:10'b0)|
    ((_net_1007)?data_in_org111:10'b0);
   assign  _add_map_x_52_moto_org_near3 = ((_net_4998)?data_in_org176:10'b0)|
    ((_net_1006)?data_in_org175:10'b0);
   assign  _add_map_x_52_moto_org = ((_net_4997)?data_in_org144:10'b0)|
    ((_net_1005)?data_in_org143:10'b0);
   assign  _add_map_x_52_sg_up = ((_net_4996)?sg_in143:2'b0)|
    ((_net_1004)?sg_in144:2'b0);
   assign  _add_map_x_52_sg_down = ((_net_4995)?sg_in145:2'b0)|
    ((_net_1003)?sg_in142:2'b0);
   assign  _add_map_x_52_sg_left = ((_net_4993)?sg_in176:2'b0)|
    ((_net_1001)?sg_in175:2'b0);
   assign  _add_map_x_52_sg_right = ((_net_4994)?sg_in112:2'b0)|
    ((_net_1002)?sg_in111:2'b0);
   assign  _add_map_x_52_wall_t_in = dig_w;
   assign  _add_map_x_52_moto = ((_net_4991)?data_in144:10'b0)|
    ((_net_999)?data_in143:10'b0);
   assign  _add_map_x_52_up = ((_net_4990)?data_in143:10'b0)|
    ((_net_998)?data_in144:10'b0);
   assign  _add_map_x_52_right = ((_net_4989)?data_in145:10'b0)|
    ((_net_997)?data_in142:10'b0);
   assign  _add_map_x_52_down = ((_net_4988)?data_in112:10'b0)|
    ((_net_996)?data_in111:10'b0);
   assign  _add_map_x_52_left = ((_net_4987)?data_in176:10'b0)|
    ((_net_995)?data_in175:10'b0);
   assign  _add_map_x_52_start = start;
   assign  _add_map_x_52_goal = goal;
   assign  _add_map_x_52_now = ((_net_4984)?10'b0010010000:10'b0)|
    ((_net_992)?10'b0010001111:10'b0);
   assign  _add_map_x_52_add_exe = (_net_4983|_net_991);
   assign  _add_map_x_52_p_reset = p_reset;
   assign  _add_map_x_52_m_clock = m_clock;
   assign  _add_map_x_51_moto_org_near = ((_net_4982)?data_in_org141:10'b0)|
    ((_net_990)?data_in_org142:10'b0);
   assign  _add_map_x_51_moto_org_near1 = ((_net_4981)?data_in_org143:10'b0)|
    ((_net_989)?data_in_org140:10'b0);
   assign  _add_map_x_51_moto_org_near2 = ((_net_4980)?data_in_org110:10'b0)|
    ((_net_988)?data_in_org109:10'b0);
   assign  _add_map_x_51_moto_org_near3 = ((_net_4979)?data_in_org174:10'b0)|
    ((_net_987)?data_in_org173:10'b0);
   assign  _add_map_x_51_moto_org = ((_net_4978)?data_in_org142:10'b0)|
    ((_net_986)?data_in_org141:10'b0);
   assign  _add_map_x_51_sg_up = ((_net_4977)?sg_in141:2'b0)|
    ((_net_985)?sg_in142:2'b0);
   assign  _add_map_x_51_sg_down = ((_net_4976)?sg_in143:2'b0)|
    ((_net_984)?sg_in140:2'b0);
   assign  _add_map_x_51_sg_left = ((_net_4974)?sg_in174:2'b0)|
    ((_net_982)?sg_in173:2'b0);
   assign  _add_map_x_51_sg_right = ((_net_4975)?sg_in110:2'b0)|
    ((_net_983)?sg_in109:2'b0);
   assign  _add_map_x_51_wall_t_in = dig_w;
   assign  _add_map_x_51_moto = ((_net_4972)?data_in142:10'b0)|
    ((_net_980)?data_in141:10'b0);
   assign  _add_map_x_51_up = ((_net_4971)?data_in141:10'b0)|
    ((_net_979)?data_in142:10'b0);
   assign  _add_map_x_51_right = ((_net_4970)?data_in143:10'b0)|
    ((_net_978)?data_in140:10'b0);
   assign  _add_map_x_51_down = ((_net_4969)?data_in110:10'b0)|
    ((_net_977)?data_in109:10'b0);
   assign  _add_map_x_51_left = ((_net_4968)?data_in174:10'b0)|
    ((_net_976)?data_in173:10'b0);
   assign  _add_map_x_51_start = start;
   assign  _add_map_x_51_goal = goal;
   assign  _add_map_x_51_now = ((_net_4965)?10'b0010001110:10'b0)|
    ((_net_973)?10'b0010001101:10'b0);
   assign  _add_map_x_51_add_exe = (_net_4964|_net_972);
   assign  _add_map_x_51_p_reset = p_reset;
   assign  _add_map_x_51_m_clock = m_clock;
   assign  _add_map_x_50_moto_org_near = ((_net_4963)?data_in_org139:10'b0)|
    ((_net_971)?data_in_org140:10'b0);
   assign  _add_map_x_50_moto_org_near1 = ((_net_4962)?data_in_org141:10'b0)|
    ((_net_970)?data_in_org138:10'b0);
   assign  _add_map_x_50_moto_org_near2 = ((_net_4961)?data_in_org108:10'b0)|
    ((_net_969)?data_in_org107:10'b0);
   assign  _add_map_x_50_moto_org_near3 = ((_net_4960)?data_in_org172:10'b0)|
    ((_net_968)?data_in_org171:10'b0);
   assign  _add_map_x_50_moto_org = ((_net_4959)?data_in_org140:10'b0)|
    ((_net_967)?data_in_org139:10'b0);
   assign  _add_map_x_50_sg_up = ((_net_4958)?sg_in139:2'b0)|
    ((_net_966)?sg_in140:2'b0);
   assign  _add_map_x_50_sg_down = ((_net_4957)?sg_in141:2'b0)|
    ((_net_965)?sg_in138:2'b0);
   assign  _add_map_x_50_sg_left = ((_net_4955)?sg_in172:2'b0)|
    ((_net_963)?sg_in171:2'b0);
   assign  _add_map_x_50_sg_right = ((_net_4956)?sg_in108:2'b0)|
    ((_net_964)?sg_in107:2'b0);
   assign  _add_map_x_50_wall_t_in = dig_w;
   assign  _add_map_x_50_moto = ((_net_4953)?data_in140:10'b0)|
    ((_net_961)?data_in139:10'b0);
   assign  _add_map_x_50_up = ((_net_4952)?data_in139:10'b0)|
    ((_net_960)?data_in140:10'b0);
   assign  _add_map_x_50_right = ((_net_4951)?data_in141:10'b0)|
    ((_net_959)?data_in138:10'b0);
   assign  _add_map_x_50_down = ((_net_4950)?data_in108:10'b0)|
    ((_net_958)?data_in107:10'b0);
   assign  _add_map_x_50_left = ((_net_4949)?data_in172:10'b0)|
    ((_net_957)?data_in171:10'b0);
   assign  _add_map_x_50_start = start;
   assign  _add_map_x_50_goal = goal;
   assign  _add_map_x_50_now = ((_net_4946)?10'b0010001100:10'b0)|
    ((_net_954)?10'b0010001011:10'b0);
   assign  _add_map_x_50_add_exe = (_net_4945|_net_953);
   assign  _add_map_x_50_p_reset = p_reset;
   assign  _add_map_x_50_m_clock = m_clock;
   assign  _add_map_x_49_moto_org_near = ((_net_4944)?data_in_org137:10'b0)|
    ((_net_952)?data_in_org138:10'b0);
   assign  _add_map_x_49_moto_org_near1 = ((_net_4943)?data_in_org139:10'b0)|
    ((_net_951)?data_in_org136:10'b0);
   assign  _add_map_x_49_moto_org_near2 = ((_net_4942)?data_in_org106:10'b0)|
    ((_net_950)?data_in_org105:10'b0);
   assign  _add_map_x_49_moto_org_near3 = ((_net_4941)?data_in_org170:10'b0)|
    ((_net_949)?data_in_org169:10'b0);
   assign  _add_map_x_49_moto_org = ((_net_4940)?data_in_org138:10'b0)|
    ((_net_948)?data_in_org137:10'b0);
   assign  _add_map_x_49_sg_up = ((_net_4939)?sg_in137:2'b0)|
    ((_net_947)?sg_in138:2'b0);
   assign  _add_map_x_49_sg_down = ((_net_4938)?sg_in139:2'b0)|
    ((_net_946)?sg_in136:2'b0);
   assign  _add_map_x_49_sg_left = ((_net_4936)?sg_in170:2'b0)|
    ((_net_944)?sg_in169:2'b0);
   assign  _add_map_x_49_sg_right = ((_net_4937)?sg_in106:2'b0)|
    ((_net_945)?sg_in105:2'b0);
   assign  _add_map_x_49_wall_t_in = dig_w;
   assign  _add_map_x_49_moto = ((_net_4934)?data_in138:10'b0)|
    ((_net_942)?data_in137:10'b0);
   assign  _add_map_x_49_up = ((_net_4933)?data_in137:10'b0)|
    ((_net_941)?data_in138:10'b0);
   assign  _add_map_x_49_right = ((_net_4932)?data_in139:10'b0)|
    ((_net_940)?data_in136:10'b0);
   assign  _add_map_x_49_down = ((_net_4931)?data_in106:10'b0)|
    ((_net_939)?data_in105:10'b0);
   assign  _add_map_x_49_left = ((_net_4930)?data_in170:10'b0)|
    ((_net_938)?data_in169:10'b0);
   assign  _add_map_x_49_start = start;
   assign  _add_map_x_49_goal = goal;
   assign  _add_map_x_49_now = ((_net_4927)?10'b0010001010:10'b0)|
    ((_net_935)?10'b0010001001:10'b0);
   assign  _add_map_x_49_add_exe = (_net_4926|_net_934);
   assign  _add_map_x_49_p_reset = p_reset;
   assign  _add_map_x_49_m_clock = m_clock;
   assign  _add_map_x_48_moto_org_near = ((_net_4925)?data_in_org135:10'b0)|
    ((_net_933)?data_in_org136:10'b0);
   assign  _add_map_x_48_moto_org_near1 = ((_net_4924)?data_in_org137:10'b0)|
    ((_net_932)?data_in_org134:10'b0);
   assign  _add_map_x_48_moto_org_near2 = ((_net_4923)?data_in_org104:10'b0)|
    ((_net_931)?data_in_org103:10'b0);
   assign  _add_map_x_48_moto_org_near3 = ((_net_4922)?data_in_org168:10'b0)|
    ((_net_930)?data_in_org167:10'b0);
   assign  _add_map_x_48_moto_org = ((_net_4921)?data_in_org136:10'b0)|
    ((_net_929)?data_in_org135:10'b0);
   assign  _add_map_x_48_sg_up = ((_net_4920)?sg_in135:2'b0)|
    ((_net_928)?sg_in136:2'b0);
   assign  _add_map_x_48_sg_down = ((_net_4919)?sg_in137:2'b0)|
    ((_net_927)?sg_in134:2'b0);
   assign  _add_map_x_48_sg_left = ((_net_4917)?sg_in168:2'b0)|
    ((_net_925)?sg_in167:2'b0);
   assign  _add_map_x_48_sg_right = ((_net_4918)?sg_in104:2'b0)|
    ((_net_926)?sg_in103:2'b0);
   assign  _add_map_x_48_wall_t_in = dig_w;
   assign  _add_map_x_48_moto = ((_net_4915)?data_in136:10'b0)|
    ((_net_923)?data_in135:10'b0);
   assign  _add_map_x_48_up = ((_net_4914)?data_in135:10'b0)|
    ((_net_922)?data_in136:10'b0);
   assign  _add_map_x_48_right = ((_net_4913)?data_in137:10'b0)|
    ((_net_921)?data_in134:10'b0);
   assign  _add_map_x_48_down = ((_net_4912)?data_in104:10'b0)|
    ((_net_920)?data_in103:10'b0);
   assign  _add_map_x_48_left = ((_net_4911)?data_in168:10'b0)|
    ((_net_919)?data_in167:10'b0);
   assign  _add_map_x_48_start = start;
   assign  _add_map_x_48_goal = goal;
   assign  _add_map_x_48_now = ((_net_4908)?10'b0010001000:10'b0)|
    ((_net_916)?10'b0010000111:10'b0);
   assign  _add_map_x_48_add_exe = (_net_4907|_net_915);
   assign  _add_map_x_48_p_reset = p_reset;
   assign  _add_map_x_48_m_clock = m_clock;
   assign  _add_map_x_47_moto_org_near = ((_net_4906)?data_in_org133:10'b0)|
    ((_net_914)?data_in_org134:10'b0);
   assign  _add_map_x_47_moto_org_near1 = ((_net_4905)?data_in_org135:10'b0)|
    ((_net_913)?data_in_org132:10'b0);
   assign  _add_map_x_47_moto_org_near2 = ((_net_4904)?data_in_org102:10'b0)|
    ((_net_912)?data_in_org101:10'b0);
   assign  _add_map_x_47_moto_org_near3 = ((_net_4903)?data_in_org166:10'b0)|
    ((_net_911)?data_in_org165:10'b0);
   assign  _add_map_x_47_moto_org = ((_net_4902)?data_in_org134:10'b0)|
    ((_net_910)?data_in_org133:10'b0);
   assign  _add_map_x_47_sg_up = ((_net_4901)?sg_in133:2'b0)|
    ((_net_909)?sg_in134:2'b0);
   assign  _add_map_x_47_sg_down = ((_net_4900)?sg_in135:2'b0)|
    ((_net_908)?sg_in132:2'b0);
   assign  _add_map_x_47_sg_left = ((_net_4898)?sg_in166:2'b0)|
    ((_net_906)?sg_in165:2'b0);
   assign  _add_map_x_47_sg_right = ((_net_4899)?sg_in102:2'b0)|
    ((_net_907)?sg_in101:2'b0);
   assign  _add_map_x_47_wall_t_in = dig_w;
   assign  _add_map_x_47_moto = ((_net_4896)?data_in134:10'b0)|
    ((_net_904)?data_in133:10'b0);
   assign  _add_map_x_47_up = ((_net_4895)?data_in133:10'b0)|
    ((_net_903)?data_in134:10'b0);
   assign  _add_map_x_47_right = ((_net_4894)?data_in135:10'b0)|
    ((_net_902)?data_in132:10'b0);
   assign  _add_map_x_47_down = ((_net_4893)?data_in102:10'b0)|
    ((_net_901)?data_in101:10'b0);
   assign  _add_map_x_47_left = ((_net_4892)?data_in166:10'b0)|
    ((_net_900)?data_in165:10'b0);
   assign  _add_map_x_47_start = start;
   assign  _add_map_x_47_goal = goal;
   assign  _add_map_x_47_now = ((_net_4889)?10'b0010000110:10'b0)|
    ((_net_897)?10'b0010000101:10'b0);
   assign  _add_map_x_47_add_exe = (_net_4888|_net_896);
   assign  _add_map_x_47_p_reset = p_reset;
   assign  _add_map_x_47_m_clock = m_clock;
   assign  _add_map_x_46_moto_org_near = ((_net_4887)?data_in_org131:10'b0)|
    ((_net_895)?data_in_org132:10'b0);
   assign  _add_map_x_46_moto_org_near1 = ((_net_4886)?data_in_org133:10'b0)|
    ((_net_894)?data_in_org130:10'b0);
   assign  _add_map_x_46_moto_org_near2 = ((_net_4885)?data_in_org100:10'b0)|
    ((_net_893)?data_in_org99:10'b0);
   assign  _add_map_x_46_moto_org_near3 = ((_net_4884)?data_in_org164:10'b0)|
    ((_net_892)?data_in_org163:10'b0);
   assign  _add_map_x_46_moto_org = ((_net_4883)?data_in_org132:10'b0)|
    ((_net_891)?data_in_org131:10'b0);
   assign  _add_map_x_46_sg_up = ((_net_4882)?sg_in131:2'b0)|
    ((_net_890)?sg_in132:2'b0);
   assign  _add_map_x_46_sg_down = ((_net_4881)?sg_in133:2'b0)|
    ((_net_889)?sg_in130:2'b0);
   assign  _add_map_x_46_sg_left = ((_net_4879)?sg_in164:2'b0)|
    ((_net_887)?sg_in163:2'b0);
   assign  _add_map_x_46_sg_right = ((_net_4880)?sg_in100:2'b0)|
    ((_net_888)?sg_in99:2'b0);
   assign  _add_map_x_46_wall_t_in = dig_w;
   assign  _add_map_x_46_moto = ((_net_4877)?data_in132:10'b0)|
    ((_net_885)?data_in131:10'b0);
   assign  _add_map_x_46_up = ((_net_4876)?data_in131:10'b0)|
    ((_net_884)?data_in132:10'b0);
   assign  _add_map_x_46_right = ((_net_4875)?data_in133:10'b0)|
    ((_net_883)?data_in130:10'b0);
   assign  _add_map_x_46_down = ((_net_4874)?data_in100:10'b0)|
    ((_net_882)?data_in99:10'b0);
   assign  _add_map_x_46_left = ((_net_4873)?data_in164:10'b0)|
    ((_net_881)?data_in163:10'b0);
   assign  _add_map_x_46_start = start;
   assign  _add_map_x_46_goal = goal;
   assign  _add_map_x_46_now = ((_net_4870)?10'b0010000100:10'b0)|
    ((_net_878)?10'b0010000011:10'b0);
   assign  _add_map_x_46_add_exe = (_net_4869|_net_877);
   assign  _add_map_x_46_p_reset = p_reset;
   assign  _add_map_x_46_m_clock = m_clock;
   assign  _add_map_x_45_moto_org_near = ((_net_4868)?data_in_org129:10'b0)|
    ((_net_876)?data_in_org130:10'b0);
   assign  _add_map_x_45_moto_org_near1 = ((_net_4867)?data_in_org131:10'b0)|
    ((_net_875)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_45_moto_org_near2 = ((_net_4866)?data_in_org98:10'b0)|
    ((_net_874)?data_in_org97:10'b0);
   assign  _add_map_x_45_moto_org_near3 = ((_net_4865)?data_in_org162:10'b0)|
    ((_net_873)?data_in_org161:10'b0);
   assign  _add_map_x_45_moto_org = ((_net_4864)?data_in_org130:10'b0)|
    ((_net_872)?data_in_org129:10'b0);
   assign  _add_map_x_45_sg_up = ((_net_4863)?sg_in129:2'b0)|
    ((_net_871)?sg_in130:2'b0);
   assign  _add_map_x_45_sg_down = ((_net_4862)?sg_in131:2'b0)|
    ((_net_870)?3'b000:2'b0);
   assign  _add_map_x_45_sg_left = ((_net_4860)?sg_in162:2'b0)|
    ((_net_868)?sg_in161:2'b0);
   assign  _add_map_x_45_sg_right = ((_net_4861)?sg_in98:2'b0)|
    ((_net_869)?sg_in97:2'b0);
   assign  _add_map_x_45_wall_t_in = dig_w;
   assign  _add_map_x_45_moto = ((_net_4858)?data_in130:10'b0)|
    ((_net_866)?data_in129:10'b0);
   assign  _add_map_x_45_up = ((_net_4857)?data_in129:10'b0)|
    ((_net_865)?data_in130:10'b0);
   assign  _add_map_x_45_right = ((_net_4856)?data_in131:10'b0)|
    ((_net_864)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_45_down = ((_net_4855)?data_in98:10'b0)|
    ((_net_863)?data_in97:10'b0);
   assign  _add_map_x_45_left = ((_net_4854)?data_in162:10'b0)|
    ((_net_862)?data_in161:10'b0);
   assign  _add_map_x_45_start = start;
   assign  _add_map_x_45_goal = goal;
   assign  _add_map_x_45_now = ((_net_4851)?10'b0010000010:10'b0)|
    ((_net_859)?10'b0010000001:10'b0);
   assign  _add_map_x_45_add_exe = (_net_4850|_net_858);
   assign  _add_map_x_45_p_reset = p_reset;
   assign  _add_map_x_45_m_clock = m_clock;
   assign  _add_map_x_44_moto_org_near = ((_net_4849)?data_in_org126:10'b0)|
    ((_net_857)?data_in_org125:10'b0);
   assign  _add_map_x_44_moto_org_near1 = ((_net_4848)?data_in_org124:10'b0)|
    ((_net_856)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_44_moto_org_near2 = ((_net_4847)?data_in_org93:10'b0)|
    ((_net_855)?data_in_org94:10'b0);
   assign  _add_map_x_44_moto_org_near3 = ((_net_4846)?data_in_org157:10'b0)|
    ((_net_854)?data_in_org158:10'b0);
   assign  _add_map_x_44_moto_org = ((_net_4845)?data_in_org125:10'b0)|
    ((_net_853)?data_in_org126:10'b0);
   assign  _add_map_x_44_sg_up = ((_net_4844)?sg_in126:2'b0)|
    ((_net_852)?sg_in125:2'b0);
   assign  _add_map_x_44_sg_down = ((_net_4843)?sg_in93:2'b0)|
    ((_net_851)?3'b000:2'b0);
   assign  _add_map_x_44_sg_left = ((_net_4841)?sg_in157:2'b0)|
    ((_net_849)?sg_in158:2'b0);
   assign  _add_map_x_44_sg_right = ((_net_4842)?sg_in124:2'b0)|
    ((_net_850)?sg_in94:2'b0);
   assign  _add_map_x_44_wall_t_in = dig_w;
   assign  _add_map_x_44_moto = ((_net_4839)?data_in125:10'b0)|
    ((_net_847)?data_in126:10'b0);
   assign  _add_map_x_44_up = ((_net_4838)?data_in126:10'b0)|
    ((_net_846)?data_in125:10'b0);
   assign  _add_map_x_44_right = ((_net_4837)?data_in124:10'b0)|
    ((_net_845)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_44_down = ((_net_4836)?data_in93:10'b0)|
    ((_net_844)?data_in94:10'b0);
   assign  _add_map_x_44_left = ((_net_4835)?data_in157:10'b0)|
    ((_net_843)?data_in158:10'b0);
   assign  _add_map_x_44_start = start;
   assign  _add_map_x_44_goal = goal;
   assign  _add_map_x_44_now = ((_net_4832)?10'b0001111101:10'b0)|
    ((_net_840)?10'b0001111110:10'b0);
   assign  _add_map_x_44_add_exe = (_net_4831|_net_839);
   assign  _add_map_x_44_p_reset = p_reset;
   assign  _add_map_x_44_m_clock = m_clock;
   assign  _add_map_x_43_moto_org_near = ((_net_4830)?data_in_org124:10'b0)|
    ((_net_838)?data_in_org123:10'b0);
   assign  _add_map_x_43_moto_org_near1 = ((_net_4829)?data_in_org122:10'b0)|
    ((_net_837)?data_in_org125:10'b0);
   assign  _add_map_x_43_moto_org_near2 = ((_net_4828)?data_in_org91:10'b0)|
    ((_net_836)?data_in_org92:10'b0);
   assign  _add_map_x_43_moto_org_near3 = ((_net_4827)?data_in_org155:10'b0)|
    ((_net_835)?data_in_org156:10'b0);
   assign  _add_map_x_43_moto_org = ((_net_4826)?data_in_org123:10'b0)|
    ((_net_834)?data_in_org124:10'b0);
   assign  _add_map_x_43_sg_up = ((_net_4825)?sg_in124:2'b0)|
    ((_net_833)?sg_in123:2'b0);
   assign  _add_map_x_43_sg_down = ((_net_4824)?sg_in91:2'b0)|
    ((_net_832)?sg_in125:2'b0);
   assign  _add_map_x_43_sg_left = ((_net_4822)?sg_in155:2'b0)|
    ((_net_830)?sg_in156:2'b0);
   assign  _add_map_x_43_sg_right = ((_net_4823)?sg_in122:2'b0)|
    ((_net_831)?sg_in92:2'b0);
   assign  _add_map_x_43_wall_t_in = dig_w;
   assign  _add_map_x_43_moto = ((_net_4820)?data_in123:10'b0)|
    ((_net_828)?data_in124:10'b0);
   assign  _add_map_x_43_up = ((_net_4819)?data_in124:10'b0)|
    ((_net_827)?data_in123:10'b0);
   assign  _add_map_x_43_right = ((_net_4818)?data_in122:10'b0)|
    ((_net_826)?data_in125:10'b0);
   assign  _add_map_x_43_down = ((_net_4817)?data_in91:10'b0)|
    ((_net_825)?data_in92:10'b0);
   assign  _add_map_x_43_left = ((_net_4816)?data_in155:10'b0)|
    ((_net_824)?data_in156:10'b0);
   assign  _add_map_x_43_start = start;
   assign  _add_map_x_43_goal = goal;
   assign  _add_map_x_43_now = ((_net_4813)?10'b0001111011:10'b0)|
    ((_net_821)?10'b0001111100:10'b0);
   assign  _add_map_x_43_add_exe = (_net_4812|_net_820);
   assign  _add_map_x_43_p_reset = p_reset;
   assign  _add_map_x_43_m_clock = m_clock;
   assign  _add_map_x_42_moto_org_near = ((_net_4811)?data_in_org122:10'b0)|
    ((_net_819)?data_in_org121:10'b0);
   assign  _add_map_x_42_moto_org_near1 = ((_net_4810)?data_in_org120:10'b0)|
    ((_net_818)?data_in_org123:10'b0);
   assign  _add_map_x_42_moto_org_near2 = ((_net_4809)?data_in_org89:10'b0)|
    ((_net_817)?data_in_org90:10'b0);
   assign  _add_map_x_42_moto_org_near3 = ((_net_4808)?data_in_org153:10'b0)|
    ((_net_816)?data_in_org154:10'b0);
   assign  _add_map_x_42_moto_org = ((_net_4807)?data_in_org121:10'b0)|
    ((_net_815)?data_in_org122:10'b0);
   assign  _add_map_x_42_sg_up = ((_net_4806)?sg_in122:2'b0)|
    ((_net_814)?sg_in121:2'b0);
   assign  _add_map_x_42_sg_down = ((_net_4805)?sg_in89:2'b0)|
    ((_net_813)?sg_in123:2'b0);
   assign  _add_map_x_42_sg_left = ((_net_4803)?sg_in153:2'b0)|
    ((_net_811)?sg_in154:2'b0);
   assign  _add_map_x_42_sg_right = ((_net_4804)?sg_in120:2'b0)|
    ((_net_812)?sg_in90:2'b0);
   assign  _add_map_x_42_wall_t_in = dig_w;
   assign  _add_map_x_42_moto = ((_net_4801)?data_in121:10'b0)|
    ((_net_809)?data_in122:10'b0);
   assign  _add_map_x_42_up = ((_net_4800)?data_in122:10'b0)|
    ((_net_808)?data_in121:10'b0);
   assign  _add_map_x_42_right = ((_net_4799)?data_in120:10'b0)|
    ((_net_807)?data_in123:10'b0);
   assign  _add_map_x_42_down = ((_net_4798)?data_in89:10'b0)|
    ((_net_806)?data_in90:10'b0);
   assign  _add_map_x_42_left = ((_net_4797)?data_in153:10'b0)|
    ((_net_805)?data_in154:10'b0);
   assign  _add_map_x_42_start = start;
   assign  _add_map_x_42_goal = goal;
   assign  _add_map_x_42_now = ((_net_4794)?10'b0001111001:10'b0)|
    ((_net_802)?10'b0001111010:10'b0);
   assign  _add_map_x_42_add_exe = (_net_4793|_net_801);
   assign  _add_map_x_42_p_reset = p_reset;
   assign  _add_map_x_42_m_clock = m_clock;
   assign  _add_map_x_41_moto_org_near = ((_net_4792)?data_in_org120:10'b0)|
    ((_net_800)?data_in_org119:10'b0);
   assign  _add_map_x_41_moto_org_near1 = ((_net_4791)?data_in_org118:10'b0)|
    ((_net_799)?data_in_org121:10'b0);
   assign  _add_map_x_41_moto_org_near2 = ((_net_4790)?data_in_org87:10'b0)|
    ((_net_798)?data_in_org88:10'b0);
   assign  _add_map_x_41_moto_org_near3 = ((_net_4789)?data_in_org151:10'b0)|
    ((_net_797)?data_in_org152:10'b0);
   assign  _add_map_x_41_moto_org = ((_net_4788)?data_in_org119:10'b0)|
    ((_net_796)?data_in_org120:10'b0);
   assign  _add_map_x_41_sg_up = ((_net_4787)?sg_in120:2'b0)|
    ((_net_795)?sg_in119:2'b0);
   assign  _add_map_x_41_sg_down = ((_net_4786)?sg_in87:2'b0)|
    ((_net_794)?sg_in121:2'b0);
   assign  _add_map_x_41_sg_left = ((_net_4784)?sg_in151:2'b0)|
    ((_net_792)?sg_in152:2'b0);
   assign  _add_map_x_41_sg_right = ((_net_4785)?sg_in118:2'b0)|
    ((_net_793)?sg_in88:2'b0);
   assign  _add_map_x_41_wall_t_in = dig_w;
   assign  _add_map_x_41_moto = ((_net_4782)?data_in119:10'b0)|
    ((_net_790)?data_in120:10'b0);
   assign  _add_map_x_41_up = ((_net_4781)?data_in120:10'b0)|
    ((_net_789)?data_in119:10'b0);
   assign  _add_map_x_41_right = ((_net_4780)?data_in118:10'b0)|
    ((_net_788)?data_in121:10'b0);
   assign  _add_map_x_41_down = ((_net_4779)?data_in87:10'b0)|
    ((_net_787)?data_in88:10'b0);
   assign  _add_map_x_41_left = ((_net_4778)?data_in151:10'b0)|
    ((_net_786)?data_in152:10'b0);
   assign  _add_map_x_41_start = start;
   assign  _add_map_x_41_goal = goal;
   assign  _add_map_x_41_now = ((_net_4775)?10'b0001110111:10'b0)|
    ((_net_783)?10'b0001111000:10'b0);
   assign  _add_map_x_41_add_exe = (_net_4774|_net_782);
   assign  _add_map_x_41_p_reset = p_reset;
   assign  _add_map_x_41_m_clock = m_clock;
   assign  _add_map_x_40_moto_org_near = ((_net_4773)?data_in_org118:10'b0)|
    ((_net_781)?data_in_org117:10'b0);
   assign  _add_map_x_40_moto_org_near1 = ((_net_4772)?data_in_org116:10'b0)|
    ((_net_780)?data_in_org119:10'b0);
   assign  _add_map_x_40_moto_org_near2 = ((_net_4771)?data_in_org85:10'b0)|
    ((_net_779)?data_in_org86:10'b0);
   assign  _add_map_x_40_moto_org_near3 = ((_net_4770)?data_in_org149:10'b0)|
    ((_net_778)?data_in_org150:10'b0);
   assign  _add_map_x_40_moto_org = ((_net_4769)?data_in_org117:10'b0)|
    ((_net_777)?data_in_org118:10'b0);
   assign  _add_map_x_40_sg_up = ((_net_4768)?sg_in118:2'b0)|
    ((_net_776)?sg_in117:2'b0);
   assign  _add_map_x_40_sg_down = ((_net_4767)?sg_in85:2'b0)|
    ((_net_775)?sg_in119:2'b0);
   assign  _add_map_x_40_sg_left = ((_net_4765)?sg_in149:2'b0)|
    ((_net_773)?sg_in150:2'b0);
   assign  _add_map_x_40_sg_right = ((_net_4766)?sg_in116:2'b0)|
    ((_net_774)?sg_in86:2'b0);
   assign  _add_map_x_40_wall_t_in = dig_w;
   assign  _add_map_x_40_moto = ((_net_4763)?data_in117:10'b0)|
    ((_net_771)?data_in118:10'b0);
   assign  _add_map_x_40_up = ((_net_4762)?data_in118:10'b0)|
    ((_net_770)?data_in117:10'b0);
   assign  _add_map_x_40_right = ((_net_4761)?data_in116:10'b0)|
    ((_net_769)?data_in119:10'b0);
   assign  _add_map_x_40_down = ((_net_4760)?data_in85:10'b0)|
    ((_net_768)?data_in86:10'b0);
   assign  _add_map_x_40_left = ((_net_4759)?data_in149:10'b0)|
    ((_net_767)?data_in150:10'b0);
   assign  _add_map_x_40_start = start;
   assign  _add_map_x_40_goal = goal;
   assign  _add_map_x_40_now = ((_net_4756)?10'b0001110101:10'b0)|
    ((_net_764)?10'b0001110110:10'b0);
   assign  _add_map_x_40_add_exe = (_net_4755|_net_763);
   assign  _add_map_x_40_p_reset = p_reset;
   assign  _add_map_x_40_m_clock = m_clock;
   assign  _add_map_x_39_moto_org_near = ((_net_4754)?data_in_org116:10'b0)|
    ((_net_762)?data_in_org115:10'b0);
   assign  _add_map_x_39_moto_org_near1 = ((_net_4753)?data_in_org114:10'b0)|
    ((_net_761)?data_in_org117:10'b0);
   assign  _add_map_x_39_moto_org_near2 = ((_net_4752)?data_in_org83:10'b0)|
    ((_net_760)?data_in_org84:10'b0);
   assign  _add_map_x_39_moto_org_near3 = ((_net_4751)?data_in_org147:10'b0)|
    ((_net_759)?data_in_org148:10'b0);
   assign  _add_map_x_39_moto_org = ((_net_4750)?data_in_org115:10'b0)|
    ((_net_758)?data_in_org116:10'b0);
   assign  _add_map_x_39_sg_up = ((_net_4749)?sg_in116:2'b0)|
    ((_net_757)?sg_in115:2'b0);
   assign  _add_map_x_39_sg_down = ((_net_4748)?sg_in83:2'b0)|
    ((_net_756)?sg_in117:2'b0);
   assign  _add_map_x_39_sg_left = ((_net_4746)?sg_in147:2'b0)|
    ((_net_754)?sg_in148:2'b0);
   assign  _add_map_x_39_sg_right = ((_net_4747)?sg_in114:2'b0)|
    ((_net_755)?sg_in84:2'b0);
   assign  _add_map_x_39_wall_t_in = dig_w;
   assign  _add_map_x_39_moto = ((_net_4744)?data_in115:10'b0)|
    ((_net_752)?data_in116:10'b0);
   assign  _add_map_x_39_up = ((_net_4743)?data_in116:10'b0)|
    ((_net_751)?data_in115:10'b0);
   assign  _add_map_x_39_right = ((_net_4742)?data_in114:10'b0)|
    ((_net_750)?data_in117:10'b0);
   assign  _add_map_x_39_down = ((_net_4741)?data_in83:10'b0)|
    ((_net_749)?data_in84:10'b0);
   assign  _add_map_x_39_left = ((_net_4740)?data_in147:10'b0)|
    ((_net_748)?data_in148:10'b0);
   assign  _add_map_x_39_start = start;
   assign  _add_map_x_39_goal = goal;
   assign  _add_map_x_39_now = ((_net_4737)?10'b0001110011:10'b0)|
    ((_net_745)?10'b0001110100:10'b0);
   assign  _add_map_x_39_add_exe = (_net_4736|_net_744);
   assign  _add_map_x_39_p_reset = p_reset;
   assign  _add_map_x_39_m_clock = m_clock;
   assign  _add_map_x_38_moto_org_near = ((_net_4735)?data_in_org114:10'b0)|
    ((_net_743)?data_in_org113:10'b0);
   assign  _add_map_x_38_moto_org_near1 = ((_net_4734)?data_in_org112:10'b0)|
    ((_net_742)?data_in_org115:10'b0);
   assign  _add_map_x_38_moto_org_near2 = ((_net_4733)?data_in_org81:10'b0)|
    ((_net_741)?data_in_org82:10'b0);
   assign  _add_map_x_38_moto_org_near3 = ((_net_4732)?data_in_org145:10'b0)|
    ((_net_740)?data_in_org146:10'b0);
   assign  _add_map_x_38_moto_org = ((_net_4731)?data_in_org113:10'b0)|
    ((_net_739)?data_in_org114:10'b0);
   assign  _add_map_x_38_sg_up = ((_net_4730)?sg_in114:2'b0)|
    ((_net_738)?sg_in113:2'b0);
   assign  _add_map_x_38_sg_down = ((_net_4729)?sg_in81:2'b0)|
    ((_net_737)?sg_in115:2'b0);
   assign  _add_map_x_38_sg_left = ((_net_4727)?sg_in145:2'b0)|
    ((_net_735)?sg_in146:2'b0);
   assign  _add_map_x_38_sg_right = ((_net_4728)?sg_in112:2'b0)|
    ((_net_736)?sg_in82:2'b0);
   assign  _add_map_x_38_wall_t_in = dig_w;
   assign  _add_map_x_38_moto = ((_net_4725)?data_in113:10'b0)|
    ((_net_733)?data_in114:10'b0);
   assign  _add_map_x_38_up = ((_net_4724)?data_in114:10'b0)|
    ((_net_732)?data_in113:10'b0);
   assign  _add_map_x_38_right = ((_net_4723)?data_in112:10'b0)|
    ((_net_731)?data_in115:10'b0);
   assign  _add_map_x_38_down = ((_net_4722)?data_in81:10'b0)|
    ((_net_730)?data_in82:10'b0);
   assign  _add_map_x_38_left = ((_net_4721)?data_in145:10'b0)|
    ((_net_729)?data_in146:10'b0);
   assign  _add_map_x_38_start = start;
   assign  _add_map_x_38_goal = goal;
   assign  _add_map_x_38_now = ((_net_4718)?10'b0001110001:10'b0)|
    ((_net_726)?10'b0001110010:10'b0);
   assign  _add_map_x_38_add_exe = (_net_4717|_net_725);
   assign  _add_map_x_38_p_reset = p_reset;
   assign  _add_map_x_38_m_clock = m_clock;
   assign  _add_map_x_37_moto_org_near = ((_net_4716)?data_in_org112:10'b0)|
    ((_net_724)?data_in_org111:10'b0);
   assign  _add_map_x_37_moto_org_near1 = ((_net_4715)?data_in_org110:10'b0)|
    ((_net_723)?data_in_org113:10'b0);
   assign  _add_map_x_37_moto_org_near2 = ((_net_4714)?data_in_org79:10'b0)|
    ((_net_722)?data_in_org80:10'b0);
   assign  _add_map_x_37_moto_org_near3 = ((_net_4713)?data_in_org143:10'b0)|
    ((_net_721)?data_in_org144:10'b0);
   assign  _add_map_x_37_moto_org = ((_net_4712)?data_in_org111:10'b0)|
    ((_net_720)?data_in_org112:10'b0);
   assign  _add_map_x_37_sg_up = ((_net_4711)?sg_in112:2'b0)|
    ((_net_719)?sg_in111:2'b0);
   assign  _add_map_x_37_sg_down = ((_net_4710)?sg_in79:2'b0)|
    ((_net_718)?sg_in113:2'b0);
   assign  _add_map_x_37_sg_left = ((_net_4708)?sg_in143:2'b0)|
    ((_net_716)?sg_in144:2'b0);
   assign  _add_map_x_37_sg_right = ((_net_4709)?sg_in110:2'b0)|
    ((_net_717)?sg_in80:2'b0);
   assign  _add_map_x_37_wall_t_in = dig_w;
   assign  _add_map_x_37_moto = ((_net_4706)?data_in111:10'b0)|
    ((_net_714)?data_in112:10'b0);
   assign  _add_map_x_37_up = ((_net_4705)?data_in112:10'b0)|
    ((_net_713)?data_in111:10'b0);
   assign  _add_map_x_37_right = ((_net_4704)?data_in110:10'b0)|
    ((_net_712)?data_in113:10'b0);
   assign  _add_map_x_37_down = ((_net_4703)?data_in79:10'b0)|
    ((_net_711)?data_in80:10'b0);
   assign  _add_map_x_37_left = ((_net_4702)?data_in143:10'b0)|
    ((_net_710)?data_in144:10'b0);
   assign  _add_map_x_37_start = start;
   assign  _add_map_x_37_goal = goal;
   assign  _add_map_x_37_now = ((_net_4699)?10'b0001101111:10'b0)|
    ((_net_707)?10'b0001110000:10'b0);
   assign  _add_map_x_37_add_exe = (_net_4698|_net_706);
   assign  _add_map_x_37_p_reset = p_reset;
   assign  _add_map_x_37_m_clock = m_clock;
   assign  _add_map_x_36_moto_org_near = ((_net_4697)?data_in_org110:10'b0)|
    ((_net_705)?data_in_org109:10'b0);
   assign  _add_map_x_36_moto_org_near1 = ((_net_4696)?data_in_org108:10'b0)|
    ((_net_704)?data_in_org111:10'b0);
   assign  _add_map_x_36_moto_org_near2 = ((_net_4695)?data_in_org77:10'b0)|
    ((_net_703)?data_in_org78:10'b0);
   assign  _add_map_x_36_moto_org_near3 = ((_net_4694)?data_in_org141:10'b0)|
    ((_net_702)?data_in_org142:10'b0);
   assign  _add_map_x_36_moto_org = ((_net_4693)?data_in_org109:10'b0)|
    ((_net_701)?data_in_org110:10'b0);
   assign  _add_map_x_36_sg_up = ((_net_4692)?sg_in110:2'b0)|
    ((_net_700)?sg_in109:2'b0);
   assign  _add_map_x_36_sg_down = ((_net_4691)?sg_in77:2'b0)|
    ((_net_699)?sg_in111:2'b0);
   assign  _add_map_x_36_sg_left = ((_net_4689)?sg_in141:2'b0)|
    ((_net_697)?sg_in142:2'b0);
   assign  _add_map_x_36_sg_right = ((_net_4690)?sg_in108:2'b0)|
    ((_net_698)?sg_in78:2'b0);
   assign  _add_map_x_36_wall_t_in = dig_w;
   assign  _add_map_x_36_moto = ((_net_4687)?data_in109:10'b0)|
    ((_net_695)?data_in110:10'b0);
   assign  _add_map_x_36_up = ((_net_4686)?data_in110:10'b0)|
    ((_net_694)?data_in109:10'b0);
   assign  _add_map_x_36_right = ((_net_4685)?data_in108:10'b0)|
    ((_net_693)?data_in111:10'b0);
   assign  _add_map_x_36_down = ((_net_4684)?data_in77:10'b0)|
    ((_net_692)?data_in78:10'b0);
   assign  _add_map_x_36_left = ((_net_4683)?data_in141:10'b0)|
    ((_net_691)?data_in142:10'b0);
   assign  _add_map_x_36_start = start;
   assign  _add_map_x_36_goal = goal;
   assign  _add_map_x_36_now = ((_net_4680)?10'b0001101101:10'b0)|
    ((_net_688)?10'b0001101110:10'b0);
   assign  _add_map_x_36_add_exe = (_net_4679|_net_687);
   assign  _add_map_x_36_p_reset = p_reset;
   assign  _add_map_x_36_m_clock = m_clock;
   assign  _add_map_x_35_moto_org_near = ((_net_4678)?data_in_org108:10'b0)|
    ((_net_686)?data_in_org107:10'b0);
   assign  _add_map_x_35_moto_org_near1 = ((_net_4677)?data_in_org106:10'b0)|
    ((_net_685)?data_in_org109:10'b0);
   assign  _add_map_x_35_moto_org_near2 = ((_net_4676)?data_in_org75:10'b0)|
    ((_net_684)?data_in_org76:10'b0);
   assign  _add_map_x_35_moto_org_near3 = ((_net_4675)?data_in_org139:10'b0)|
    ((_net_683)?data_in_org140:10'b0);
   assign  _add_map_x_35_moto_org = ((_net_4674)?data_in_org107:10'b0)|
    ((_net_682)?data_in_org108:10'b0);
   assign  _add_map_x_35_sg_up = ((_net_4673)?sg_in108:2'b0)|
    ((_net_681)?sg_in107:2'b0);
   assign  _add_map_x_35_sg_down = ((_net_4672)?sg_in75:2'b0)|
    ((_net_680)?sg_in109:2'b0);
   assign  _add_map_x_35_sg_left = ((_net_4670)?sg_in139:2'b0)|
    ((_net_678)?sg_in140:2'b0);
   assign  _add_map_x_35_sg_right = ((_net_4671)?sg_in106:2'b0)|
    ((_net_679)?sg_in76:2'b0);
   assign  _add_map_x_35_wall_t_in = dig_w;
   assign  _add_map_x_35_moto = ((_net_4668)?data_in107:10'b0)|
    ((_net_676)?data_in108:10'b0);
   assign  _add_map_x_35_up = ((_net_4667)?data_in108:10'b0)|
    ((_net_675)?data_in107:10'b0);
   assign  _add_map_x_35_right = ((_net_4666)?data_in106:10'b0)|
    ((_net_674)?data_in109:10'b0);
   assign  _add_map_x_35_down = ((_net_4665)?data_in75:10'b0)|
    ((_net_673)?data_in76:10'b0);
   assign  _add_map_x_35_left = ((_net_4664)?data_in139:10'b0)|
    ((_net_672)?data_in140:10'b0);
   assign  _add_map_x_35_start = start;
   assign  _add_map_x_35_goal = goal;
   assign  _add_map_x_35_now = ((_net_4661)?10'b0001101011:10'b0)|
    ((_net_669)?10'b0001101100:10'b0);
   assign  _add_map_x_35_add_exe = (_net_4660|_net_668);
   assign  _add_map_x_35_p_reset = p_reset;
   assign  _add_map_x_35_m_clock = m_clock;
   assign  _add_map_x_34_moto_org_near = ((_net_4659)?data_in_org106:10'b0)|
    ((_net_667)?data_in_org105:10'b0);
   assign  _add_map_x_34_moto_org_near1 = ((_net_4658)?data_in_org104:10'b0)|
    ((_net_666)?data_in_org107:10'b0);
   assign  _add_map_x_34_moto_org_near2 = ((_net_4657)?data_in_org73:10'b0)|
    ((_net_665)?data_in_org74:10'b0);
   assign  _add_map_x_34_moto_org_near3 = ((_net_4656)?data_in_org137:10'b0)|
    ((_net_664)?data_in_org138:10'b0);
   assign  _add_map_x_34_moto_org = ((_net_4655)?data_in_org105:10'b0)|
    ((_net_663)?data_in_org106:10'b0);
   assign  _add_map_x_34_sg_up = ((_net_4654)?sg_in106:2'b0)|
    ((_net_662)?sg_in105:2'b0);
   assign  _add_map_x_34_sg_down = ((_net_4653)?sg_in73:2'b0)|
    ((_net_661)?sg_in107:2'b0);
   assign  _add_map_x_34_sg_left = ((_net_4651)?sg_in137:2'b0)|
    ((_net_659)?sg_in138:2'b0);
   assign  _add_map_x_34_sg_right = ((_net_4652)?sg_in104:2'b0)|
    ((_net_660)?sg_in74:2'b0);
   assign  _add_map_x_34_wall_t_in = dig_w;
   assign  _add_map_x_34_moto = ((_net_4649)?data_in105:10'b0)|
    ((_net_657)?data_in106:10'b0);
   assign  _add_map_x_34_up = ((_net_4648)?data_in106:10'b0)|
    ((_net_656)?data_in105:10'b0);
   assign  _add_map_x_34_right = ((_net_4647)?data_in104:10'b0)|
    ((_net_655)?data_in107:10'b0);
   assign  _add_map_x_34_down = ((_net_4646)?data_in73:10'b0)|
    ((_net_654)?data_in74:10'b0);
   assign  _add_map_x_34_left = ((_net_4645)?data_in137:10'b0)|
    ((_net_653)?data_in138:10'b0);
   assign  _add_map_x_34_start = start;
   assign  _add_map_x_34_goal = goal;
   assign  _add_map_x_34_now = ((_net_4642)?10'b0001101001:10'b0)|
    ((_net_650)?10'b0001101010:10'b0);
   assign  _add_map_x_34_add_exe = (_net_4641|_net_649);
   assign  _add_map_x_34_p_reset = p_reset;
   assign  _add_map_x_34_m_clock = m_clock;
   assign  _add_map_x_33_moto_org_near = ((_net_4640)?data_in_org104:10'b0)|
    ((_net_648)?data_in_org103:10'b0);
   assign  _add_map_x_33_moto_org_near1 = ((_net_4639)?data_in_org102:10'b0)|
    ((_net_647)?data_in_org105:10'b0);
   assign  _add_map_x_33_moto_org_near2 = ((_net_4638)?data_in_org71:10'b0)|
    ((_net_646)?data_in_org72:10'b0);
   assign  _add_map_x_33_moto_org_near3 = ((_net_4637)?data_in_org135:10'b0)|
    ((_net_645)?data_in_org136:10'b0);
   assign  _add_map_x_33_moto_org = ((_net_4636)?data_in_org103:10'b0)|
    ((_net_644)?data_in_org104:10'b0);
   assign  _add_map_x_33_sg_up = ((_net_4635)?sg_in104:2'b0)|
    ((_net_643)?sg_in103:2'b0);
   assign  _add_map_x_33_sg_down = ((_net_4634)?sg_in71:2'b0)|
    ((_net_642)?sg_in105:2'b0);
   assign  _add_map_x_33_sg_left = ((_net_4632)?sg_in135:2'b0)|
    ((_net_640)?sg_in136:2'b0);
   assign  _add_map_x_33_sg_right = ((_net_4633)?sg_in102:2'b0)|
    ((_net_641)?sg_in72:2'b0);
   assign  _add_map_x_33_wall_t_in = dig_w;
   assign  _add_map_x_33_moto = ((_net_4630)?data_in103:10'b0)|
    ((_net_638)?data_in104:10'b0);
   assign  _add_map_x_33_up = ((_net_4629)?data_in104:10'b0)|
    ((_net_637)?data_in103:10'b0);
   assign  _add_map_x_33_right = ((_net_4628)?data_in102:10'b0)|
    ((_net_636)?data_in105:10'b0);
   assign  _add_map_x_33_down = ((_net_4627)?data_in71:10'b0)|
    ((_net_635)?data_in72:10'b0);
   assign  _add_map_x_33_left = ((_net_4626)?data_in135:10'b0)|
    ((_net_634)?data_in136:10'b0);
   assign  _add_map_x_33_start = start;
   assign  _add_map_x_33_goal = goal;
   assign  _add_map_x_33_now = ((_net_4623)?10'b0001100111:10'b0)|
    ((_net_631)?10'b0001101000:10'b0);
   assign  _add_map_x_33_add_exe = (_net_4622|_net_630);
   assign  _add_map_x_33_p_reset = p_reset;
   assign  _add_map_x_33_m_clock = m_clock;
   assign  _add_map_x_32_moto_org_near = ((_net_4621)?data_in_org102:10'b0)|
    ((_net_629)?data_in_org101:10'b0);
   assign  _add_map_x_32_moto_org_near1 = ((_net_4620)?data_in_org100:10'b0)|
    ((_net_628)?data_in_org103:10'b0);
   assign  _add_map_x_32_moto_org_near2 = ((_net_4619)?data_in_org69:10'b0)|
    ((_net_627)?data_in_org70:10'b0);
   assign  _add_map_x_32_moto_org_near3 = ((_net_4618)?data_in_org133:10'b0)|
    ((_net_626)?data_in_org134:10'b0);
   assign  _add_map_x_32_moto_org = ((_net_4617)?data_in_org101:10'b0)|
    ((_net_625)?data_in_org102:10'b0);
   assign  _add_map_x_32_sg_up = ((_net_4616)?sg_in102:2'b0)|
    ((_net_624)?sg_in101:2'b0);
   assign  _add_map_x_32_sg_down = ((_net_4615)?sg_in69:2'b0)|
    ((_net_623)?sg_in103:2'b0);
   assign  _add_map_x_32_sg_left = ((_net_4613)?sg_in133:2'b0)|
    ((_net_621)?sg_in134:2'b0);
   assign  _add_map_x_32_sg_right = ((_net_4614)?sg_in100:2'b0)|
    ((_net_622)?sg_in70:2'b0);
   assign  _add_map_x_32_wall_t_in = dig_w;
   assign  _add_map_x_32_moto = ((_net_4611)?data_in101:10'b0)|
    ((_net_619)?data_in102:10'b0);
   assign  _add_map_x_32_up = ((_net_4610)?data_in102:10'b0)|
    ((_net_618)?data_in101:10'b0);
   assign  _add_map_x_32_right = ((_net_4609)?data_in100:10'b0)|
    ((_net_617)?data_in103:10'b0);
   assign  _add_map_x_32_down = ((_net_4608)?data_in69:10'b0)|
    ((_net_616)?data_in70:10'b0);
   assign  _add_map_x_32_left = ((_net_4607)?data_in133:10'b0)|
    ((_net_615)?data_in134:10'b0);
   assign  _add_map_x_32_start = start;
   assign  _add_map_x_32_goal = goal;
   assign  _add_map_x_32_now = ((_net_4604)?10'b0001100101:10'b0)|
    ((_net_612)?10'b0001100110:10'b0);
   assign  _add_map_x_32_add_exe = (_net_4603|_net_611);
   assign  _add_map_x_32_p_reset = p_reset;
   assign  _add_map_x_32_m_clock = m_clock;
   assign  _add_map_x_31_moto_org_near = ((_net_4602)?data_in_org100:10'b0)|
    ((_net_610)?data_in_org99:10'b0);
   assign  _add_map_x_31_moto_org_near1 = ((_net_4601)?data_in_org98:10'b0)|
    ((_net_609)?data_in_org101:10'b0);
   assign  _add_map_x_31_moto_org_near2 = ((_net_4600)?data_in_org67:10'b0)|
    ((_net_608)?data_in_org68:10'b0);
   assign  _add_map_x_31_moto_org_near3 = ((_net_4599)?data_in_org131:10'b0)|
    ((_net_607)?data_in_org132:10'b0);
   assign  _add_map_x_31_moto_org = ((_net_4598)?data_in_org99:10'b0)|
    ((_net_606)?data_in_org100:10'b0);
   assign  _add_map_x_31_sg_up = ((_net_4597)?sg_in100:2'b0)|
    ((_net_605)?sg_in99:2'b0);
   assign  _add_map_x_31_sg_down = ((_net_4596)?sg_in67:2'b0)|
    ((_net_604)?sg_in101:2'b0);
   assign  _add_map_x_31_sg_left = ((_net_4594)?sg_in131:2'b0)|
    ((_net_602)?sg_in132:2'b0);
   assign  _add_map_x_31_sg_right = ((_net_4595)?sg_in98:2'b0)|
    ((_net_603)?sg_in68:2'b0);
   assign  _add_map_x_31_wall_t_in = dig_w;
   assign  _add_map_x_31_moto = ((_net_4592)?data_in99:10'b0)|
    ((_net_600)?data_in100:10'b0);
   assign  _add_map_x_31_up = ((_net_4591)?data_in100:10'b0)|
    ((_net_599)?data_in99:10'b0);
   assign  _add_map_x_31_right = ((_net_4590)?data_in98:10'b0)|
    ((_net_598)?data_in101:10'b0);
   assign  _add_map_x_31_down = ((_net_4589)?data_in67:10'b0)|
    ((_net_597)?data_in68:10'b0);
   assign  _add_map_x_31_left = ((_net_4588)?data_in131:10'b0)|
    ((_net_596)?data_in132:10'b0);
   assign  _add_map_x_31_start = start;
   assign  _add_map_x_31_goal = goal;
   assign  _add_map_x_31_now = ((_net_4585)?10'b0001100011:10'b0)|
    ((_net_593)?10'b0001100100:10'b0);
   assign  _add_map_x_31_add_exe = (_net_4584|_net_592);
   assign  _add_map_x_31_p_reset = p_reset;
   assign  _add_map_x_31_m_clock = m_clock;
   assign  _add_map_x_30_moto_org_near = ((_net_4583)?data_in_org98:10'b0)|
    ((_net_591)?data_in_org97:10'b0);
   assign  _add_map_x_30_moto_org_near1 = ((_net_4582)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_590)?data_in_org99:10'b0);
   assign  _add_map_x_30_moto_org_near2 = ((_net_4581)?data_in_org65:10'b0)|
    ((_net_589)?data_in_org66:10'b0);
   assign  _add_map_x_30_moto_org_near3 = ((_net_4580)?data_in_org129:10'b0)|
    ((_net_588)?data_in_org130:10'b0);
   assign  _add_map_x_30_moto_org = ((_net_4579)?data_in_org97:10'b0)|
    ((_net_587)?data_in_org98:10'b0);
   assign  _add_map_x_30_sg_up = ((_net_4578)?sg_in98:2'b0)|
    ((_net_586)?sg_in97:2'b0);
   assign  _add_map_x_30_sg_down = ((_net_4577)?sg_in65:2'b0)|
    ((_net_585)?sg_in99:2'b0);
   assign  _add_map_x_30_sg_left = ((_net_4575)?sg_in129:2'b0)|
    ((_net_583)?sg_in130:2'b0);
   assign  _add_map_x_30_sg_right = ((_net_4576)?3'b000:2'b0)|
    ((_net_584)?sg_in66:2'b0);
   assign  _add_map_x_30_wall_t_in = dig_w;
   assign  _add_map_x_30_moto = ((_net_4573)?data_in97:10'b0)|
    ((_net_581)?data_in98:10'b0);
   assign  _add_map_x_30_up = ((_net_4572)?data_in98:10'b0)|
    ((_net_580)?data_in97:10'b0);
   assign  _add_map_x_30_right = ((_net_4571)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_579)?data_in99:10'b0);
   assign  _add_map_x_30_down = ((_net_4570)?data_in65:10'b0)|
    ((_net_578)?data_in66:10'b0);
   assign  _add_map_x_30_left = ((_net_4569)?data_in129:10'b0)|
    ((_net_577)?data_in130:10'b0);
   assign  _add_map_x_30_start = start;
   assign  _add_map_x_30_goal = goal;
   assign  _add_map_x_30_now = ((_net_4566)?10'b0001100001:10'b0)|
    ((_net_574)?10'b0001100010:10'b0);
   assign  _add_map_x_30_add_exe = (_net_4565|_net_573);
   assign  _add_map_x_30_p_reset = p_reset;
   assign  _add_map_x_30_m_clock = m_clock;
   assign  _add_map_x_29_moto_org_near = ((_net_4564)?data_in_org93:10'b0)|
    ((_net_572)?data_in_org94:10'b0);
   assign  _add_map_x_29_moto_org_near1 = ((_net_4563)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_571)?data_in_org92:10'b0);
   assign  _add_map_x_29_moto_org_near2 = ((_net_4562)?data_in_org62:10'b0)|
    ((_net_570)?data_in_org61:10'b0);
   assign  _add_map_x_29_moto_org_near3 = ((_net_4561)?data_in_org126:10'b0)|
    ((_net_569)?data_in_org125:10'b0);
   assign  _add_map_x_29_moto_org = ((_net_4560)?data_in_org94:10'b0)|
    ((_net_568)?data_in_org93:10'b0);
   assign  _add_map_x_29_sg_up = ((_net_4559)?sg_in93:2'b0)|
    ((_net_567)?sg_in94:2'b0);
   assign  _add_map_x_29_sg_down = ((_net_4558)?3'b000:2'b0)|
    ((_net_566)?sg_in92:2'b0);
   assign  _add_map_x_29_sg_left = ((_net_4556)?sg_in126:2'b0)|
    ((_net_564)?sg_in125:2'b0);
   assign  _add_map_x_29_sg_right = ((_net_4557)?sg_in62:2'b0)|
    ((_net_565)?sg_in61:2'b0);
   assign  _add_map_x_29_wall_t_in = dig_w;
   assign  _add_map_x_29_moto = ((_net_4554)?data_in94:10'b0)|
    ((_net_562)?data_in93:10'b0);
   assign  _add_map_x_29_up = ((_net_4553)?data_in93:10'b0)|
    ((_net_561)?data_in94:10'b0);
   assign  _add_map_x_29_right = ((_net_4552)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0)|
    ((_net_560)?data_in92:10'b0);
   assign  _add_map_x_29_down = ((_net_4551)?data_in62:10'b0)|
    ((_net_559)?data_in61:10'b0);
   assign  _add_map_x_29_left = ((_net_4550)?data_in126:10'b0)|
    ((_net_558)?data_in125:10'b0);
   assign  _add_map_x_29_start = start;
   assign  _add_map_x_29_goal = goal;
   assign  _add_map_x_29_now = ((_net_4547)?10'b0001011110:10'b0)|
    ((_net_555)?10'b0001011101:10'b0);
   assign  _add_map_x_29_add_exe = (_net_4546|_net_554);
   assign  _add_map_x_29_p_reset = p_reset;
   assign  _add_map_x_29_m_clock = m_clock;
   assign  _add_map_x_28_moto_org_near = ((_net_4545)?data_in_org91:10'b0)|
    ((_net_553)?data_in_org92:10'b0);
   assign  _add_map_x_28_moto_org_near1 = ((_net_4544)?data_in_org93:10'b0)|
    ((_net_552)?data_in_org90:10'b0);
   assign  _add_map_x_28_moto_org_near2 = ((_net_4543)?data_in_org60:10'b0)|
    ((_net_551)?data_in_org59:10'b0);
   assign  _add_map_x_28_moto_org_near3 = ((_net_4542)?data_in_org124:10'b0)|
    ((_net_550)?data_in_org123:10'b0);
   assign  _add_map_x_28_moto_org = ((_net_4541)?data_in_org92:10'b0)|
    ((_net_549)?data_in_org91:10'b0);
   assign  _add_map_x_28_sg_up = ((_net_4540)?sg_in91:2'b0)|
    ((_net_548)?sg_in92:2'b0);
   assign  _add_map_x_28_sg_down = ((_net_4539)?sg_in93:2'b0)|
    ((_net_547)?sg_in90:2'b0);
   assign  _add_map_x_28_sg_left = ((_net_4537)?sg_in124:2'b0)|
    ((_net_545)?sg_in123:2'b0);
   assign  _add_map_x_28_sg_right = ((_net_4538)?sg_in60:2'b0)|
    ((_net_546)?sg_in59:2'b0);
   assign  _add_map_x_28_wall_t_in = dig_w;
   assign  _add_map_x_28_moto = ((_net_4535)?data_in92:10'b0)|
    ((_net_543)?data_in91:10'b0);
   assign  _add_map_x_28_up = ((_net_4534)?data_in91:10'b0)|
    ((_net_542)?data_in92:10'b0);
   assign  _add_map_x_28_right = ((_net_4533)?data_in93:10'b0)|
    ((_net_541)?data_in90:10'b0);
   assign  _add_map_x_28_down = ((_net_4532)?data_in60:10'b0)|
    ((_net_540)?data_in59:10'b0);
   assign  _add_map_x_28_left = ((_net_4531)?data_in124:10'b0)|
    ((_net_539)?data_in123:10'b0);
   assign  _add_map_x_28_start = start;
   assign  _add_map_x_28_goal = goal;
   assign  _add_map_x_28_now = ((_net_4528)?10'b0001011100:10'b0)|
    ((_net_536)?10'b0001011011:10'b0);
   assign  _add_map_x_28_add_exe = (_net_4527|_net_535);
   assign  _add_map_x_28_p_reset = p_reset;
   assign  _add_map_x_28_m_clock = m_clock;
   assign  _add_map_x_27_moto_org_near = ((_net_4526)?data_in_org89:10'b0)|
    ((_net_534)?data_in_org90:10'b0);
   assign  _add_map_x_27_moto_org_near1 = ((_net_4525)?data_in_org91:10'b0)|
    ((_net_533)?data_in_org88:10'b0);
   assign  _add_map_x_27_moto_org_near2 = ((_net_4524)?data_in_org58:10'b0)|
    ((_net_532)?data_in_org57:10'b0);
   assign  _add_map_x_27_moto_org_near3 = ((_net_4523)?data_in_org122:10'b0)|
    ((_net_531)?data_in_org121:10'b0);
   assign  _add_map_x_27_moto_org = ((_net_4522)?data_in_org90:10'b0)|
    ((_net_530)?data_in_org89:10'b0);
   assign  _add_map_x_27_sg_up = ((_net_4521)?sg_in89:2'b0)|
    ((_net_529)?sg_in90:2'b0);
   assign  _add_map_x_27_sg_down = ((_net_4520)?sg_in91:2'b0)|
    ((_net_528)?sg_in88:2'b0);
   assign  _add_map_x_27_sg_left = ((_net_4518)?sg_in122:2'b0)|
    ((_net_526)?sg_in121:2'b0);
   assign  _add_map_x_27_sg_right = ((_net_4519)?sg_in58:2'b0)|
    ((_net_527)?sg_in57:2'b0);
   assign  _add_map_x_27_wall_t_in = dig_w;
   assign  _add_map_x_27_moto = ((_net_4516)?data_in90:10'b0)|
    ((_net_524)?data_in89:10'b0);
   assign  _add_map_x_27_up = ((_net_4515)?data_in89:10'b0)|
    ((_net_523)?data_in90:10'b0);
   assign  _add_map_x_27_right = ((_net_4514)?data_in91:10'b0)|
    ((_net_522)?data_in88:10'b0);
   assign  _add_map_x_27_down = ((_net_4513)?data_in58:10'b0)|
    ((_net_521)?data_in57:10'b0);
   assign  _add_map_x_27_left = ((_net_4512)?data_in122:10'b0)|
    ((_net_520)?data_in121:10'b0);
   assign  _add_map_x_27_start = start;
   assign  _add_map_x_27_goal = goal;
   assign  _add_map_x_27_now = ((_net_4509)?10'b0001011010:10'b0)|
    ((_net_517)?10'b0001011001:10'b0);
   assign  _add_map_x_27_add_exe = (_net_4508|_net_516);
   assign  _add_map_x_27_p_reset = p_reset;
   assign  _add_map_x_27_m_clock = m_clock;
   assign  _add_map_x_26_moto_org_near = ((_net_4507)?data_in_org87:10'b0)|
    ((_net_515)?data_in_org88:10'b0);
   assign  _add_map_x_26_moto_org_near1 = ((_net_4506)?data_in_org89:10'b0)|
    ((_net_514)?data_in_org86:10'b0);
   assign  _add_map_x_26_moto_org_near2 = ((_net_4505)?data_in_org56:10'b0)|
    ((_net_513)?data_in_org55:10'b0);
   assign  _add_map_x_26_moto_org_near3 = ((_net_4504)?data_in_org120:10'b0)|
    ((_net_512)?data_in_org119:10'b0);
   assign  _add_map_x_26_moto_org = ((_net_4503)?data_in_org88:10'b0)|
    ((_net_511)?data_in_org87:10'b0);
   assign  _add_map_x_26_sg_up = ((_net_4502)?sg_in87:2'b0)|
    ((_net_510)?sg_in88:2'b0);
   assign  _add_map_x_26_sg_down = ((_net_4501)?sg_in89:2'b0)|
    ((_net_509)?sg_in86:2'b0);
   assign  _add_map_x_26_sg_left = ((_net_4499)?sg_in120:2'b0)|
    ((_net_507)?sg_in119:2'b0);
   assign  _add_map_x_26_sg_right = ((_net_4500)?sg_in56:2'b0)|
    ((_net_508)?sg_in55:2'b0);
   assign  _add_map_x_26_wall_t_in = dig_w;
   assign  _add_map_x_26_moto = ((_net_4497)?data_in88:10'b0)|
    ((_net_505)?data_in87:10'b0);
   assign  _add_map_x_26_up = ((_net_4496)?data_in87:10'b0)|
    ((_net_504)?data_in88:10'b0);
   assign  _add_map_x_26_right = ((_net_4495)?data_in89:10'b0)|
    ((_net_503)?data_in86:10'b0);
   assign  _add_map_x_26_down = ((_net_4494)?data_in56:10'b0)|
    ((_net_502)?data_in55:10'b0);
   assign  _add_map_x_26_left = ((_net_4493)?data_in120:10'b0)|
    ((_net_501)?data_in119:10'b0);
   assign  _add_map_x_26_start = start;
   assign  _add_map_x_26_goal = goal;
   assign  _add_map_x_26_now = ((_net_4490)?10'b0001011000:10'b0)|
    ((_net_498)?10'b0001010111:10'b0);
   assign  _add_map_x_26_add_exe = (_net_4489|_net_497);
   assign  _add_map_x_26_p_reset = p_reset;
   assign  _add_map_x_26_m_clock = m_clock;
   assign  _add_map_x_25_moto_org_near = ((_net_4488)?data_in_org85:10'b0)|
    ((_net_496)?data_in_org86:10'b0);
   assign  _add_map_x_25_moto_org_near1 = ((_net_4487)?data_in_org87:10'b0)|
    ((_net_495)?data_in_org84:10'b0);
   assign  _add_map_x_25_moto_org_near2 = ((_net_4486)?data_in_org54:10'b0)|
    ((_net_494)?data_in_org53:10'b0);
   assign  _add_map_x_25_moto_org_near3 = ((_net_4485)?data_in_org118:10'b0)|
    ((_net_493)?data_in_org117:10'b0);
   assign  _add_map_x_25_moto_org = ((_net_4484)?data_in_org86:10'b0)|
    ((_net_492)?data_in_org85:10'b0);
   assign  _add_map_x_25_sg_up = ((_net_4483)?sg_in85:2'b0)|
    ((_net_491)?sg_in86:2'b0);
   assign  _add_map_x_25_sg_down = ((_net_4482)?sg_in87:2'b0)|
    ((_net_490)?sg_in84:2'b0);
   assign  _add_map_x_25_sg_left = ((_net_4480)?sg_in118:2'b0)|
    ((_net_488)?sg_in117:2'b0);
   assign  _add_map_x_25_sg_right = ((_net_4481)?sg_in54:2'b0)|
    ((_net_489)?sg_in53:2'b0);
   assign  _add_map_x_25_wall_t_in = dig_w;
   assign  _add_map_x_25_moto = ((_net_4478)?data_in86:10'b0)|
    ((_net_486)?data_in85:10'b0);
   assign  _add_map_x_25_up = ((_net_4477)?data_in85:10'b0)|
    ((_net_485)?data_in86:10'b0);
   assign  _add_map_x_25_right = ((_net_4476)?data_in87:10'b0)|
    ((_net_484)?data_in84:10'b0);
   assign  _add_map_x_25_down = ((_net_4475)?data_in54:10'b0)|
    ((_net_483)?data_in53:10'b0);
   assign  _add_map_x_25_left = ((_net_4474)?data_in118:10'b0)|
    ((_net_482)?data_in117:10'b0);
   assign  _add_map_x_25_start = start;
   assign  _add_map_x_25_goal = goal;
   assign  _add_map_x_25_now = ((_net_4471)?10'b0001010110:10'b0)|
    ((_net_479)?10'b0001010101:10'b0);
   assign  _add_map_x_25_add_exe = (_net_4470|_net_478);
   assign  _add_map_x_25_p_reset = p_reset;
   assign  _add_map_x_25_m_clock = m_clock;
   assign  _add_map_x_24_moto_org_near = ((_net_4469)?data_in_org83:10'b0)|
    ((_net_477)?data_in_org84:10'b0);
   assign  _add_map_x_24_moto_org_near1 = ((_net_4468)?data_in_org85:10'b0)|
    ((_net_476)?data_in_org82:10'b0);
   assign  _add_map_x_24_moto_org_near2 = ((_net_4467)?data_in_org52:10'b0)|
    ((_net_475)?data_in_org51:10'b0);
   assign  _add_map_x_24_moto_org_near3 = ((_net_4466)?data_in_org116:10'b0)|
    ((_net_474)?data_in_org115:10'b0);
   assign  _add_map_x_24_moto_org = ((_net_4465)?data_in_org84:10'b0)|
    ((_net_473)?data_in_org83:10'b0);
   assign  _add_map_x_24_sg_up = ((_net_4464)?sg_in83:2'b0)|
    ((_net_472)?sg_in84:2'b0);
   assign  _add_map_x_24_sg_down = ((_net_4463)?sg_in85:2'b0)|
    ((_net_471)?sg_in82:2'b0);
   assign  _add_map_x_24_sg_left = ((_net_4461)?sg_in116:2'b0)|
    ((_net_469)?sg_in115:2'b0);
   assign  _add_map_x_24_sg_right = ((_net_4462)?sg_in52:2'b0)|
    ((_net_470)?sg_in51:2'b0);
   assign  _add_map_x_24_wall_t_in = dig_w;
   assign  _add_map_x_24_moto = ((_net_4459)?data_in84:10'b0)|
    ((_net_467)?data_in83:10'b0);
   assign  _add_map_x_24_up = ((_net_4458)?data_in83:10'b0)|
    ((_net_466)?data_in84:10'b0);
   assign  _add_map_x_24_right = ((_net_4457)?data_in85:10'b0)|
    ((_net_465)?data_in82:10'b0);
   assign  _add_map_x_24_down = ((_net_4456)?data_in52:10'b0)|
    ((_net_464)?data_in51:10'b0);
   assign  _add_map_x_24_left = ((_net_4455)?data_in116:10'b0)|
    ((_net_463)?data_in115:10'b0);
   assign  _add_map_x_24_start = start;
   assign  _add_map_x_24_goal = goal;
   assign  _add_map_x_24_now = ((_net_4452)?10'b0001010100:10'b0)|
    ((_net_460)?10'b0001010011:10'b0);
   assign  _add_map_x_24_add_exe = (_net_4451|_net_459);
   assign  _add_map_x_24_p_reset = p_reset;
   assign  _add_map_x_24_m_clock = m_clock;
   assign  _add_map_x_23_moto_org_near = ((_net_4450)?data_in_org81:10'b0)|
    ((_net_458)?data_in_org82:10'b0);
   assign  _add_map_x_23_moto_org_near1 = ((_net_4449)?data_in_org83:10'b0)|
    ((_net_457)?data_in_org80:10'b0);
   assign  _add_map_x_23_moto_org_near2 = ((_net_4448)?data_in_org50:10'b0)|
    ((_net_456)?data_in_org49:10'b0);
   assign  _add_map_x_23_moto_org_near3 = ((_net_4447)?data_in_org114:10'b0)|
    ((_net_455)?data_in_org113:10'b0);
   assign  _add_map_x_23_moto_org = ((_net_4446)?data_in_org82:10'b0)|
    ((_net_454)?data_in_org81:10'b0);
   assign  _add_map_x_23_sg_up = ((_net_4445)?sg_in81:2'b0)|
    ((_net_453)?sg_in82:2'b0);
   assign  _add_map_x_23_sg_down = ((_net_4444)?sg_in83:2'b0)|
    ((_net_452)?sg_in80:2'b0);
   assign  _add_map_x_23_sg_left = ((_net_4442)?sg_in114:2'b0)|
    ((_net_450)?sg_in113:2'b0);
   assign  _add_map_x_23_sg_right = ((_net_4443)?sg_in50:2'b0)|
    ((_net_451)?sg_in49:2'b0);
   assign  _add_map_x_23_wall_t_in = dig_w;
   assign  _add_map_x_23_moto = ((_net_4440)?data_in82:10'b0)|
    ((_net_448)?data_in81:10'b0);
   assign  _add_map_x_23_up = ((_net_4439)?data_in81:10'b0)|
    ((_net_447)?data_in82:10'b0);
   assign  _add_map_x_23_right = ((_net_4438)?data_in83:10'b0)|
    ((_net_446)?data_in80:10'b0);
   assign  _add_map_x_23_down = ((_net_4437)?data_in50:10'b0)|
    ((_net_445)?data_in49:10'b0);
   assign  _add_map_x_23_left = ((_net_4436)?data_in114:10'b0)|
    ((_net_444)?data_in113:10'b0);
   assign  _add_map_x_23_start = start;
   assign  _add_map_x_23_goal = goal;
   assign  _add_map_x_23_now = ((_net_4433)?10'b0001010010:10'b0)|
    ((_net_441)?10'b0001010001:10'b0);
   assign  _add_map_x_23_add_exe = (_net_4432|_net_440);
   assign  _add_map_x_23_p_reset = p_reset;
   assign  _add_map_x_23_m_clock = m_clock;
   assign  _add_map_x_22_moto_org_near = ((_net_4431)?data_in_org79:10'b0)|
    ((_net_439)?data_in_org80:10'b0);
   assign  _add_map_x_22_moto_org_near1 = ((_net_4430)?data_in_org81:10'b0)|
    ((_net_438)?data_in_org78:10'b0);
   assign  _add_map_x_22_moto_org_near2 = ((_net_4429)?data_in_org48:10'b0)|
    ((_net_437)?data_in_org47:10'b0);
   assign  _add_map_x_22_moto_org_near3 = ((_net_4428)?data_in_org112:10'b0)|
    ((_net_436)?data_in_org111:10'b0);
   assign  _add_map_x_22_moto_org = ((_net_4427)?data_in_org80:10'b0)|
    ((_net_435)?data_in_org79:10'b0);
   assign  _add_map_x_22_sg_up = ((_net_4426)?sg_in79:2'b0)|
    ((_net_434)?sg_in80:2'b0);
   assign  _add_map_x_22_sg_down = ((_net_4425)?sg_in81:2'b0)|
    ((_net_433)?sg_in78:2'b0);
   assign  _add_map_x_22_sg_left = ((_net_4423)?sg_in112:2'b0)|
    ((_net_431)?sg_in111:2'b0);
   assign  _add_map_x_22_sg_right = ((_net_4424)?sg_in48:2'b0)|
    ((_net_432)?sg_in47:2'b0);
   assign  _add_map_x_22_wall_t_in = dig_w;
   assign  _add_map_x_22_moto = ((_net_4421)?data_in80:10'b0)|
    ((_net_429)?data_in79:10'b0);
   assign  _add_map_x_22_up = ((_net_4420)?data_in79:10'b0)|
    ((_net_428)?data_in80:10'b0);
   assign  _add_map_x_22_right = ((_net_4419)?data_in81:10'b0)|
    ((_net_427)?data_in78:10'b0);
   assign  _add_map_x_22_down = ((_net_4418)?data_in48:10'b0)|
    ((_net_426)?data_in47:10'b0);
   assign  _add_map_x_22_left = ((_net_4417)?data_in112:10'b0)|
    ((_net_425)?data_in111:10'b0);
   assign  _add_map_x_22_start = start;
   assign  _add_map_x_22_goal = goal;
   assign  _add_map_x_22_now = ((_net_4414)?10'b0001010000:10'b0)|
    ((_net_422)?10'b0001001111:10'b0);
   assign  _add_map_x_22_add_exe = (_net_4413|_net_421);
   assign  _add_map_x_22_p_reset = p_reset;
   assign  _add_map_x_22_m_clock = m_clock;
   assign  _add_map_x_21_moto_org_near = ((_net_4412)?data_in_org77:10'b0)|
    ((_net_420)?data_in_org78:10'b0);
   assign  _add_map_x_21_moto_org_near1 = ((_net_4411)?data_in_org79:10'b0)|
    ((_net_419)?data_in_org76:10'b0);
   assign  _add_map_x_21_moto_org_near2 = ((_net_4410)?data_in_org46:10'b0)|
    ((_net_418)?data_in_org45:10'b0);
   assign  _add_map_x_21_moto_org_near3 = ((_net_4409)?data_in_org110:10'b0)|
    ((_net_417)?data_in_org109:10'b0);
   assign  _add_map_x_21_moto_org = ((_net_4408)?data_in_org78:10'b0)|
    ((_net_416)?data_in_org77:10'b0);
   assign  _add_map_x_21_sg_up = ((_net_4407)?sg_in77:2'b0)|
    ((_net_415)?sg_in78:2'b0);
   assign  _add_map_x_21_sg_down = ((_net_4406)?sg_in79:2'b0)|
    ((_net_414)?sg_in76:2'b0);
   assign  _add_map_x_21_sg_left = ((_net_4404)?sg_in110:2'b0)|
    ((_net_412)?sg_in109:2'b0);
   assign  _add_map_x_21_sg_right = ((_net_4405)?sg_in46:2'b0)|
    ((_net_413)?sg_in45:2'b0);
   assign  _add_map_x_21_wall_t_in = dig_w;
   assign  _add_map_x_21_moto = ((_net_4402)?data_in78:10'b0)|
    ((_net_410)?data_in77:10'b0);
   assign  _add_map_x_21_up = ((_net_4401)?data_in77:10'b0)|
    ((_net_409)?data_in78:10'b0);
   assign  _add_map_x_21_right = ((_net_4400)?data_in79:10'b0)|
    ((_net_408)?data_in76:10'b0);
   assign  _add_map_x_21_down = ((_net_4399)?data_in46:10'b0)|
    ((_net_407)?data_in45:10'b0);
   assign  _add_map_x_21_left = ((_net_4398)?data_in110:10'b0)|
    ((_net_406)?data_in109:10'b0);
   assign  _add_map_x_21_start = start;
   assign  _add_map_x_21_goal = goal;
   assign  _add_map_x_21_now = ((_net_4395)?10'b0001001110:10'b0)|
    ((_net_403)?10'b0001001101:10'b0);
   assign  _add_map_x_21_add_exe = (_net_4394|_net_402);
   assign  _add_map_x_21_p_reset = p_reset;
   assign  _add_map_x_21_m_clock = m_clock;
   assign  _add_map_x_20_moto_org_near = ((_net_4393)?data_in_org75:10'b0)|
    ((_net_401)?data_in_org76:10'b0);
   assign  _add_map_x_20_moto_org_near1 = ((_net_4392)?data_in_org77:10'b0)|
    ((_net_400)?data_in_org74:10'b0);
   assign  _add_map_x_20_moto_org_near2 = ((_net_4391)?data_in_org44:10'b0)|
    ((_net_399)?data_in_org43:10'b0);
   assign  _add_map_x_20_moto_org_near3 = ((_net_4390)?data_in_org108:10'b0)|
    ((_net_398)?data_in_org107:10'b0);
   assign  _add_map_x_20_moto_org = ((_net_4389)?data_in_org76:10'b0)|
    ((_net_397)?data_in_org75:10'b0);
   assign  _add_map_x_20_sg_up = ((_net_4388)?sg_in75:2'b0)|
    ((_net_396)?sg_in76:2'b0);
   assign  _add_map_x_20_sg_down = ((_net_4387)?sg_in77:2'b0)|
    ((_net_395)?sg_in74:2'b0);
   assign  _add_map_x_20_sg_left = ((_net_4385)?sg_in108:2'b0)|
    ((_net_393)?sg_in107:2'b0);
   assign  _add_map_x_20_sg_right = ((_net_4386)?sg_in44:2'b0)|
    ((_net_394)?sg_in43:2'b0);
   assign  _add_map_x_20_wall_t_in = dig_w;
   assign  _add_map_x_20_moto = ((_net_4383)?data_in76:10'b0)|
    ((_net_391)?data_in75:10'b0);
   assign  _add_map_x_20_up = ((_net_4382)?data_in75:10'b0)|
    ((_net_390)?data_in76:10'b0);
   assign  _add_map_x_20_right = ((_net_4381)?data_in77:10'b0)|
    ((_net_389)?data_in74:10'b0);
   assign  _add_map_x_20_down = ((_net_4380)?data_in44:10'b0)|
    ((_net_388)?data_in43:10'b0);
   assign  _add_map_x_20_left = ((_net_4379)?data_in108:10'b0)|
    ((_net_387)?data_in107:10'b0);
   assign  _add_map_x_20_start = start;
   assign  _add_map_x_20_goal = goal;
   assign  _add_map_x_20_now = ((_net_4376)?10'b0001001100:10'b0)|
    ((_net_384)?10'b0001001011:10'b0);
   assign  _add_map_x_20_add_exe = (_net_4375|_net_383);
   assign  _add_map_x_20_p_reset = p_reset;
   assign  _add_map_x_20_m_clock = m_clock;
   assign  _add_map_x_19_moto_org_near = ((_net_4374)?data_in_org73:10'b0)|
    ((_net_382)?data_in_org74:10'b0);
   assign  _add_map_x_19_moto_org_near1 = ((_net_4373)?data_in_org75:10'b0)|
    ((_net_381)?data_in_org72:10'b0);
   assign  _add_map_x_19_moto_org_near2 = ((_net_4372)?data_in_org42:10'b0)|
    ((_net_380)?data_in_org41:10'b0);
   assign  _add_map_x_19_moto_org_near3 = ((_net_4371)?data_in_org106:10'b0)|
    ((_net_379)?data_in_org105:10'b0);
   assign  _add_map_x_19_moto_org = ((_net_4370)?data_in_org74:10'b0)|
    ((_net_378)?data_in_org73:10'b0);
   assign  _add_map_x_19_sg_up = ((_net_4369)?sg_in73:2'b0)|
    ((_net_377)?sg_in74:2'b0);
   assign  _add_map_x_19_sg_down = ((_net_4368)?sg_in75:2'b0)|
    ((_net_376)?sg_in72:2'b0);
   assign  _add_map_x_19_sg_left = ((_net_4366)?sg_in106:2'b0)|
    ((_net_374)?sg_in105:2'b0);
   assign  _add_map_x_19_sg_right = ((_net_4367)?sg_in42:2'b0)|
    ((_net_375)?sg_in41:2'b0);
   assign  _add_map_x_19_wall_t_in = dig_w;
   assign  _add_map_x_19_moto = ((_net_4364)?data_in74:10'b0)|
    ((_net_372)?data_in73:10'b0);
   assign  _add_map_x_19_up = ((_net_4363)?data_in73:10'b0)|
    ((_net_371)?data_in74:10'b0);
   assign  _add_map_x_19_right = ((_net_4362)?data_in75:10'b0)|
    ((_net_370)?data_in72:10'b0);
   assign  _add_map_x_19_down = ((_net_4361)?data_in42:10'b0)|
    ((_net_369)?data_in41:10'b0);
   assign  _add_map_x_19_left = ((_net_4360)?data_in106:10'b0)|
    ((_net_368)?data_in105:10'b0);
   assign  _add_map_x_19_start = start;
   assign  _add_map_x_19_goal = goal;
   assign  _add_map_x_19_now = ((_net_4357)?10'b0001001010:10'b0)|
    ((_net_365)?10'b0001001001:10'b0);
   assign  _add_map_x_19_add_exe = (_net_4356|_net_364);
   assign  _add_map_x_19_p_reset = p_reset;
   assign  _add_map_x_19_m_clock = m_clock;
   assign  _add_map_x_18_moto_org_near = ((_net_4355)?data_in_org71:10'b0)|
    ((_net_363)?data_in_org72:10'b0);
   assign  _add_map_x_18_moto_org_near1 = ((_net_4354)?data_in_org73:10'b0)|
    ((_net_362)?data_in_org70:10'b0);
   assign  _add_map_x_18_moto_org_near2 = ((_net_4353)?data_in_org40:10'b0)|
    ((_net_361)?data_in_org39:10'b0);
   assign  _add_map_x_18_moto_org_near3 = ((_net_4352)?data_in_org104:10'b0)|
    ((_net_360)?data_in_org103:10'b0);
   assign  _add_map_x_18_moto_org = ((_net_4351)?data_in_org72:10'b0)|
    ((_net_359)?data_in_org71:10'b0);
   assign  _add_map_x_18_sg_up = ((_net_4350)?sg_in71:2'b0)|
    ((_net_358)?sg_in72:2'b0);
   assign  _add_map_x_18_sg_down = ((_net_4349)?sg_in73:2'b0)|
    ((_net_357)?sg_in70:2'b0);
   assign  _add_map_x_18_sg_left = ((_net_4347)?sg_in104:2'b0)|
    ((_net_355)?sg_in103:2'b0);
   assign  _add_map_x_18_sg_right = ((_net_4348)?sg_in40:2'b0)|
    ((_net_356)?sg_in39:2'b0);
   assign  _add_map_x_18_wall_t_in = dig_w;
   assign  _add_map_x_18_moto = ((_net_4345)?data_in72:10'b0)|
    ((_net_353)?data_in71:10'b0);
   assign  _add_map_x_18_up = ((_net_4344)?data_in71:10'b0)|
    ((_net_352)?data_in72:10'b0);
   assign  _add_map_x_18_right = ((_net_4343)?data_in73:10'b0)|
    ((_net_351)?data_in70:10'b0);
   assign  _add_map_x_18_down = ((_net_4342)?data_in40:10'b0)|
    ((_net_350)?data_in39:10'b0);
   assign  _add_map_x_18_left = ((_net_4341)?data_in104:10'b0)|
    ((_net_349)?data_in103:10'b0);
   assign  _add_map_x_18_start = start;
   assign  _add_map_x_18_goal = goal;
   assign  _add_map_x_18_now = ((_net_4338)?10'b0001001000:10'b0)|
    ((_net_346)?10'b0001000111:10'b0);
   assign  _add_map_x_18_add_exe = (_net_4337|_net_345);
   assign  _add_map_x_18_p_reset = p_reset;
   assign  _add_map_x_18_m_clock = m_clock;
   assign  _add_map_x_17_moto_org_near = ((_net_4336)?data_in_org69:10'b0)|
    ((_net_344)?data_in_org70:10'b0);
   assign  _add_map_x_17_moto_org_near1 = ((_net_4335)?data_in_org71:10'b0)|
    ((_net_343)?data_in_org68:10'b0);
   assign  _add_map_x_17_moto_org_near2 = ((_net_4334)?data_in_org38:10'b0)|
    ((_net_342)?data_in_org37:10'b0);
   assign  _add_map_x_17_moto_org_near3 = ((_net_4333)?data_in_org102:10'b0)|
    ((_net_341)?data_in_org101:10'b0);
   assign  _add_map_x_17_moto_org = ((_net_4332)?data_in_org70:10'b0)|
    ((_net_340)?data_in_org69:10'b0);
   assign  _add_map_x_17_sg_up = ((_net_4331)?sg_in69:2'b0)|
    ((_net_339)?sg_in70:2'b0);
   assign  _add_map_x_17_sg_down = ((_net_4330)?sg_in71:2'b0)|
    ((_net_338)?sg_in68:2'b0);
   assign  _add_map_x_17_sg_left = ((_net_4328)?sg_in102:2'b0)|
    ((_net_336)?sg_in101:2'b0);
   assign  _add_map_x_17_sg_right = ((_net_4329)?sg_in38:2'b0)|
    ((_net_337)?sg_in37:2'b0);
   assign  _add_map_x_17_wall_t_in = dig_w;
   assign  _add_map_x_17_moto = ((_net_4326)?data_in70:10'b0)|
    ((_net_334)?data_in69:10'b0);
   assign  _add_map_x_17_up = ((_net_4325)?data_in69:10'b0)|
    ((_net_333)?data_in70:10'b0);
   assign  _add_map_x_17_right = ((_net_4324)?data_in71:10'b0)|
    ((_net_332)?data_in68:10'b0);
   assign  _add_map_x_17_down = ((_net_4323)?data_in38:10'b0)|
    ((_net_331)?data_in37:10'b0);
   assign  _add_map_x_17_left = ((_net_4322)?data_in102:10'b0)|
    ((_net_330)?data_in101:10'b0);
   assign  _add_map_x_17_start = start;
   assign  _add_map_x_17_goal = goal;
   assign  _add_map_x_17_now = ((_net_4319)?10'b0001000110:10'b0)|
    ((_net_327)?10'b0001000101:10'b0);
   assign  _add_map_x_17_add_exe = (_net_4318|_net_326);
   assign  _add_map_x_17_p_reset = p_reset;
   assign  _add_map_x_17_m_clock = m_clock;
   assign  _add_map_x_16_moto_org_near = ((_net_4317)?data_in_org67:10'b0)|
    ((_net_325)?data_in_org68:10'b0);
   assign  _add_map_x_16_moto_org_near1 = ((_net_4316)?data_in_org69:10'b0)|
    ((_net_324)?data_in_org66:10'b0);
   assign  _add_map_x_16_moto_org_near2 = ((_net_4315)?data_in_org36:10'b0)|
    ((_net_323)?data_in_org35:10'b0);
   assign  _add_map_x_16_moto_org_near3 = ((_net_4314)?data_in_org100:10'b0)|
    ((_net_322)?data_in_org99:10'b0);
   assign  _add_map_x_16_moto_org = ((_net_4313)?data_in_org68:10'b0)|
    ((_net_321)?data_in_org67:10'b0);
   assign  _add_map_x_16_sg_up = ((_net_4312)?sg_in67:2'b0)|
    ((_net_320)?sg_in68:2'b0);
   assign  _add_map_x_16_sg_down = ((_net_4311)?sg_in69:2'b0)|
    ((_net_319)?sg_in66:2'b0);
   assign  _add_map_x_16_sg_left = ((_net_4309)?sg_in100:2'b0)|
    ((_net_317)?sg_in99:2'b0);
   assign  _add_map_x_16_sg_right = ((_net_4310)?sg_in36:2'b0)|
    ((_net_318)?sg_in35:2'b0);
   assign  _add_map_x_16_wall_t_in = dig_w;
   assign  _add_map_x_16_moto = ((_net_4307)?data_in68:10'b0)|
    ((_net_315)?data_in67:10'b0);
   assign  _add_map_x_16_up = ((_net_4306)?data_in67:10'b0)|
    ((_net_314)?data_in68:10'b0);
   assign  _add_map_x_16_right = ((_net_4305)?data_in69:10'b0)|
    ((_net_313)?data_in66:10'b0);
   assign  _add_map_x_16_down = ((_net_4304)?data_in36:10'b0)|
    ((_net_312)?data_in35:10'b0);
   assign  _add_map_x_16_left = ((_net_4303)?data_in100:10'b0)|
    ((_net_311)?data_in99:10'b0);
   assign  _add_map_x_16_start = start;
   assign  _add_map_x_16_goal = goal;
   assign  _add_map_x_16_now = ((_net_4300)?10'b0001000100:10'b0)|
    ((_net_308)?10'b0001000011:10'b0);
   assign  _add_map_x_16_add_exe = (_net_4299|_net_307);
   assign  _add_map_x_16_p_reset = p_reset;
   assign  _add_map_x_16_m_clock = m_clock;
   assign  _add_map_x_15_moto_org_near = ((_net_4298)?data_in_org65:10'b0)|
    ((_net_306)?data_in_org66:10'b0);
   assign  _add_map_x_15_moto_org_near1 = ((_net_4297)?data_in_org67:10'b0)|
    ((_net_305)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_15_moto_org_near2 = ((_net_4296)?data_in_org34:10'b0)|
    ((_net_304)?data_in_org33:10'b0);
   assign  _add_map_x_15_moto_org_near3 = ((_net_4295)?data_in_org98:10'b0)|
    ((_net_303)?data_in_org97:10'b0);
   assign  _add_map_x_15_moto_org = ((_net_4294)?data_in_org66:10'b0)|
    ((_net_302)?data_in_org65:10'b0);
   assign  _add_map_x_15_sg_up = ((_net_4293)?sg_in65:2'b0)|
    ((_net_301)?sg_in66:2'b0);
   assign  _add_map_x_15_sg_down = ((_net_4292)?sg_in67:2'b0)|
    ((_net_300)?3'b000:2'b0);
   assign  _add_map_x_15_sg_left = ((_net_4290)?sg_in98:2'b0)|
    ((_net_298)?sg_in97:2'b0);
   assign  _add_map_x_15_sg_right = ((_net_4291)?sg_in34:2'b0)|
    ((_net_299)?sg_in33:2'b0);
   assign  _add_map_x_15_wall_t_in = dig_w;
   assign  _add_map_x_15_moto = ((_net_4288)?data_in66:10'b0)|
    ((_net_296)?data_in65:10'b0);
   assign  _add_map_x_15_up = ((_net_4287)?data_in65:10'b0)|
    ((_net_295)?data_in66:10'b0);
   assign  _add_map_x_15_right = ((_net_4286)?data_in67:10'b0)|
    ((_net_294)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_15_down = ((_net_4285)?data_in34:10'b0)|
    ((_net_293)?data_in33:10'b0);
   assign  _add_map_x_15_left = ((_net_4284)?data_in98:10'b0)|
    ((_net_292)?data_in97:10'b0);
   assign  _add_map_x_15_start = start;
   assign  _add_map_x_15_goal = goal;
   assign  _add_map_x_15_now = ((_net_4281)?10'b0001000010:10'b0)|
    ((_net_289)?10'b0001000001:10'b0);
   assign  _add_map_x_15_add_exe = (_net_4280|_net_288);
   assign  _add_map_x_15_p_reset = p_reset;
   assign  _add_map_x_15_m_clock = m_clock;
   assign  _add_map_x_14_moto_org_near = ((_net_4279)?data_in_org62:10'b0)|
    ((_net_287)?data_in_org61:10'b0);
   assign  _add_map_x_14_moto_org_near1 = ((_net_4278)?data_in_org60:10'b0)|
    ((_net_286)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_14_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_14_moto_org_near3 = ((_net_4276)?data_in_org93:10'b0)|
    ((_net_284)?data_in_org94:10'b0);
   assign  _add_map_x_14_moto_org = ((_net_4275)?data_in_org61:10'b0)|
    ((_net_283)?data_in_org62:10'b0);
   assign  _add_map_x_14_sg_up = ((_net_4274)?sg_in62:2'b0)|
    ((_net_282)?sg_in61:2'b0);
   assign  _add_map_x_14_sg_down = 3'b000;
   assign  _add_map_x_14_sg_left = ((_net_4271)?sg_in93:2'b0)|
    ((_net_279)?sg_in94:2'b0);
   assign  _add_map_x_14_sg_right = ((_net_4272)?sg_in60:2'b0)|
    ((_net_280)?3'b000:2'b0);
   assign  _add_map_x_14_wall_t_in = dig_w;
   assign  _add_map_x_14_moto = ((_net_4269)?data_in61:10'b0)|
    ((_net_277)?data_in62:10'b0);
   assign  _add_map_x_14_up = ((_net_4268)?data_in62:10'b0)|
    ((_net_276)?data_in61:10'b0);
   assign  _add_map_x_14_right = ((_net_4267)?data_in60:10'b0)|
    ((_net_275)?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):10'b0);
   assign  _add_map_x_14_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_14_left = ((_net_4265)?data_in93:10'b0)|
    ((_net_273)?data_in94:10'b0);
   assign  _add_map_x_14_start = start;
   assign  _add_map_x_14_goal = goal;
   assign  _add_map_x_14_now = ((_net_4262)?10'b0000111101:10'b0)|
    ((_net_270)?10'b0000111110:10'b0);
   assign  _add_map_x_14_add_exe = (_net_4261|_net_269);
   assign  _add_map_x_14_p_reset = p_reset;
   assign  _add_map_x_14_m_clock = m_clock;
   assign  _add_map_x_13_moto_org_near = ((_net_4260)?data_in_org60:10'b0)|
    ((_net_268)?data_in_org59:10'b0);
   assign  _add_map_x_13_moto_org_near1 = ((_net_4259)?data_in_org58:10'b0)|
    ((_net_267)?data_in_org61:10'b0);
   assign  _add_map_x_13_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_13_moto_org_near3 = ((_net_4257)?data_in_org91:10'b0)|
    ((_net_265)?data_in_org92:10'b0);
   assign  _add_map_x_13_moto_org = ((_net_4256)?data_in_org59:10'b0)|
    ((_net_264)?data_in_org60:10'b0);
   assign  _add_map_x_13_sg_up = ((_net_4255)?sg_in60:2'b0)|
    ((_net_263)?sg_in59:2'b0);
   assign  _add_map_x_13_sg_down = ((_net_4254)?3'b000:2'b0)|
    ((_net_262)?sg_in61:2'b0);
   assign  _add_map_x_13_sg_left = ((_net_4252)?sg_in91:2'b0)|
    ((_net_260)?sg_in92:2'b0);
   assign  _add_map_x_13_sg_right = ((_net_4253)?sg_in58:2'b0)|
    ((_net_261)?3'b000:2'b0);
   assign  _add_map_x_13_wall_t_in = dig_w;
   assign  _add_map_x_13_moto = ((_net_4250)?data_in59:10'b0)|
    ((_net_258)?data_in60:10'b0);
   assign  _add_map_x_13_up = ((_net_4249)?data_in60:10'b0)|
    ((_net_257)?data_in59:10'b0);
   assign  _add_map_x_13_right = ((_net_4248)?data_in58:10'b0)|
    ((_net_256)?data_in61:10'b0);
   assign  _add_map_x_13_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_13_left = ((_net_4246)?data_in91:10'b0)|
    ((_net_254)?data_in92:10'b0);
   assign  _add_map_x_13_start = start;
   assign  _add_map_x_13_goal = goal;
   assign  _add_map_x_13_now = ((_net_4243)?10'b0000111011:10'b0)|
    ((_net_251)?10'b0000111100:10'b0);
   assign  _add_map_x_13_add_exe = (_net_4242|_net_250);
   assign  _add_map_x_13_p_reset = p_reset;
   assign  _add_map_x_13_m_clock = m_clock;
   assign  _add_map_x_12_moto_org_near = ((_net_4241)?data_in_org58:10'b0)|
    ((_net_249)?data_in_org57:10'b0);
   assign  _add_map_x_12_moto_org_near1 = ((_net_4240)?data_in_org56:10'b0)|
    ((_net_248)?data_in_org59:10'b0);
   assign  _add_map_x_12_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_12_moto_org_near3 = ((_net_4238)?data_in_org89:10'b0)|
    ((_net_246)?data_in_org90:10'b0);
   assign  _add_map_x_12_moto_org = ((_net_4237)?data_in_org57:10'b0)|
    ((_net_245)?data_in_org58:10'b0);
   assign  _add_map_x_12_sg_up = ((_net_4236)?sg_in58:2'b0)|
    ((_net_244)?sg_in57:2'b0);
   assign  _add_map_x_12_sg_down = ((_net_4235)?3'b000:2'b0)|
    ((_net_243)?sg_in59:2'b0);
   assign  _add_map_x_12_sg_left = ((_net_4233)?sg_in89:2'b0)|
    ((_net_241)?sg_in90:2'b0);
   assign  _add_map_x_12_sg_right = ((_net_4234)?sg_in56:2'b0)|
    ((_net_242)?3'b000:2'b0);
   assign  _add_map_x_12_wall_t_in = dig_w;
   assign  _add_map_x_12_moto = ((_net_4231)?data_in57:10'b0)|
    ((_net_239)?data_in58:10'b0);
   assign  _add_map_x_12_up = ((_net_4230)?data_in58:10'b0)|
    ((_net_238)?data_in57:10'b0);
   assign  _add_map_x_12_right = ((_net_4229)?data_in56:10'b0)|
    ((_net_237)?data_in59:10'b0);
   assign  _add_map_x_12_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_12_left = ((_net_4227)?data_in89:10'b0)|
    ((_net_235)?data_in90:10'b0);
   assign  _add_map_x_12_start = start;
   assign  _add_map_x_12_goal = goal;
   assign  _add_map_x_12_now = ((_net_4224)?10'b0000111001:10'b0)|
    ((_net_232)?10'b0000111010:10'b0);
   assign  _add_map_x_12_add_exe = (_net_4223|_net_231);
   assign  _add_map_x_12_p_reset = p_reset;
   assign  _add_map_x_12_m_clock = m_clock;
   assign  _add_map_x_11_moto_org_near = ((_net_4222)?data_in_org56:10'b0)|
    ((_net_230)?data_in_org55:10'b0);
   assign  _add_map_x_11_moto_org_near1 = ((_net_4221)?data_in_org54:10'b0)|
    ((_net_229)?data_in_org57:10'b0);
   assign  _add_map_x_11_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_11_moto_org_near3 = ((_net_4219)?data_in_org87:10'b0)|
    ((_net_227)?data_in_org88:10'b0);
   assign  _add_map_x_11_moto_org = ((_net_4218)?data_in_org55:10'b0)|
    ((_net_226)?data_in_org56:10'b0);
   assign  _add_map_x_11_sg_up = ((_net_4217)?sg_in56:2'b0)|
    ((_net_225)?sg_in55:2'b0);
   assign  _add_map_x_11_sg_down = ((_net_4216)?3'b000:2'b0)|
    ((_net_224)?sg_in57:2'b0);
   assign  _add_map_x_11_sg_left = ((_net_4214)?sg_in87:2'b0)|
    ((_net_222)?sg_in88:2'b0);
   assign  _add_map_x_11_sg_right = ((_net_4215)?sg_in54:2'b0)|
    ((_net_223)?3'b000:2'b0);
   assign  _add_map_x_11_wall_t_in = dig_w;
   assign  _add_map_x_11_moto = ((_net_4212)?data_in55:10'b0)|
    ((_net_220)?data_in56:10'b0);
   assign  _add_map_x_11_up = ((_net_4211)?data_in56:10'b0)|
    ((_net_219)?data_in55:10'b0);
   assign  _add_map_x_11_right = ((_net_4210)?data_in54:10'b0)|
    ((_net_218)?data_in57:10'b0);
   assign  _add_map_x_11_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_11_left = ((_net_4208)?data_in87:10'b0)|
    ((_net_216)?data_in88:10'b0);
   assign  _add_map_x_11_start = start;
   assign  _add_map_x_11_goal = goal;
   assign  _add_map_x_11_now = ((_net_4205)?10'b0000110111:10'b0)|
    ((_net_213)?10'b0000111000:10'b0);
   assign  _add_map_x_11_add_exe = (_net_4204|_net_212);
   assign  _add_map_x_11_p_reset = p_reset;
   assign  _add_map_x_11_m_clock = m_clock;
   assign  _add_map_x_10_moto_org_near = ((_net_4203)?data_in_org54:10'b0)|
    ((_net_211)?data_in_org53:10'b0);
   assign  _add_map_x_10_moto_org_near1 = ((_net_4202)?data_in_org52:10'b0)|
    ((_net_210)?data_in_org55:10'b0);
   assign  _add_map_x_10_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_10_moto_org_near3 = ((_net_4200)?data_in_org85:10'b0)|
    ((_net_208)?data_in_org86:10'b0);
   assign  _add_map_x_10_moto_org = ((_net_4199)?data_in_org53:10'b0)|
    ((_net_207)?data_in_org54:10'b0);
   assign  _add_map_x_10_sg_up = ((_net_4198)?sg_in54:2'b0)|
    ((_net_206)?sg_in53:2'b0);
   assign  _add_map_x_10_sg_down = ((_net_4197)?3'b000:2'b0)|
    ((_net_205)?sg_in55:2'b0);
   assign  _add_map_x_10_sg_left = ((_net_4195)?sg_in85:2'b0)|
    ((_net_203)?sg_in86:2'b0);
   assign  _add_map_x_10_sg_right = ((_net_4196)?sg_in52:2'b0)|
    ((_net_204)?3'b000:2'b0);
   assign  _add_map_x_10_wall_t_in = dig_w;
   assign  _add_map_x_10_moto = ((_net_4193)?data_in53:10'b0)|
    ((_net_201)?data_in54:10'b0);
   assign  _add_map_x_10_up = ((_net_4192)?data_in54:10'b0)|
    ((_net_200)?data_in53:10'b0);
   assign  _add_map_x_10_right = ((_net_4191)?data_in52:10'b0)|
    ((_net_199)?data_in55:10'b0);
   assign  _add_map_x_10_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_10_left = ((_net_4189)?data_in85:10'b0)|
    ((_net_197)?data_in86:10'b0);
   assign  _add_map_x_10_start = start;
   assign  _add_map_x_10_goal = goal;
   assign  _add_map_x_10_now = ((_net_4186)?10'b0000110101:10'b0)|
    ((_net_194)?10'b0000110110:10'b0);
   assign  _add_map_x_10_add_exe = (_net_4185|_net_193);
   assign  _add_map_x_10_p_reset = p_reset;
   assign  _add_map_x_10_m_clock = m_clock;
   assign  _add_map_x_9_moto_org_near = ((_net_4184)?data_in_org52:10'b0)|
    ((_net_192)?data_in_org51:10'b0);
   assign  _add_map_x_9_moto_org_near1 = ((_net_4183)?data_in_org50:10'b0)|
    ((_net_191)?data_in_org53:10'b0);
   assign  _add_map_x_9_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_9_moto_org_near3 = ((_net_4181)?data_in_org83:10'b0)|
    ((_net_189)?data_in_org84:10'b0);
   assign  _add_map_x_9_moto_org = ((_net_4180)?data_in_org51:10'b0)|
    ((_net_188)?data_in_org52:10'b0);
   assign  _add_map_x_9_sg_up = ((_net_4179)?sg_in52:2'b0)|
    ((_net_187)?sg_in51:2'b0);
   assign  _add_map_x_9_sg_down = ((_net_4178)?3'b000:2'b0)|
    ((_net_186)?sg_in53:2'b0);
   assign  _add_map_x_9_sg_left = ((_net_4176)?sg_in83:2'b0)|
    ((_net_184)?sg_in84:2'b0);
   assign  _add_map_x_9_sg_right = ((_net_4177)?sg_in50:2'b0)|
    ((_net_185)?3'b000:2'b0);
   assign  _add_map_x_9_wall_t_in = dig_w;
   assign  _add_map_x_9_moto = ((_net_4174)?data_in51:10'b0)|
    ((_net_182)?data_in52:10'b0);
   assign  _add_map_x_9_up = ((_net_4173)?data_in52:10'b0)|
    ((_net_181)?data_in51:10'b0);
   assign  _add_map_x_9_right = ((_net_4172)?data_in50:10'b0)|
    ((_net_180)?data_in53:10'b0);
   assign  _add_map_x_9_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_9_left = ((_net_4170)?data_in83:10'b0)|
    ((_net_178)?data_in84:10'b0);
   assign  _add_map_x_9_start = start;
   assign  _add_map_x_9_goal = goal;
   assign  _add_map_x_9_now = ((_net_4167)?10'b0000110011:10'b0)|
    ((_net_175)?10'b0000110100:10'b0);
   assign  _add_map_x_9_add_exe = (_net_4166|_net_174);
   assign  _add_map_x_9_p_reset = p_reset;
   assign  _add_map_x_9_m_clock = m_clock;
   assign  _add_map_x_8_moto_org_near = ((_net_4165)?data_in_org50:10'b0)|
    ((_net_173)?data_in_org49:10'b0);
   assign  _add_map_x_8_moto_org_near1 = ((_net_4164)?data_in_org48:10'b0)|
    ((_net_172)?data_in_org51:10'b0);
   assign  _add_map_x_8_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_8_moto_org_near3 = ((_net_4162)?data_in_org81:10'b0)|
    ((_net_170)?data_in_org82:10'b0);
   assign  _add_map_x_8_moto_org = ((_net_4161)?data_in_org49:10'b0)|
    ((_net_169)?data_in_org50:10'b0);
   assign  _add_map_x_8_sg_up = ((_net_4160)?sg_in50:2'b0)|
    ((_net_168)?sg_in49:2'b0);
   assign  _add_map_x_8_sg_down = ((_net_4159)?3'b000:2'b0)|
    ((_net_167)?sg_in51:2'b0);
   assign  _add_map_x_8_sg_left = ((_net_4157)?sg_in81:2'b0)|
    ((_net_165)?sg_in82:2'b0);
   assign  _add_map_x_8_sg_right = ((_net_4158)?sg_in48:2'b0)|
    ((_net_166)?3'b000:2'b0);
   assign  _add_map_x_8_wall_t_in = dig_w;
   assign  _add_map_x_8_moto = ((_net_4155)?data_in49:10'b0)|
    ((_net_163)?data_in50:10'b0);
   assign  _add_map_x_8_up = ((_net_4154)?data_in50:10'b0)|
    ((_net_162)?data_in49:10'b0);
   assign  _add_map_x_8_right = ((_net_4153)?data_in48:10'b0)|
    ((_net_161)?data_in51:10'b0);
   assign  _add_map_x_8_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_8_left = ((_net_4151)?data_in81:10'b0)|
    ((_net_159)?data_in82:10'b0);
   assign  _add_map_x_8_start = start;
   assign  _add_map_x_8_goal = goal;
   assign  _add_map_x_8_now = ((_net_4148)?10'b0000110001:10'b0)|
    ((_net_156)?10'b0000110010:10'b0);
   assign  _add_map_x_8_add_exe = (_net_4147|_net_155);
   assign  _add_map_x_8_p_reset = p_reset;
   assign  _add_map_x_8_m_clock = m_clock;
   assign  _add_map_x_7_moto_org_near = ((_net_4146)?data_in_org48:10'b0)|
    ((_net_154)?data_in_org47:10'b0);
   assign  _add_map_x_7_moto_org_near1 = ((_net_4145)?data_in_org46:10'b0)|
    ((_net_153)?data_in_org49:10'b0);
   assign  _add_map_x_7_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_7_moto_org_near3 = ((_net_4143)?data_in_org79:10'b0)|
    ((_net_151)?data_in_org80:10'b0);
   assign  _add_map_x_7_moto_org = ((_net_4142)?data_in_org47:10'b0)|
    ((_net_150)?data_in_org48:10'b0);
   assign  _add_map_x_7_sg_up = ((_net_4141)?sg_in48:2'b0)|
    ((_net_149)?sg_in47:2'b0);
   assign  _add_map_x_7_sg_down = ((_net_4140)?3'b000:2'b0)|
    ((_net_148)?sg_in49:2'b0);
   assign  _add_map_x_7_sg_left = ((_net_4138)?sg_in79:2'b0)|
    ((_net_146)?sg_in80:2'b0);
   assign  _add_map_x_7_sg_right = ((_net_4139)?sg_in46:2'b0)|
    ((_net_147)?3'b000:2'b0);
   assign  _add_map_x_7_wall_t_in = dig_w;
   assign  _add_map_x_7_moto = ((_net_4136)?data_in47:10'b0)|
    ((_net_144)?data_in48:10'b0);
   assign  _add_map_x_7_up = ((_net_4135)?data_in48:10'b0)|
    ((_net_143)?data_in47:10'b0);
   assign  _add_map_x_7_right = ((_net_4134)?data_in46:10'b0)|
    ((_net_142)?data_in49:10'b0);
   assign  _add_map_x_7_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_7_left = ((_net_4132)?data_in79:10'b0)|
    ((_net_140)?data_in80:10'b0);
   assign  _add_map_x_7_start = start;
   assign  _add_map_x_7_goal = goal;
   assign  _add_map_x_7_now = ((_net_4129)?10'b0000101111:10'b0)|
    ((_net_137)?10'b0000110000:10'b0);
   assign  _add_map_x_7_add_exe = (_net_4128|_net_136);
   assign  _add_map_x_7_p_reset = p_reset;
   assign  _add_map_x_7_m_clock = m_clock;
   assign  _add_map_x_6_moto_org_near = ((_net_4127)?data_in_org46:10'b0)|
    ((_net_135)?data_in_org45:10'b0);
   assign  _add_map_x_6_moto_org_near1 = ((_net_4126)?data_in_org44:10'b0)|
    ((_net_134)?data_in_org47:10'b0);
   assign  _add_map_x_6_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_6_moto_org_near3 = ((_net_4124)?data_in_org77:10'b0)|
    ((_net_132)?data_in_org78:10'b0);
   assign  _add_map_x_6_moto_org = ((_net_4123)?data_in_org45:10'b0)|
    ((_net_131)?data_in_org46:10'b0);
   assign  _add_map_x_6_sg_up = ((_net_4122)?sg_in46:2'b0)|
    ((_net_130)?sg_in45:2'b0);
   assign  _add_map_x_6_sg_down = ((_net_4121)?3'b000:2'b0)|
    ((_net_129)?sg_in47:2'b0);
   assign  _add_map_x_6_sg_left = ((_net_4119)?sg_in77:2'b0)|
    ((_net_127)?sg_in78:2'b0);
   assign  _add_map_x_6_sg_right = ((_net_4120)?sg_in44:2'b0)|
    ((_net_128)?3'b000:2'b0);
   assign  _add_map_x_6_wall_t_in = dig_w;
   assign  _add_map_x_6_moto = ((_net_4117)?data_in45:10'b0)|
    ((_net_125)?data_in46:10'b0);
   assign  _add_map_x_6_up = ((_net_4116)?data_in46:10'b0)|
    ((_net_124)?data_in45:10'b0);
   assign  _add_map_x_6_right = ((_net_4115)?data_in44:10'b0)|
    ((_net_123)?data_in47:10'b0);
   assign  _add_map_x_6_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_6_left = ((_net_4113)?data_in77:10'b0)|
    ((_net_121)?data_in78:10'b0);
   assign  _add_map_x_6_start = start;
   assign  _add_map_x_6_goal = goal;
   assign  _add_map_x_6_now = ((_net_4110)?10'b0000101101:10'b0)|
    ((_net_118)?10'b0000101110:10'b0);
   assign  _add_map_x_6_add_exe = (_net_4109|_net_117);
   assign  _add_map_x_6_p_reset = p_reset;
   assign  _add_map_x_6_m_clock = m_clock;
   assign  _add_map_x_5_moto_org_near = ((_net_4108)?data_in_org44:10'b0)|
    ((_net_116)?data_in_org43:10'b0);
   assign  _add_map_x_5_moto_org_near1 = ((_net_4107)?data_in_org42:10'b0)|
    ((_net_115)?data_in_org45:10'b0);
   assign  _add_map_x_5_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_5_moto_org_near3 = ((_net_4105)?data_in_org75:10'b0)|
    ((_net_113)?data_in_org76:10'b0);
   assign  _add_map_x_5_moto_org = ((_net_4104)?data_in_org43:10'b0)|
    ((_net_112)?data_in_org44:10'b0);
   assign  _add_map_x_5_sg_up = ((_net_4103)?sg_in44:2'b0)|
    ((_net_111)?sg_in43:2'b0);
   assign  _add_map_x_5_sg_down = ((_net_4102)?3'b000:2'b0)|
    ((_net_110)?sg_in45:2'b0);
   assign  _add_map_x_5_sg_left = ((_net_4100)?sg_in75:2'b0)|
    ((_net_108)?sg_in76:2'b0);
   assign  _add_map_x_5_sg_right = ((_net_4101)?sg_in42:2'b0)|
    ((_net_109)?3'b000:2'b0);
   assign  _add_map_x_5_wall_t_in = dig_w;
   assign  _add_map_x_5_moto = ((_net_4098)?data_in43:10'b0)|
    ((_net_106)?data_in44:10'b0);
   assign  _add_map_x_5_up = ((_net_4097)?data_in44:10'b0)|
    ((_net_105)?data_in43:10'b0);
   assign  _add_map_x_5_right = ((_net_4096)?data_in42:10'b0)|
    ((_net_104)?data_in45:10'b0);
   assign  _add_map_x_5_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_5_left = ((_net_4094)?data_in75:10'b0)|
    ((_net_102)?data_in76:10'b0);
   assign  _add_map_x_5_start = start;
   assign  _add_map_x_5_goal = goal;
   assign  _add_map_x_5_now = ((_net_4091)?10'b0000101011:10'b0)|
    ((_net_99)?10'b0000101100:10'b0);
   assign  _add_map_x_5_add_exe = (_net_4090|_net_98);
   assign  _add_map_x_5_p_reset = p_reset;
   assign  _add_map_x_5_m_clock = m_clock;
   assign  _add_map_x_4_moto_org_near = ((_net_4089)?data_in_org42:10'b0)|
    ((_net_97)?data_in_org41:10'b0);
   assign  _add_map_x_4_moto_org_near1 = ((_net_4088)?data_in_org40:10'b0)|
    ((_net_96)?data_in_org43:10'b0);
   assign  _add_map_x_4_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_4_moto_org_near3 = ((_net_4086)?data_in_org73:10'b0)|
    ((_net_94)?data_in_org74:10'b0);
   assign  _add_map_x_4_moto_org = ((_net_4085)?data_in_org41:10'b0)|
    ((_net_93)?data_in_org42:10'b0);
   assign  _add_map_x_4_sg_up = ((_net_4084)?sg_in42:2'b0)|
    ((_net_92)?sg_in41:2'b0);
   assign  _add_map_x_4_sg_down = ((_net_4083)?3'b000:2'b0)|
    ((_net_91)?sg_in43:2'b0);
   assign  _add_map_x_4_sg_left = ((_net_4081)?sg_in73:2'b0)|
    ((_net_89)?sg_in74:2'b0);
   assign  _add_map_x_4_sg_right = ((_net_4082)?sg_in40:2'b0)|
    ((_net_90)?3'b000:2'b0);
   assign  _add_map_x_4_wall_t_in = dig_w;
   assign  _add_map_x_4_moto = ((_net_4079)?data_in41:10'b0)|
    ((_net_87)?data_in42:10'b0);
   assign  _add_map_x_4_up = ((_net_4078)?data_in42:10'b0)|
    ((_net_86)?data_in41:10'b0);
   assign  _add_map_x_4_right = ((_net_4077)?data_in40:10'b0)|
    ((_net_85)?data_in43:10'b0);
   assign  _add_map_x_4_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_4_left = ((_net_4075)?data_in73:10'b0)|
    ((_net_83)?data_in74:10'b0);
   assign  _add_map_x_4_start = start;
   assign  _add_map_x_4_goal = goal;
   assign  _add_map_x_4_now = ((_net_4072)?10'b0000101001:10'b0)|
    ((_net_80)?10'b0000101010:10'b0);
   assign  _add_map_x_4_add_exe = (_net_4071|_net_79);
   assign  _add_map_x_4_p_reset = p_reset;
   assign  _add_map_x_4_m_clock = m_clock;
   assign  _add_map_x_3_moto_org_near = ((_net_4070)?data_in_org40:10'b0)|
    ((_net_78)?data_in_org39:10'b0);
   assign  _add_map_x_3_moto_org_near1 = ((_net_4069)?data_in_org38:10'b0)|
    ((_net_77)?data_in_org41:10'b0);
   assign  _add_map_x_3_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_3_moto_org_near3 = ((_net_4067)?data_in_org71:10'b0)|
    ((_net_75)?data_in_org72:10'b0);
   assign  _add_map_x_3_moto_org = ((_net_4066)?data_in_org39:10'b0)|
    ((_net_74)?data_in_org40:10'b0);
   assign  _add_map_x_3_sg_up = ((_net_4065)?sg_in40:2'b0)|
    ((_net_73)?sg_in39:2'b0);
   assign  _add_map_x_3_sg_down = ((_net_4064)?3'b000:2'b0)|
    ((_net_72)?sg_in41:2'b0);
   assign  _add_map_x_3_sg_left = ((_net_4062)?sg_in71:2'b0)|
    ((_net_70)?sg_in72:2'b0);
   assign  _add_map_x_3_sg_right = ((_net_4063)?sg_in38:2'b0)|
    ((_net_71)?3'b000:2'b0);
   assign  _add_map_x_3_wall_t_in = dig_w;
   assign  _add_map_x_3_moto = ((_net_4060)?data_in39:10'b0)|
    ((_net_68)?data_in40:10'b0);
   assign  _add_map_x_3_up = ((_net_4059)?data_in40:10'b0)|
    ((_net_67)?data_in39:10'b0);
   assign  _add_map_x_3_right = ((_net_4058)?data_in38:10'b0)|
    ((_net_66)?data_in41:10'b0);
   assign  _add_map_x_3_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_3_left = ((_net_4056)?data_in71:10'b0)|
    ((_net_64)?data_in72:10'b0);
   assign  _add_map_x_3_start = start;
   assign  _add_map_x_3_goal = goal;
   assign  _add_map_x_3_now = ((_net_4053)?10'b0000100111:10'b0)|
    ((_net_61)?10'b0000101000:10'b0);
   assign  _add_map_x_3_add_exe = (_net_4052|_net_60);
   assign  _add_map_x_3_p_reset = p_reset;
   assign  _add_map_x_3_m_clock = m_clock;
   assign  _add_map_x_2_moto_org_near = ((_net_4051)?data_in_org38:10'b0)|
    ((_net_59)?data_in_org37:10'b0);
   assign  _add_map_x_2_moto_org_near1 = ((_net_4050)?data_in_org36:10'b0)|
    ((_net_58)?data_in_org39:10'b0);
   assign  _add_map_x_2_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_2_moto_org_near3 = ((_net_4048)?data_in_org69:10'b0)|
    ((_net_56)?data_in_org70:10'b0);
   assign  _add_map_x_2_moto_org = ((_net_4047)?data_in_org37:10'b0)|
    ((_net_55)?data_in_org38:10'b0);
   assign  _add_map_x_2_sg_up = ((_net_4046)?sg_in38:2'b0)|
    ((_net_54)?sg_in37:2'b0);
   assign  _add_map_x_2_sg_down = ((_net_4045)?3'b000:2'b0)|
    ((_net_53)?sg_in39:2'b0);
   assign  _add_map_x_2_sg_left = ((_net_4043)?sg_in69:2'b0)|
    ((_net_51)?sg_in70:2'b0);
   assign  _add_map_x_2_sg_right = ((_net_4044)?sg_in36:2'b0)|
    ((_net_52)?3'b000:2'b0);
   assign  _add_map_x_2_wall_t_in = dig_w;
   assign  _add_map_x_2_moto = ((_net_4041)?data_in37:10'b0)|
    ((_net_49)?data_in38:10'b0);
   assign  _add_map_x_2_up = ((_net_4040)?data_in38:10'b0)|
    ((_net_48)?data_in37:10'b0);
   assign  _add_map_x_2_right = ((_net_4039)?data_in36:10'b0)|
    ((_net_47)?data_in39:10'b0);
   assign  _add_map_x_2_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_2_left = ((_net_4037)?data_in69:10'b0)|
    ((_net_45)?data_in70:10'b0);
   assign  _add_map_x_2_start = start;
   assign  _add_map_x_2_goal = goal;
   assign  _add_map_x_2_now = ((_net_4034)?10'b0000100101:10'b0)|
    ((_net_42)?10'b0000100110:10'b0);
   assign  _add_map_x_2_add_exe = (_net_4033|_net_41);
   assign  _add_map_x_2_p_reset = p_reset;
   assign  _add_map_x_2_m_clock = m_clock;
   assign  _add_map_x_1_moto_org_near = ((_net_4032)?data_in_org36:10'b0)|
    ((_net_40)?data_in_org35:10'b0);
   assign  _add_map_x_1_moto_org_near1 = ((_net_4031)?data_in_org34:10'b0)|
    ((_net_39)?data_in_org37:10'b0);
   assign  _add_map_x_1_moto_org_near2 = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_1_moto_org_near3 = ((_net_4029)?data_in_org67:10'b0)|
    ((_net_37)?data_in_org68:10'b0);
   assign  _add_map_x_1_moto_org = ((_net_4028)?data_in_org35:10'b0)|
    ((_net_36)?data_in_org36:10'b0);
   assign  _add_map_x_1_sg_up = ((_net_4027)?sg_in36:2'b0)|
    ((_net_35)?sg_in35:2'b0);
   assign  _add_map_x_1_sg_down = ((_net_4026)?3'b000:2'b0)|
    ((_net_34)?sg_in37:2'b0);
   assign  _add_map_x_1_sg_left = ((_net_4024)?sg_in67:2'b0)|
    ((_net_32)?sg_in68:2'b0);
   assign  _add_map_x_1_sg_right = ((_net_4025)?sg_in34:2'b0)|
    ((_net_33)?3'b000:2'b0);
   assign  _add_map_x_1_wall_t_in = dig_w;
   assign  _add_map_x_1_moto = ((_net_4022)?data_in35:10'b0)|
    ((_net_30)?data_in36:10'b0);
   assign  _add_map_x_1_up = ((_net_4021)?data_in36:10'b0)|
    ((_net_29)?data_in35:10'b0);
   assign  _add_map_x_1_right = ((_net_4020)?data_in34:10'b0)|
    ((_net_28)?data_in37:10'b0);
   assign  _add_map_x_1_down = ({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1});
   assign  _add_map_x_1_left = ((_net_4018)?data_in67:10'b0)|
    ((_net_26)?data_in68:10'b0);
   assign  _add_map_x_1_start = start;
   assign  _add_map_x_1_goal = goal;
   assign  _add_map_x_1_now = ((_net_4015)?10'b0000100011:10'b0)|
    ((_net_23)?10'b0000100100:10'b0);
   assign  _add_map_x_1_add_exe = (_net_4014|_net_22);
   assign  _add_map_x_1_p_reset = p_reset;
   assign  _add_map_x_1_m_clock = m_clock;
   assign  _net_0 = (sig_reg==1'b0);
   assign  _net_1 = (sig_reg==1'b1);
   assign  _net_2 = (sig==1'b1);
   assign  _net_3 = (in_do&_net_2);
   assign  _net_4 = (in_do&_net_2);
   assign  _net_5 = (in_do&_net_2);
   assign  _net_6 = (in_do&_net_2);
   assign  _net_7 = (in_do&_net_2);
   assign  _net_8 = (in_do&_net_2);
   assign  _net_9 = (in_do&_net_2);
   assign  _net_10 = (in_do&_net_2);
   assign  _net_11 = (in_do&_net_2);
   assign  _net_12 = (in_do&_net_2);
   assign  _net_13 = (in_do&_net_2);
   assign  _net_14 = (in_do&_net_2);
   assign  _net_15 = (in_do&_net_2);
   assign  _net_16 = (in_do&_net_2);
   assign  _net_17 = (in_do&_net_2);
   assign  _net_18 = (in_do&_net_2);
   assign  _net_19 = (in_do&_net_2);
   assign  _net_20 = (in_do&_net_2);
   assign  _net_21 = (in_do&_net_2);
   assign  _net_22 = (in_do&_net_2);
   assign  _net_23 = (in_do&_net_2);
   assign  _net_24 = (in_do&_net_2);
   assign  _net_25 = (in_do&_net_2);
   assign  _net_26 = (in_do&_net_2);
   assign  _net_27 = (in_do&_net_2);
   assign  _net_28 = (in_do&_net_2);
   assign  _net_29 = (in_do&_net_2);
   assign  _net_30 = (in_do&_net_2);
   assign  _net_31 = (in_do&_net_2);
   assign  _net_32 = (in_do&_net_2);
   assign  _net_33 = (in_do&_net_2);
   assign  _net_34 = (in_do&_net_2);
   assign  _net_35 = (in_do&_net_2);
   assign  _net_36 = (in_do&_net_2);
   assign  _net_37 = (in_do&_net_2);
   assign  _net_38 = (in_do&_net_2);
   assign  _net_39 = (in_do&_net_2);
   assign  _net_40 = (in_do&_net_2);
   assign  _net_41 = (in_do&_net_2);
   assign  _net_42 = (in_do&_net_2);
   assign  _net_43 = (in_do&_net_2);
   assign  _net_44 = (in_do&_net_2);
   assign  _net_45 = (in_do&_net_2);
   assign  _net_46 = (in_do&_net_2);
   assign  _net_47 = (in_do&_net_2);
   assign  _net_48 = (in_do&_net_2);
   assign  _net_49 = (in_do&_net_2);
   assign  _net_50 = (in_do&_net_2);
   assign  _net_51 = (in_do&_net_2);
   assign  _net_52 = (in_do&_net_2);
   assign  _net_53 = (in_do&_net_2);
   assign  _net_54 = (in_do&_net_2);
   assign  _net_55 = (in_do&_net_2);
   assign  _net_56 = (in_do&_net_2);
   assign  _net_57 = (in_do&_net_2);
   assign  _net_58 = (in_do&_net_2);
   assign  _net_59 = (in_do&_net_2);
   assign  _net_60 = (in_do&_net_2);
   assign  _net_61 = (in_do&_net_2);
   assign  _net_62 = (in_do&_net_2);
   assign  _net_63 = (in_do&_net_2);
   assign  _net_64 = (in_do&_net_2);
   assign  _net_65 = (in_do&_net_2);
   assign  _net_66 = (in_do&_net_2);
   assign  _net_67 = (in_do&_net_2);
   assign  _net_68 = (in_do&_net_2);
   assign  _net_69 = (in_do&_net_2);
   assign  _net_70 = (in_do&_net_2);
   assign  _net_71 = (in_do&_net_2);
   assign  _net_72 = (in_do&_net_2);
   assign  _net_73 = (in_do&_net_2);
   assign  _net_74 = (in_do&_net_2);
   assign  _net_75 = (in_do&_net_2);
   assign  _net_76 = (in_do&_net_2);
   assign  _net_77 = (in_do&_net_2);
   assign  _net_78 = (in_do&_net_2);
   assign  _net_79 = (in_do&_net_2);
   assign  _net_80 = (in_do&_net_2);
   assign  _net_81 = (in_do&_net_2);
   assign  _net_82 = (in_do&_net_2);
   assign  _net_83 = (in_do&_net_2);
   assign  _net_84 = (in_do&_net_2);
   assign  _net_85 = (in_do&_net_2);
   assign  _net_86 = (in_do&_net_2);
   assign  _net_87 = (in_do&_net_2);
   assign  _net_88 = (in_do&_net_2);
   assign  _net_89 = (in_do&_net_2);
   assign  _net_90 = (in_do&_net_2);
   assign  _net_91 = (in_do&_net_2);
   assign  _net_92 = (in_do&_net_2);
   assign  _net_93 = (in_do&_net_2);
   assign  _net_94 = (in_do&_net_2);
   assign  _net_95 = (in_do&_net_2);
   assign  _net_96 = (in_do&_net_2);
   assign  _net_97 = (in_do&_net_2);
   assign  _net_98 = (in_do&_net_2);
   assign  _net_99 = (in_do&_net_2);
   assign  _net_100 = (in_do&_net_2);
   assign  _net_101 = (in_do&_net_2);
   assign  _net_102 = (in_do&_net_2);
   assign  _net_103 = (in_do&_net_2);
   assign  _net_104 = (in_do&_net_2);
   assign  _net_105 = (in_do&_net_2);
   assign  _net_106 = (in_do&_net_2);
   assign  _net_107 = (in_do&_net_2);
   assign  _net_108 = (in_do&_net_2);
   assign  _net_109 = (in_do&_net_2);
   assign  _net_110 = (in_do&_net_2);
   assign  _net_111 = (in_do&_net_2);
   assign  _net_112 = (in_do&_net_2);
   assign  _net_113 = (in_do&_net_2);
   assign  _net_114 = (in_do&_net_2);
   assign  _net_115 = (in_do&_net_2);
   assign  _net_116 = (in_do&_net_2);
   assign  _net_117 = (in_do&_net_2);
   assign  _net_118 = (in_do&_net_2);
   assign  _net_119 = (in_do&_net_2);
   assign  _net_120 = (in_do&_net_2);
   assign  _net_121 = (in_do&_net_2);
   assign  _net_122 = (in_do&_net_2);
   assign  _net_123 = (in_do&_net_2);
   assign  _net_124 = (in_do&_net_2);
   assign  _net_125 = (in_do&_net_2);
   assign  _net_126 = (in_do&_net_2);
   assign  _net_127 = (in_do&_net_2);
   assign  _net_128 = (in_do&_net_2);
   assign  _net_129 = (in_do&_net_2);
   assign  _net_130 = (in_do&_net_2);
   assign  _net_131 = (in_do&_net_2);
   assign  _net_132 = (in_do&_net_2);
   assign  _net_133 = (in_do&_net_2);
   assign  _net_134 = (in_do&_net_2);
   assign  _net_135 = (in_do&_net_2);
   assign  _net_136 = (in_do&_net_2);
   assign  _net_137 = (in_do&_net_2);
   assign  _net_138 = (in_do&_net_2);
   assign  _net_139 = (in_do&_net_2);
   assign  _net_140 = (in_do&_net_2);
   assign  _net_141 = (in_do&_net_2);
   assign  _net_142 = (in_do&_net_2);
   assign  _net_143 = (in_do&_net_2);
   assign  _net_144 = (in_do&_net_2);
   assign  _net_145 = (in_do&_net_2);
   assign  _net_146 = (in_do&_net_2);
   assign  _net_147 = (in_do&_net_2);
   assign  _net_148 = (in_do&_net_2);
   assign  _net_149 = (in_do&_net_2);
   assign  _net_150 = (in_do&_net_2);
   assign  _net_151 = (in_do&_net_2);
   assign  _net_152 = (in_do&_net_2);
   assign  _net_153 = (in_do&_net_2);
   assign  _net_154 = (in_do&_net_2);
   assign  _net_155 = (in_do&_net_2);
   assign  _net_156 = (in_do&_net_2);
   assign  _net_157 = (in_do&_net_2);
   assign  _net_158 = (in_do&_net_2);
   assign  _net_159 = (in_do&_net_2);
   assign  _net_160 = (in_do&_net_2);
   assign  _net_161 = (in_do&_net_2);
   assign  _net_162 = (in_do&_net_2);
   assign  _net_163 = (in_do&_net_2);
   assign  _net_164 = (in_do&_net_2);
   assign  _net_165 = (in_do&_net_2);
   assign  _net_166 = (in_do&_net_2);
   assign  _net_167 = (in_do&_net_2);
   assign  _net_168 = (in_do&_net_2);
   assign  _net_169 = (in_do&_net_2);
   assign  _net_170 = (in_do&_net_2);
   assign  _net_171 = (in_do&_net_2);
   assign  _net_172 = (in_do&_net_2);
   assign  _net_173 = (in_do&_net_2);
   assign  _net_174 = (in_do&_net_2);
   assign  _net_175 = (in_do&_net_2);
   assign  _net_176 = (in_do&_net_2);
   assign  _net_177 = (in_do&_net_2);
   assign  _net_178 = (in_do&_net_2);
   assign  _net_179 = (in_do&_net_2);
   assign  _net_180 = (in_do&_net_2);
   assign  _net_181 = (in_do&_net_2);
   assign  _net_182 = (in_do&_net_2);
   assign  _net_183 = (in_do&_net_2);
   assign  _net_184 = (in_do&_net_2);
   assign  _net_185 = (in_do&_net_2);
   assign  _net_186 = (in_do&_net_2);
   assign  _net_187 = (in_do&_net_2);
   assign  _net_188 = (in_do&_net_2);
   assign  _net_189 = (in_do&_net_2);
   assign  _net_190 = (in_do&_net_2);
   assign  _net_191 = (in_do&_net_2);
   assign  _net_192 = (in_do&_net_2);
   assign  _net_193 = (in_do&_net_2);
   assign  _net_194 = (in_do&_net_2);
   assign  _net_195 = (in_do&_net_2);
   assign  _net_196 = (in_do&_net_2);
   assign  _net_197 = (in_do&_net_2);
   assign  _net_198 = (in_do&_net_2);
   assign  _net_199 = (in_do&_net_2);
   assign  _net_200 = (in_do&_net_2);
   assign  _net_201 = (in_do&_net_2);
   assign  _net_202 = (in_do&_net_2);
   assign  _net_203 = (in_do&_net_2);
   assign  _net_204 = (in_do&_net_2);
   assign  _net_205 = (in_do&_net_2);
   assign  _net_206 = (in_do&_net_2);
   assign  _net_207 = (in_do&_net_2);
   assign  _net_208 = (in_do&_net_2);
   assign  _net_209 = (in_do&_net_2);
   assign  _net_210 = (in_do&_net_2);
   assign  _net_211 = (in_do&_net_2);
   assign  _net_212 = (in_do&_net_2);
   assign  _net_213 = (in_do&_net_2);
   assign  _net_214 = (in_do&_net_2);
   assign  _net_215 = (in_do&_net_2);
   assign  _net_216 = (in_do&_net_2);
   assign  _net_217 = (in_do&_net_2);
   assign  _net_218 = (in_do&_net_2);
   assign  _net_219 = (in_do&_net_2);
   assign  _net_220 = (in_do&_net_2);
   assign  _net_221 = (in_do&_net_2);
   assign  _net_222 = (in_do&_net_2);
   assign  _net_223 = (in_do&_net_2);
   assign  _net_224 = (in_do&_net_2);
   assign  _net_225 = (in_do&_net_2);
   assign  _net_226 = (in_do&_net_2);
   assign  _net_227 = (in_do&_net_2);
   assign  _net_228 = (in_do&_net_2);
   assign  _net_229 = (in_do&_net_2);
   assign  _net_230 = (in_do&_net_2);
   assign  _net_231 = (in_do&_net_2);
   assign  _net_232 = (in_do&_net_2);
   assign  _net_233 = (in_do&_net_2);
   assign  _net_234 = (in_do&_net_2);
   assign  _net_235 = (in_do&_net_2);
   assign  _net_236 = (in_do&_net_2);
   assign  _net_237 = (in_do&_net_2);
   assign  _net_238 = (in_do&_net_2);
   assign  _net_239 = (in_do&_net_2);
   assign  _net_240 = (in_do&_net_2);
   assign  _net_241 = (in_do&_net_2);
   assign  _net_242 = (in_do&_net_2);
   assign  _net_243 = (in_do&_net_2);
   assign  _net_244 = (in_do&_net_2);
   assign  _net_245 = (in_do&_net_2);
   assign  _net_246 = (in_do&_net_2);
   assign  _net_247 = (in_do&_net_2);
   assign  _net_248 = (in_do&_net_2);
   assign  _net_249 = (in_do&_net_2);
   assign  _net_250 = (in_do&_net_2);
   assign  _net_251 = (in_do&_net_2);
   assign  _net_252 = (in_do&_net_2);
   assign  _net_253 = (in_do&_net_2);
   assign  _net_254 = (in_do&_net_2);
   assign  _net_255 = (in_do&_net_2);
   assign  _net_256 = (in_do&_net_2);
   assign  _net_257 = (in_do&_net_2);
   assign  _net_258 = (in_do&_net_2);
   assign  _net_259 = (in_do&_net_2);
   assign  _net_260 = (in_do&_net_2);
   assign  _net_261 = (in_do&_net_2);
   assign  _net_262 = (in_do&_net_2);
   assign  _net_263 = (in_do&_net_2);
   assign  _net_264 = (in_do&_net_2);
   assign  _net_265 = (in_do&_net_2);
   assign  _net_266 = (in_do&_net_2);
   assign  _net_267 = (in_do&_net_2);
   assign  _net_268 = (in_do&_net_2);
   assign  _net_269 = (in_do&_net_2);
   assign  _net_270 = (in_do&_net_2);
   assign  _net_271 = (in_do&_net_2);
   assign  _net_272 = (in_do&_net_2);
   assign  _net_273 = (in_do&_net_2);
   assign  _net_274 = (in_do&_net_2);
   assign  _net_275 = (in_do&_net_2);
   assign  _net_276 = (in_do&_net_2);
   assign  _net_277 = (in_do&_net_2);
   assign  _net_278 = (in_do&_net_2);
   assign  _net_279 = (in_do&_net_2);
   assign  _net_280 = (in_do&_net_2);
   assign  _net_281 = (in_do&_net_2);
   assign  _net_282 = (in_do&_net_2);
   assign  _net_283 = (in_do&_net_2);
   assign  _net_284 = (in_do&_net_2);
   assign  _net_285 = (in_do&_net_2);
   assign  _net_286 = (in_do&_net_2);
   assign  _net_287 = (in_do&_net_2);
   assign  _net_288 = (in_do&_net_2);
   assign  _net_289 = (in_do&_net_2);
   assign  _net_290 = (in_do&_net_2);
   assign  _net_291 = (in_do&_net_2);
   assign  _net_292 = (in_do&_net_2);
   assign  _net_293 = (in_do&_net_2);
   assign  _net_294 = (in_do&_net_2);
   assign  _net_295 = (in_do&_net_2);
   assign  _net_296 = (in_do&_net_2);
   assign  _net_297 = (in_do&_net_2);
   assign  _net_298 = (in_do&_net_2);
   assign  _net_299 = (in_do&_net_2);
   assign  _net_300 = (in_do&_net_2);
   assign  _net_301 = (in_do&_net_2);
   assign  _net_302 = (in_do&_net_2);
   assign  _net_303 = (in_do&_net_2);
   assign  _net_304 = (in_do&_net_2);
   assign  _net_305 = (in_do&_net_2);
   assign  _net_306 = (in_do&_net_2);
   assign  _net_307 = (in_do&_net_2);
   assign  _net_308 = (in_do&_net_2);
   assign  _net_309 = (in_do&_net_2);
   assign  _net_310 = (in_do&_net_2);
   assign  _net_311 = (in_do&_net_2);
   assign  _net_312 = (in_do&_net_2);
   assign  _net_313 = (in_do&_net_2);
   assign  _net_314 = (in_do&_net_2);
   assign  _net_315 = (in_do&_net_2);
   assign  _net_316 = (in_do&_net_2);
   assign  _net_317 = (in_do&_net_2);
   assign  _net_318 = (in_do&_net_2);
   assign  _net_319 = (in_do&_net_2);
   assign  _net_320 = (in_do&_net_2);
   assign  _net_321 = (in_do&_net_2);
   assign  _net_322 = (in_do&_net_2);
   assign  _net_323 = (in_do&_net_2);
   assign  _net_324 = (in_do&_net_2);
   assign  _net_325 = (in_do&_net_2);
   assign  _net_326 = (in_do&_net_2);
   assign  _net_327 = (in_do&_net_2);
   assign  _net_328 = (in_do&_net_2);
   assign  _net_329 = (in_do&_net_2);
   assign  _net_330 = (in_do&_net_2);
   assign  _net_331 = (in_do&_net_2);
   assign  _net_332 = (in_do&_net_2);
   assign  _net_333 = (in_do&_net_2);
   assign  _net_334 = (in_do&_net_2);
   assign  _net_335 = (in_do&_net_2);
   assign  _net_336 = (in_do&_net_2);
   assign  _net_337 = (in_do&_net_2);
   assign  _net_338 = (in_do&_net_2);
   assign  _net_339 = (in_do&_net_2);
   assign  _net_340 = (in_do&_net_2);
   assign  _net_341 = (in_do&_net_2);
   assign  _net_342 = (in_do&_net_2);
   assign  _net_343 = (in_do&_net_2);
   assign  _net_344 = (in_do&_net_2);
   assign  _net_345 = (in_do&_net_2);
   assign  _net_346 = (in_do&_net_2);
   assign  _net_347 = (in_do&_net_2);
   assign  _net_348 = (in_do&_net_2);
   assign  _net_349 = (in_do&_net_2);
   assign  _net_350 = (in_do&_net_2);
   assign  _net_351 = (in_do&_net_2);
   assign  _net_352 = (in_do&_net_2);
   assign  _net_353 = (in_do&_net_2);
   assign  _net_354 = (in_do&_net_2);
   assign  _net_355 = (in_do&_net_2);
   assign  _net_356 = (in_do&_net_2);
   assign  _net_357 = (in_do&_net_2);
   assign  _net_358 = (in_do&_net_2);
   assign  _net_359 = (in_do&_net_2);
   assign  _net_360 = (in_do&_net_2);
   assign  _net_361 = (in_do&_net_2);
   assign  _net_362 = (in_do&_net_2);
   assign  _net_363 = (in_do&_net_2);
   assign  _net_364 = (in_do&_net_2);
   assign  _net_365 = (in_do&_net_2);
   assign  _net_366 = (in_do&_net_2);
   assign  _net_367 = (in_do&_net_2);
   assign  _net_368 = (in_do&_net_2);
   assign  _net_369 = (in_do&_net_2);
   assign  _net_370 = (in_do&_net_2);
   assign  _net_371 = (in_do&_net_2);
   assign  _net_372 = (in_do&_net_2);
   assign  _net_373 = (in_do&_net_2);
   assign  _net_374 = (in_do&_net_2);
   assign  _net_375 = (in_do&_net_2);
   assign  _net_376 = (in_do&_net_2);
   assign  _net_377 = (in_do&_net_2);
   assign  _net_378 = (in_do&_net_2);
   assign  _net_379 = (in_do&_net_2);
   assign  _net_380 = (in_do&_net_2);
   assign  _net_381 = (in_do&_net_2);
   assign  _net_382 = (in_do&_net_2);
   assign  _net_383 = (in_do&_net_2);
   assign  _net_384 = (in_do&_net_2);
   assign  _net_385 = (in_do&_net_2);
   assign  _net_386 = (in_do&_net_2);
   assign  _net_387 = (in_do&_net_2);
   assign  _net_388 = (in_do&_net_2);
   assign  _net_389 = (in_do&_net_2);
   assign  _net_390 = (in_do&_net_2);
   assign  _net_391 = (in_do&_net_2);
   assign  _net_392 = (in_do&_net_2);
   assign  _net_393 = (in_do&_net_2);
   assign  _net_394 = (in_do&_net_2);
   assign  _net_395 = (in_do&_net_2);
   assign  _net_396 = (in_do&_net_2);
   assign  _net_397 = (in_do&_net_2);
   assign  _net_398 = (in_do&_net_2);
   assign  _net_399 = (in_do&_net_2);
   assign  _net_400 = (in_do&_net_2);
   assign  _net_401 = (in_do&_net_2);
   assign  _net_402 = (in_do&_net_2);
   assign  _net_403 = (in_do&_net_2);
   assign  _net_404 = (in_do&_net_2);
   assign  _net_405 = (in_do&_net_2);
   assign  _net_406 = (in_do&_net_2);
   assign  _net_407 = (in_do&_net_2);
   assign  _net_408 = (in_do&_net_2);
   assign  _net_409 = (in_do&_net_2);
   assign  _net_410 = (in_do&_net_2);
   assign  _net_411 = (in_do&_net_2);
   assign  _net_412 = (in_do&_net_2);
   assign  _net_413 = (in_do&_net_2);
   assign  _net_414 = (in_do&_net_2);
   assign  _net_415 = (in_do&_net_2);
   assign  _net_416 = (in_do&_net_2);
   assign  _net_417 = (in_do&_net_2);
   assign  _net_418 = (in_do&_net_2);
   assign  _net_419 = (in_do&_net_2);
   assign  _net_420 = (in_do&_net_2);
   assign  _net_421 = (in_do&_net_2);
   assign  _net_422 = (in_do&_net_2);
   assign  _net_423 = (in_do&_net_2);
   assign  _net_424 = (in_do&_net_2);
   assign  _net_425 = (in_do&_net_2);
   assign  _net_426 = (in_do&_net_2);
   assign  _net_427 = (in_do&_net_2);
   assign  _net_428 = (in_do&_net_2);
   assign  _net_429 = (in_do&_net_2);
   assign  _net_430 = (in_do&_net_2);
   assign  _net_431 = (in_do&_net_2);
   assign  _net_432 = (in_do&_net_2);
   assign  _net_433 = (in_do&_net_2);
   assign  _net_434 = (in_do&_net_2);
   assign  _net_435 = (in_do&_net_2);
   assign  _net_436 = (in_do&_net_2);
   assign  _net_437 = (in_do&_net_2);
   assign  _net_438 = (in_do&_net_2);
   assign  _net_439 = (in_do&_net_2);
   assign  _net_440 = (in_do&_net_2);
   assign  _net_441 = (in_do&_net_2);
   assign  _net_442 = (in_do&_net_2);
   assign  _net_443 = (in_do&_net_2);
   assign  _net_444 = (in_do&_net_2);
   assign  _net_445 = (in_do&_net_2);
   assign  _net_446 = (in_do&_net_2);
   assign  _net_447 = (in_do&_net_2);
   assign  _net_448 = (in_do&_net_2);
   assign  _net_449 = (in_do&_net_2);
   assign  _net_450 = (in_do&_net_2);
   assign  _net_451 = (in_do&_net_2);
   assign  _net_452 = (in_do&_net_2);
   assign  _net_453 = (in_do&_net_2);
   assign  _net_454 = (in_do&_net_2);
   assign  _net_455 = (in_do&_net_2);
   assign  _net_456 = (in_do&_net_2);
   assign  _net_457 = (in_do&_net_2);
   assign  _net_458 = (in_do&_net_2);
   assign  _net_459 = (in_do&_net_2);
   assign  _net_460 = (in_do&_net_2);
   assign  _net_461 = (in_do&_net_2);
   assign  _net_462 = (in_do&_net_2);
   assign  _net_463 = (in_do&_net_2);
   assign  _net_464 = (in_do&_net_2);
   assign  _net_465 = (in_do&_net_2);
   assign  _net_466 = (in_do&_net_2);
   assign  _net_467 = (in_do&_net_2);
   assign  _net_468 = (in_do&_net_2);
   assign  _net_469 = (in_do&_net_2);
   assign  _net_470 = (in_do&_net_2);
   assign  _net_471 = (in_do&_net_2);
   assign  _net_472 = (in_do&_net_2);
   assign  _net_473 = (in_do&_net_2);
   assign  _net_474 = (in_do&_net_2);
   assign  _net_475 = (in_do&_net_2);
   assign  _net_476 = (in_do&_net_2);
   assign  _net_477 = (in_do&_net_2);
   assign  _net_478 = (in_do&_net_2);
   assign  _net_479 = (in_do&_net_2);
   assign  _net_480 = (in_do&_net_2);
   assign  _net_481 = (in_do&_net_2);
   assign  _net_482 = (in_do&_net_2);
   assign  _net_483 = (in_do&_net_2);
   assign  _net_484 = (in_do&_net_2);
   assign  _net_485 = (in_do&_net_2);
   assign  _net_486 = (in_do&_net_2);
   assign  _net_487 = (in_do&_net_2);
   assign  _net_488 = (in_do&_net_2);
   assign  _net_489 = (in_do&_net_2);
   assign  _net_490 = (in_do&_net_2);
   assign  _net_491 = (in_do&_net_2);
   assign  _net_492 = (in_do&_net_2);
   assign  _net_493 = (in_do&_net_2);
   assign  _net_494 = (in_do&_net_2);
   assign  _net_495 = (in_do&_net_2);
   assign  _net_496 = (in_do&_net_2);
   assign  _net_497 = (in_do&_net_2);
   assign  _net_498 = (in_do&_net_2);
   assign  _net_499 = (in_do&_net_2);
   assign  _net_500 = (in_do&_net_2);
   assign  _net_501 = (in_do&_net_2);
   assign  _net_502 = (in_do&_net_2);
   assign  _net_503 = (in_do&_net_2);
   assign  _net_504 = (in_do&_net_2);
   assign  _net_505 = (in_do&_net_2);
   assign  _net_506 = (in_do&_net_2);
   assign  _net_507 = (in_do&_net_2);
   assign  _net_508 = (in_do&_net_2);
   assign  _net_509 = (in_do&_net_2);
   assign  _net_510 = (in_do&_net_2);
   assign  _net_511 = (in_do&_net_2);
   assign  _net_512 = (in_do&_net_2);
   assign  _net_513 = (in_do&_net_2);
   assign  _net_514 = (in_do&_net_2);
   assign  _net_515 = (in_do&_net_2);
   assign  _net_516 = (in_do&_net_2);
   assign  _net_517 = (in_do&_net_2);
   assign  _net_518 = (in_do&_net_2);
   assign  _net_519 = (in_do&_net_2);
   assign  _net_520 = (in_do&_net_2);
   assign  _net_521 = (in_do&_net_2);
   assign  _net_522 = (in_do&_net_2);
   assign  _net_523 = (in_do&_net_2);
   assign  _net_524 = (in_do&_net_2);
   assign  _net_525 = (in_do&_net_2);
   assign  _net_526 = (in_do&_net_2);
   assign  _net_527 = (in_do&_net_2);
   assign  _net_528 = (in_do&_net_2);
   assign  _net_529 = (in_do&_net_2);
   assign  _net_530 = (in_do&_net_2);
   assign  _net_531 = (in_do&_net_2);
   assign  _net_532 = (in_do&_net_2);
   assign  _net_533 = (in_do&_net_2);
   assign  _net_534 = (in_do&_net_2);
   assign  _net_535 = (in_do&_net_2);
   assign  _net_536 = (in_do&_net_2);
   assign  _net_537 = (in_do&_net_2);
   assign  _net_538 = (in_do&_net_2);
   assign  _net_539 = (in_do&_net_2);
   assign  _net_540 = (in_do&_net_2);
   assign  _net_541 = (in_do&_net_2);
   assign  _net_542 = (in_do&_net_2);
   assign  _net_543 = (in_do&_net_2);
   assign  _net_544 = (in_do&_net_2);
   assign  _net_545 = (in_do&_net_2);
   assign  _net_546 = (in_do&_net_2);
   assign  _net_547 = (in_do&_net_2);
   assign  _net_548 = (in_do&_net_2);
   assign  _net_549 = (in_do&_net_2);
   assign  _net_550 = (in_do&_net_2);
   assign  _net_551 = (in_do&_net_2);
   assign  _net_552 = (in_do&_net_2);
   assign  _net_553 = (in_do&_net_2);
   assign  _net_554 = (in_do&_net_2);
   assign  _net_555 = (in_do&_net_2);
   assign  _net_556 = (in_do&_net_2);
   assign  _net_557 = (in_do&_net_2);
   assign  _net_558 = (in_do&_net_2);
   assign  _net_559 = (in_do&_net_2);
   assign  _net_560 = (in_do&_net_2);
   assign  _net_561 = (in_do&_net_2);
   assign  _net_562 = (in_do&_net_2);
   assign  _net_563 = (in_do&_net_2);
   assign  _net_564 = (in_do&_net_2);
   assign  _net_565 = (in_do&_net_2);
   assign  _net_566 = (in_do&_net_2);
   assign  _net_567 = (in_do&_net_2);
   assign  _net_568 = (in_do&_net_2);
   assign  _net_569 = (in_do&_net_2);
   assign  _net_570 = (in_do&_net_2);
   assign  _net_571 = (in_do&_net_2);
   assign  _net_572 = (in_do&_net_2);
   assign  _net_573 = (in_do&_net_2);
   assign  _net_574 = (in_do&_net_2);
   assign  _net_575 = (in_do&_net_2);
   assign  _net_576 = (in_do&_net_2);
   assign  _net_577 = (in_do&_net_2);
   assign  _net_578 = (in_do&_net_2);
   assign  _net_579 = (in_do&_net_2);
   assign  _net_580 = (in_do&_net_2);
   assign  _net_581 = (in_do&_net_2);
   assign  _net_582 = (in_do&_net_2);
   assign  _net_583 = (in_do&_net_2);
   assign  _net_584 = (in_do&_net_2);
   assign  _net_585 = (in_do&_net_2);
   assign  _net_586 = (in_do&_net_2);
   assign  _net_587 = (in_do&_net_2);
   assign  _net_588 = (in_do&_net_2);
   assign  _net_589 = (in_do&_net_2);
   assign  _net_590 = (in_do&_net_2);
   assign  _net_591 = (in_do&_net_2);
   assign  _net_592 = (in_do&_net_2);
   assign  _net_593 = (in_do&_net_2);
   assign  _net_594 = (in_do&_net_2);
   assign  _net_595 = (in_do&_net_2);
   assign  _net_596 = (in_do&_net_2);
   assign  _net_597 = (in_do&_net_2);
   assign  _net_598 = (in_do&_net_2);
   assign  _net_599 = (in_do&_net_2);
   assign  _net_600 = (in_do&_net_2);
   assign  _net_601 = (in_do&_net_2);
   assign  _net_602 = (in_do&_net_2);
   assign  _net_603 = (in_do&_net_2);
   assign  _net_604 = (in_do&_net_2);
   assign  _net_605 = (in_do&_net_2);
   assign  _net_606 = (in_do&_net_2);
   assign  _net_607 = (in_do&_net_2);
   assign  _net_608 = (in_do&_net_2);
   assign  _net_609 = (in_do&_net_2);
   assign  _net_610 = (in_do&_net_2);
   assign  _net_611 = (in_do&_net_2);
   assign  _net_612 = (in_do&_net_2);
   assign  _net_613 = (in_do&_net_2);
   assign  _net_614 = (in_do&_net_2);
   assign  _net_615 = (in_do&_net_2);
   assign  _net_616 = (in_do&_net_2);
   assign  _net_617 = (in_do&_net_2);
   assign  _net_618 = (in_do&_net_2);
   assign  _net_619 = (in_do&_net_2);
   assign  _net_620 = (in_do&_net_2);
   assign  _net_621 = (in_do&_net_2);
   assign  _net_622 = (in_do&_net_2);
   assign  _net_623 = (in_do&_net_2);
   assign  _net_624 = (in_do&_net_2);
   assign  _net_625 = (in_do&_net_2);
   assign  _net_626 = (in_do&_net_2);
   assign  _net_627 = (in_do&_net_2);
   assign  _net_628 = (in_do&_net_2);
   assign  _net_629 = (in_do&_net_2);
   assign  _net_630 = (in_do&_net_2);
   assign  _net_631 = (in_do&_net_2);
   assign  _net_632 = (in_do&_net_2);
   assign  _net_633 = (in_do&_net_2);
   assign  _net_634 = (in_do&_net_2);
   assign  _net_635 = (in_do&_net_2);
   assign  _net_636 = (in_do&_net_2);
   assign  _net_637 = (in_do&_net_2);
   assign  _net_638 = (in_do&_net_2);
   assign  _net_639 = (in_do&_net_2);
   assign  _net_640 = (in_do&_net_2);
   assign  _net_641 = (in_do&_net_2);
   assign  _net_642 = (in_do&_net_2);
   assign  _net_643 = (in_do&_net_2);
   assign  _net_644 = (in_do&_net_2);
   assign  _net_645 = (in_do&_net_2);
   assign  _net_646 = (in_do&_net_2);
   assign  _net_647 = (in_do&_net_2);
   assign  _net_648 = (in_do&_net_2);
   assign  _net_649 = (in_do&_net_2);
   assign  _net_650 = (in_do&_net_2);
   assign  _net_651 = (in_do&_net_2);
   assign  _net_652 = (in_do&_net_2);
   assign  _net_653 = (in_do&_net_2);
   assign  _net_654 = (in_do&_net_2);
   assign  _net_655 = (in_do&_net_2);
   assign  _net_656 = (in_do&_net_2);
   assign  _net_657 = (in_do&_net_2);
   assign  _net_658 = (in_do&_net_2);
   assign  _net_659 = (in_do&_net_2);
   assign  _net_660 = (in_do&_net_2);
   assign  _net_661 = (in_do&_net_2);
   assign  _net_662 = (in_do&_net_2);
   assign  _net_663 = (in_do&_net_2);
   assign  _net_664 = (in_do&_net_2);
   assign  _net_665 = (in_do&_net_2);
   assign  _net_666 = (in_do&_net_2);
   assign  _net_667 = (in_do&_net_2);
   assign  _net_668 = (in_do&_net_2);
   assign  _net_669 = (in_do&_net_2);
   assign  _net_670 = (in_do&_net_2);
   assign  _net_671 = (in_do&_net_2);
   assign  _net_672 = (in_do&_net_2);
   assign  _net_673 = (in_do&_net_2);
   assign  _net_674 = (in_do&_net_2);
   assign  _net_675 = (in_do&_net_2);
   assign  _net_676 = (in_do&_net_2);
   assign  _net_677 = (in_do&_net_2);
   assign  _net_678 = (in_do&_net_2);
   assign  _net_679 = (in_do&_net_2);
   assign  _net_680 = (in_do&_net_2);
   assign  _net_681 = (in_do&_net_2);
   assign  _net_682 = (in_do&_net_2);
   assign  _net_683 = (in_do&_net_2);
   assign  _net_684 = (in_do&_net_2);
   assign  _net_685 = (in_do&_net_2);
   assign  _net_686 = (in_do&_net_2);
   assign  _net_687 = (in_do&_net_2);
   assign  _net_688 = (in_do&_net_2);
   assign  _net_689 = (in_do&_net_2);
   assign  _net_690 = (in_do&_net_2);
   assign  _net_691 = (in_do&_net_2);
   assign  _net_692 = (in_do&_net_2);
   assign  _net_693 = (in_do&_net_2);
   assign  _net_694 = (in_do&_net_2);
   assign  _net_695 = (in_do&_net_2);
   assign  _net_696 = (in_do&_net_2);
   assign  _net_697 = (in_do&_net_2);
   assign  _net_698 = (in_do&_net_2);
   assign  _net_699 = (in_do&_net_2);
   assign  _net_700 = (in_do&_net_2);
   assign  _net_701 = (in_do&_net_2);
   assign  _net_702 = (in_do&_net_2);
   assign  _net_703 = (in_do&_net_2);
   assign  _net_704 = (in_do&_net_2);
   assign  _net_705 = (in_do&_net_2);
   assign  _net_706 = (in_do&_net_2);
   assign  _net_707 = (in_do&_net_2);
   assign  _net_708 = (in_do&_net_2);
   assign  _net_709 = (in_do&_net_2);
   assign  _net_710 = (in_do&_net_2);
   assign  _net_711 = (in_do&_net_2);
   assign  _net_712 = (in_do&_net_2);
   assign  _net_713 = (in_do&_net_2);
   assign  _net_714 = (in_do&_net_2);
   assign  _net_715 = (in_do&_net_2);
   assign  _net_716 = (in_do&_net_2);
   assign  _net_717 = (in_do&_net_2);
   assign  _net_718 = (in_do&_net_2);
   assign  _net_719 = (in_do&_net_2);
   assign  _net_720 = (in_do&_net_2);
   assign  _net_721 = (in_do&_net_2);
   assign  _net_722 = (in_do&_net_2);
   assign  _net_723 = (in_do&_net_2);
   assign  _net_724 = (in_do&_net_2);
   assign  _net_725 = (in_do&_net_2);
   assign  _net_726 = (in_do&_net_2);
   assign  _net_727 = (in_do&_net_2);
   assign  _net_728 = (in_do&_net_2);
   assign  _net_729 = (in_do&_net_2);
   assign  _net_730 = (in_do&_net_2);
   assign  _net_731 = (in_do&_net_2);
   assign  _net_732 = (in_do&_net_2);
   assign  _net_733 = (in_do&_net_2);
   assign  _net_734 = (in_do&_net_2);
   assign  _net_735 = (in_do&_net_2);
   assign  _net_736 = (in_do&_net_2);
   assign  _net_737 = (in_do&_net_2);
   assign  _net_738 = (in_do&_net_2);
   assign  _net_739 = (in_do&_net_2);
   assign  _net_740 = (in_do&_net_2);
   assign  _net_741 = (in_do&_net_2);
   assign  _net_742 = (in_do&_net_2);
   assign  _net_743 = (in_do&_net_2);
   assign  _net_744 = (in_do&_net_2);
   assign  _net_745 = (in_do&_net_2);
   assign  _net_746 = (in_do&_net_2);
   assign  _net_747 = (in_do&_net_2);
   assign  _net_748 = (in_do&_net_2);
   assign  _net_749 = (in_do&_net_2);
   assign  _net_750 = (in_do&_net_2);
   assign  _net_751 = (in_do&_net_2);
   assign  _net_752 = (in_do&_net_2);
   assign  _net_753 = (in_do&_net_2);
   assign  _net_754 = (in_do&_net_2);
   assign  _net_755 = (in_do&_net_2);
   assign  _net_756 = (in_do&_net_2);
   assign  _net_757 = (in_do&_net_2);
   assign  _net_758 = (in_do&_net_2);
   assign  _net_759 = (in_do&_net_2);
   assign  _net_760 = (in_do&_net_2);
   assign  _net_761 = (in_do&_net_2);
   assign  _net_762 = (in_do&_net_2);
   assign  _net_763 = (in_do&_net_2);
   assign  _net_764 = (in_do&_net_2);
   assign  _net_765 = (in_do&_net_2);
   assign  _net_766 = (in_do&_net_2);
   assign  _net_767 = (in_do&_net_2);
   assign  _net_768 = (in_do&_net_2);
   assign  _net_769 = (in_do&_net_2);
   assign  _net_770 = (in_do&_net_2);
   assign  _net_771 = (in_do&_net_2);
   assign  _net_772 = (in_do&_net_2);
   assign  _net_773 = (in_do&_net_2);
   assign  _net_774 = (in_do&_net_2);
   assign  _net_775 = (in_do&_net_2);
   assign  _net_776 = (in_do&_net_2);
   assign  _net_777 = (in_do&_net_2);
   assign  _net_778 = (in_do&_net_2);
   assign  _net_779 = (in_do&_net_2);
   assign  _net_780 = (in_do&_net_2);
   assign  _net_781 = (in_do&_net_2);
   assign  _net_782 = (in_do&_net_2);
   assign  _net_783 = (in_do&_net_2);
   assign  _net_784 = (in_do&_net_2);
   assign  _net_785 = (in_do&_net_2);
   assign  _net_786 = (in_do&_net_2);
   assign  _net_787 = (in_do&_net_2);
   assign  _net_788 = (in_do&_net_2);
   assign  _net_789 = (in_do&_net_2);
   assign  _net_790 = (in_do&_net_2);
   assign  _net_791 = (in_do&_net_2);
   assign  _net_792 = (in_do&_net_2);
   assign  _net_793 = (in_do&_net_2);
   assign  _net_794 = (in_do&_net_2);
   assign  _net_795 = (in_do&_net_2);
   assign  _net_796 = (in_do&_net_2);
   assign  _net_797 = (in_do&_net_2);
   assign  _net_798 = (in_do&_net_2);
   assign  _net_799 = (in_do&_net_2);
   assign  _net_800 = (in_do&_net_2);
   assign  _net_801 = (in_do&_net_2);
   assign  _net_802 = (in_do&_net_2);
   assign  _net_803 = (in_do&_net_2);
   assign  _net_804 = (in_do&_net_2);
   assign  _net_805 = (in_do&_net_2);
   assign  _net_806 = (in_do&_net_2);
   assign  _net_807 = (in_do&_net_2);
   assign  _net_808 = (in_do&_net_2);
   assign  _net_809 = (in_do&_net_2);
   assign  _net_810 = (in_do&_net_2);
   assign  _net_811 = (in_do&_net_2);
   assign  _net_812 = (in_do&_net_2);
   assign  _net_813 = (in_do&_net_2);
   assign  _net_814 = (in_do&_net_2);
   assign  _net_815 = (in_do&_net_2);
   assign  _net_816 = (in_do&_net_2);
   assign  _net_817 = (in_do&_net_2);
   assign  _net_818 = (in_do&_net_2);
   assign  _net_819 = (in_do&_net_2);
   assign  _net_820 = (in_do&_net_2);
   assign  _net_821 = (in_do&_net_2);
   assign  _net_822 = (in_do&_net_2);
   assign  _net_823 = (in_do&_net_2);
   assign  _net_824 = (in_do&_net_2);
   assign  _net_825 = (in_do&_net_2);
   assign  _net_826 = (in_do&_net_2);
   assign  _net_827 = (in_do&_net_2);
   assign  _net_828 = (in_do&_net_2);
   assign  _net_829 = (in_do&_net_2);
   assign  _net_830 = (in_do&_net_2);
   assign  _net_831 = (in_do&_net_2);
   assign  _net_832 = (in_do&_net_2);
   assign  _net_833 = (in_do&_net_2);
   assign  _net_834 = (in_do&_net_2);
   assign  _net_835 = (in_do&_net_2);
   assign  _net_836 = (in_do&_net_2);
   assign  _net_837 = (in_do&_net_2);
   assign  _net_838 = (in_do&_net_2);
   assign  _net_839 = (in_do&_net_2);
   assign  _net_840 = (in_do&_net_2);
   assign  _net_841 = (in_do&_net_2);
   assign  _net_842 = (in_do&_net_2);
   assign  _net_843 = (in_do&_net_2);
   assign  _net_844 = (in_do&_net_2);
   assign  _net_845 = (in_do&_net_2);
   assign  _net_846 = (in_do&_net_2);
   assign  _net_847 = (in_do&_net_2);
   assign  _net_848 = (in_do&_net_2);
   assign  _net_849 = (in_do&_net_2);
   assign  _net_850 = (in_do&_net_2);
   assign  _net_851 = (in_do&_net_2);
   assign  _net_852 = (in_do&_net_2);
   assign  _net_853 = (in_do&_net_2);
   assign  _net_854 = (in_do&_net_2);
   assign  _net_855 = (in_do&_net_2);
   assign  _net_856 = (in_do&_net_2);
   assign  _net_857 = (in_do&_net_2);
   assign  _net_858 = (in_do&_net_2);
   assign  _net_859 = (in_do&_net_2);
   assign  _net_860 = (in_do&_net_2);
   assign  _net_861 = (in_do&_net_2);
   assign  _net_862 = (in_do&_net_2);
   assign  _net_863 = (in_do&_net_2);
   assign  _net_864 = (in_do&_net_2);
   assign  _net_865 = (in_do&_net_2);
   assign  _net_866 = (in_do&_net_2);
   assign  _net_867 = (in_do&_net_2);
   assign  _net_868 = (in_do&_net_2);
   assign  _net_869 = (in_do&_net_2);
   assign  _net_870 = (in_do&_net_2);
   assign  _net_871 = (in_do&_net_2);
   assign  _net_872 = (in_do&_net_2);
   assign  _net_873 = (in_do&_net_2);
   assign  _net_874 = (in_do&_net_2);
   assign  _net_875 = (in_do&_net_2);
   assign  _net_876 = (in_do&_net_2);
   assign  _net_877 = (in_do&_net_2);
   assign  _net_878 = (in_do&_net_2);
   assign  _net_879 = (in_do&_net_2);
   assign  _net_880 = (in_do&_net_2);
   assign  _net_881 = (in_do&_net_2);
   assign  _net_882 = (in_do&_net_2);
   assign  _net_883 = (in_do&_net_2);
   assign  _net_884 = (in_do&_net_2);
   assign  _net_885 = (in_do&_net_2);
   assign  _net_886 = (in_do&_net_2);
   assign  _net_887 = (in_do&_net_2);
   assign  _net_888 = (in_do&_net_2);
   assign  _net_889 = (in_do&_net_2);
   assign  _net_890 = (in_do&_net_2);
   assign  _net_891 = (in_do&_net_2);
   assign  _net_892 = (in_do&_net_2);
   assign  _net_893 = (in_do&_net_2);
   assign  _net_894 = (in_do&_net_2);
   assign  _net_895 = (in_do&_net_2);
   assign  _net_896 = (in_do&_net_2);
   assign  _net_897 = (in_do&_net_2);
   assign  _net_898 = (in_do&_net_2);
   assign  _net_899 = (in_do&_net_2);
   assign  _net_900 = (in_do&_net_2);
   assign  _net_901 = (in_do&_net_2);
   assign  _net_902 = (in_do&_net_2);
   assign  _net_903 = (in_do&_net_2);
   assign  _net_904 = (in_do&_net_2);
   assign  _net_905 = (in_do&_net_2);
   assign  _net_906 = (in_do&_net_2);
   assign  _net_907 = (in_do&_net_2);
   assign  _net_908 = (in_do&_net_2);
   assign  _net_909 = (in_do&_net_2);
   assign  _net_910 = (in_do&_net_2);
   assign  _net_911 = (in_do&_net_2);
   assign  _net_912 = (in_do&_net_2);
   assign  _net_913 = (in_do&_net_2);
   assign  _net_914 = (in_do&_net_2);
   assign  _net_915 = (in_do&_net_2);
   assign  _net_916 = (in_do&_net_2);
   assign  _net_917 = (in_do&_net_2);
   assign  _net_918 = (in_do&_net_2);
   assign  _net_919 = (in_do&_net_2);
   assign  _net_920 = (in_do&_net_2);
   assign  _net_921 = (in_do&_net_2);
   assign  _net_922 = (in_do&_net_2);
   assign  _net_923 = (in_do&_net_2);
   assign  _net_924 = (in_do&_net_2);
   assign  _net_925 = (in_do&_net_2);
   assign  _net_926 = (in_do&_net_2);
   assign  _net_927 = (in_do&_net_2);
   assign  _net_928 = (in_do&_net_2);
   assign  _net_929 = (in_do&_net_2);
   assign  _net_930 = (in_do&_net_2);
   assign  _net_931 = (in_do&_net_2);
   assign  _net_932 = (in_do&_net_2);
   assign  _net_933 = (in_do&_net_2);
   assign  _net_934 = (in_do&_net_2);
   assign  _net_935 = (in_do&_net_2);
   assign  _net_936 = (in_do&_net_2);
   assign  _net_937 = (in_do&_net_2);
   assign  _net_938 = (in_do&_net_2);
   assign  _net_939 = (in_do&_net_2);
   assign  _net_940 = (in_do&_net_2);
   assign  _net_941 = (in_do&_net_2);
   assign  _net_942 = (in_do&_net_2);
   assign  _net_943 = (in_do&_net_2);
   assign  _net_944 = (in_do&_net_2);
   assign  _net_945 = (in_do&_net_2);
   assign  _net_946 = (in_do&_net_2);
   assign  _net_947 = (in_do&_net_2);
   assign  _net_948 = (in_do&_net_2);
   assign  _net_949 = (in_do&_net_2);
   assign  _net_950 = (in_do&_net_2);
   assign  _net_951 = (in_do&_net_2);
   assign  _net_952 = (in_do&_net_2);
   assign  _net_953 = (in_do&_net_2);
   assign  _net_954 = (in_do&_net_2);
   assign  _net_955 = (in_do&_net_2);
   assign  _net_956 = (in_do&_net_2);
   assign  _net_957 = (in_do&_net_2);
   assign  _net_958 = (in_do&_net_2);
   assign  _net_959 = (in_do&_net_2);
   assign  _net_960 = (in_do&_net_2);
   assign  _net_961 = (in_do&_net_2);
   assign  _net_962 = (in_do&_net_2);
   assign  _net_963 = (in_do&_net_2);
   assign  _net_964 = (in_do&_net_2);
   assign  _net_965 = (in_do&_net_2);
   assign  _net_966 = (in_do&_net_2);
   assign  _net_967 = (in_do&_net_2);
   assign  _net_968 = (in_do&_net_2);
   assign  _net_969 = (in_do&_net_2);
   assign  _net_970 = (in_do&_net_2);
   assign  _net_971 = (in_do&_net_2);
   assign  _net_972 = (in_do&_net_2);
   assign  _net_973 = (in_do&_net_2);
   assign  _net_974 = (in_do&_net_2);
   assign  _net_975 = (in_do&_net_2);
   assign  _net_976 = (in_do&_net_2);
   assign  _net_977 = (in_do&_net_2);
   assign  _net_978 = (in_do&_net_2);
   assign  _net_979 = (in_do&_net_2);
   assign  _net_980 = (in_do&_net_2);
   assign  _net_981 = (in_do&_net_2);
   assign  _net_982 = (in_do&_net_2);
   assign  _net_983 = (in_do&_net_2);
   assign  _net_984 = (in_do&_net_2);
   assign  _net_985 = (in_do&_net_2);
   assign  _net_986 = (in_do&_net_2);
   assign  _net_987 = (in_do&_net_2);
   assign  _net_988 = (in_do&_net_2);
   assign  _net_989 = (in_do&_net_2);
   assign  _net_990 = (in_do&_net_2);
   assign  _net_991 = (in_do&_net_2);
   assign  _net_992 = (in_do&_net_2);
   assign  _net_993 = (in_do&_net_2);
   assign  _net_994 = (in_do&_net_2);
   assign  _net_995 = (in_do&_net_2);
   assign  _net_996 = (in_do&_net_2);
   assign  _net_997 = (in_do&_net_2);
   assign  _net_998 = (in_do&_net_2);
   assign  _net_999 = (in_do&_net_2);
   assign  _net_1000 = (in_do&_net_2);
   assign  _net_1001 = (in_do&_net_2);
   assign  _net_1002 = (in_do&_net_2);
   assign  _net_1003 = (in_do&_net_2);
   assign  _net_1004 = (in_do&_net_2);
   assign  _net_1005 = (in_do&_net_2);
   assign  _net_1006 = (in_do&_net_2);
   assign  _net_1007 = (in_do&_net_2);
   assign  _net_1008 = (in_do&_net_2);
   assign  _net_1009 = (in_do&_net_2);
   assign  _net_1010 = (in_do&_net_2);
   assign  _net_1011 = (in_do&_net_2);
   assign  _net_1012 = (in_do&_net_2);
   assign  _net_1013 = (in_do&_net_2);
   assign  _net_1014 = (in_do&_net_2);
   assign  _net_1015 = (in_do&_net_2);
   assign  _net_1016 = (in_do&_net_2);
   assign  _net_1017 = (in_do&_net_2);
   assign  _net_1018 = (in_do&_net_2);
   assign  _net_1019 = (in_do&_net_2);
   assign  _net_1020 = (in_do&_net_2);
   assign  _net_1021 = (in_do&_net_2);
   assign  _net_1022 = (in_do&_net_2);
   assign  _net_1023 = (in_do&_net_2);
   assign  _net_1024 = (in_do&_net_2);
   assign  _net_1025 = (in_do&_net_2);
   assign  _net_1026 = (in_do&_net_2);
   assign  _net_1027 = (in_do&_net_2);
   assign  _net_1028 = (in_do&_net_2);
   assign  _net_1029 = (in_do&_net_2);
   assign  _net_1030 = (in_do&_net_2);
   assign  _net_1031 = (in_do&_net_2);
   assign  _net_1032 = (in_do&_net_2);
   assign  _net_1033 = (in_do&_net_2);
   assign  _net_1034 = (in_do&_net_2);
   assign  _net_1035 = (in_do&_net_2);
   assign  _net_1036 = (in_do&_net_2);
   assign  _net_1037 = (in_do&_net_2);
   assign  _net_1038 = (in_do&_net_2);
   assign  _net_1039 = (in_do&_net_2);
   assign  _net_1040 = (in_do&_net_2);
   assign  _net_1041 = (in_do&_net_2);
   assign  _net_1042 = (in_do&_net_2);
   assign  _net_1043 = (in_do&_net_2);
   assign  _net_1044 = (in_do&_net_2);
   assign  _net_1045 = (in_do&_net_2);
   assign  _net_1046 = (in_do&_net_2);
   assign  _net_1047 = (in_do&_net_2);
   assign  _net_1048 = (in_do&_net_2);
   assign  _net_1049 = (in_do&_net_2);
   assign  _net_1050 = (in_do&_net_2);
   assign  _net_1051 = (in_do&_net_2);
   assign  _net_1052 = (in_do&_net_2);
   assign  _net_1053 = (in_do&_net_2);
   assign  _net_1054 = (in_do&_net_2);
   assign  _net_1055 = (in_do&_net_2);
   assign  _net_1056 = (in_do&_net_2);
   assign  _net_1057 = (in_do&_net_2);
   assign  _net_1058 = (in_do&_net_2);
   assign  _net_1059 = (in_do&_net_2);
   assign  _net_1060 = (in_do&_net_2);
   assign  _net_1061 = (in_do&_net_2);
   assign  _net_1062 = (in_do&_net_2);
   assign  _net_1063 = (in_do&_net_2);
   assign  _net_1064 = (in_do&_net_2);
   assign  _net_1065 = (in_do&_net_2);
   assign  _net_1066 = (in_do&_net_2);
   assign  _net_1067 = (in_do&_net_2);
   assign  _net_1068 = (in_do&_net_2);
   assign  _net_1069 = (in_do&_net_2);
   assign  _net_1070 = (in_do&_net_2);
   assign  _net_1071 = (in_do&_net_2);
   assign  _net_1072 = (in_do&_net_2);
   assign  _net_1073 = (in_do&_net_2);
   assign  _net_1074 = (in_do&_net_2);
   assign  _net_1075 = (in_do&_net_2);
   assign  _net_1076 = (in_do&_net_2);
   assign  _net_1077 = (in_do&_net_2);
   assign  _net_1078 = (in_do&_net_2);
   assign  _net_1079 = (in_do&_net_2);
   assign  _net_1080 = (in_do&_net_2);
   assign  _net_1081 = (in_do&_net_2);
   assign  _net_1082 = (in_do&_net_2);
   assign  _net_1083 = (in_do&_net_2);
   assign  _net_1084 = (in_do&_net_2);
   assign  _net_1085 = (in_do&_net_2);
   assign  _net_1086 = (in_do&_net_2);
   assign  _net_1087 = (in_do&_net_2);
   assign  _net_1088 = (in_do&_net_2);
   assign  _net_1089 = (in_do&_net_2);
   assign  _net_1090 = (in_do&_net_2);
   assign  _net_1091 = (in_do&_net_2);
   assign  _net_1092 = (in_do&_net_2);
   assign  _net_1093 = (in_do&_net_2);
   assign  _net_1094 = (in_do&_net_2);
   assign  _net_1095 = (in_do&_net_2);
   assign  _net_1096 = (in_do&_net_2);
   assign  _net_1097 = (in_do&_net_2);
   assign  _net_1098 = (in_do&_net_2);
   assign  _net_1099 = (in_do&_net_2);
   assign  _net_1100 = (in_do&_net_2);
   assign  _net_1101 = (in_do&_net_2);
   assign  _net_1102 = (in_do&_net_2);
   assign  _net_1103 = (in_do&_net_2);
   assign  _net_1104 = (in_do&_net_2);
   assign  _net_1105 = (in_do&_net_2);
   assign  _net_1106 = (in_do&_net_2);
   assign  _net_1107 = (in_do&_net_2);
   assign  _net_1108 = (in_do&_net_2);
   assign  _net_1109 = (in_do&_net_2);
   assign  _net_1110 = (in_do&_net_2);
   assign  _net_1111 = (in_do&_net_2);
   assign  _net_1112 = (in_do&_net_2);
   assign  _net_1113 = (in_do&_net_2);
   assign  _net_1114 = (in_do&_net_2);
   assign  _net_1115 = (in_do&_net_2);
   assign  _net_1116 = (in_do&_net_2);
   assign  _net_1117 = (in_do&_net_2);
   assign  _net_1118 = (in_do&_net_2);
   assign  _net_1119 = (in_do&_net_2);
   assign  _net_1120 = (in_do&_net_2);
   assign  _net_1121 = (in_do&_net_2);
   assign  _net_1122 = (in_do&_net_2);
   assign  _net_1123 = (in_do&_net_2);
   assign  _net_1124 = (in_do&_net_2);
   assign  _net_1125 = (in_do&_net_2);
   assign  _net_1126 = (in_do&_net_2);
   assign  _net_1127 = (in_do&_net_2);
   assign  _net_1128 = (in_do&_net_2);
   assign  _net_1129 = (in_do&_net_2);
   assign  _net_1130 = (in_do&_net_2);
   assign  _net_1131 = (in_do&_net_2);
   assign  _net_1132 = (in_do&_net_2);
   assign  _net_1133 = (in_do&_net_2);
   assign  _net_1134 = (in_do&_net_2);
   assign  _net_1135 = (in_do&_net_2);
   assign  _net_1136 = (in_do&_net_2);
   assign  _net_1137 = (in_do&_net_2);
   assign  _net_1138 = (in_do&_net_2);
   assign  _net_1139 = (in_do&_net_2);
   assign  _net_1140 = (in_do&_net_2);
   assign  _net_1141 = (in_do&_net_2);
   assign  _net_1142 = (in_do&_net_2);
   assign  _net_1143 = (in_do&_net_2);
   assign  _net_1144 = (in_do&_net_2);
   assign  _net_1145 = (in_do&_net_2);
   assign  _net_1146 = (in_do&_net_2);
   assign  _net_1147 = (in_do&_net_2);
   assign  _net_1148 = (in_do&_net_2);
   assign  _net_1149 = (in_do&_net_2);
   assign  _net_1150 = (in_do&_net_2);
   assign  _net_1151 = (in_do&_net_2);
   assign  _net_1152 = (in_do&_net_2);
   assign  _net_1153 = (in_do&_net_2);
   assign  _net_1154 = (in_do&_net_2);
   assign  _net_1155 = (in_do&_net_2);
   assign  _net_1156 = (in_do&_net_2);
   assign  _net_1157 = (in_do&_net_2);
   assign  _net_1158 = (in_do&_net_2);
   assign  _net_1159 = (in_do&_net_2);
   assign  _net_1160 = (in_do&_net_2);
   assign  _net_1161 = (in_do&_net_2);
   assign  _net_1162 = (in_do&_net_2);
   assign  _net_1163 = (in_do&_net_2);
   assign  _net_1164 = (in_do&_net_2);
   assign  _net_1165 = (in_do&_net_2);
   assign  _net_1166 = (in_do&_net_2);
   assign  _net_1167 = (in_do&_net_2);
   assign  _net_1168 = (in_do&_net_2);
   assign  _net_1169 = (in_do&_net_2);
   assign  _net_1170 = (in_do&_net_2);
   assign  _net_1171 = (in_do&_net_2);
   assign  _net_1172 = (in_do&_net_2);
   assign  _net_1173 = (in_do&_net_2);
   assign  _net_1174 = (in_do&_net_2);
   assign  _net_1175 = (in_do&_net_2);
   assign  _net_1176 = (in_do&_net_2);
   assign  _net_1177 = (in_do&_net_2);
   assign  _net_1178 = (in_do&_net_2);
   assign  _net_1179 = (in_do&_net_2);
   assign  _net_1180 = (in_do&_net_2);
   assign  _net_1181 = (in_do&_net_2);
   assign  _net_1182 = (in_do&_net_2);
   assign  _net_1183 = (in_do&_net_2);
   assign  _net_1184 = (in_do&_net_2);
   assign  _net_1185 = (in_do&_net_2);
   assign  _net_1186 = (in_do&_net_2);
   assign  _net_1187 = (in_do&_net_2);
   assign  _net_1188 = (in_do&_net_2);
   assign  _net_1189 = (in_do&_net_2);
   assign  _net_1190 = (in_do&_net_2);
   assign  _net_1191 = (in_do&_net_2);
   assign  _net_1192 = (in_do&_net_2);
   assign  _net_1193 = (in_do&_net_2);
   assign  _net_1194 = (in_do&_net_2);
   assign  _net_1195 = (in_do&_net_2);
   assign  _net_1196 = (in_do&_net_2);
   assign  _net_1197 = (in_do&_net_2);
   assign  _net_1198 = (in_do&_net_2);
   assign  _net_1199 = (in_do&_net_2);
   assign  _net_1200 = (in_do&_net_2);
   assign  _net_1201 = (in_do&_net_2);
   assign  _net_1202 = (in_do&_net_2);
   assign  _net_1203 = (in_do&_net_2);
   assign  _net_1204 = (in_do&_net_2);
   assign  _net_1205 = (in_do&_net_2);
   assign  _net_1206 = (in_do&_net_2);
   assign  _net_1207 = (in_do&_net_2);
   assign  _net_1208 = (in_do&_net_2);
   assign  _net_1209 = (in_do&_net_2);
   assign  _net_1210 = (in_do&_net_2);
   assign  _net_1211 = (in_do&_net_2);
   assign  _net_1212 = (in_do&_net_2);
   assign  _net_1213 = (in_do&_net_2);
   assign  _net_1214 = (in_do&_net_2);
   assign  _net_1215 = (in_do&_net_2);
   assign  _net_1216 = (in_do&_net_2);
   assign  _net_1217 = (in_do&_net_2);
   assign  _net_1218 = (in_do&_net_2);
   assign  _net_1219 = (in_do&_net_2);
   assign  _net_1220 = (in_do&_net_2);
   assign  _net_1221 = (in_do&_net_2);
   assign  _net_1222 = (in_do&_net_2);
   assign  _net_1223 = (in_do&_net_2);
   assign  _net_1224 = (in_do&_net_2);
   assign  _net_1225 = (in_do&_net_2);
   assign  _net_1226 = (in_do&_net_2);
   assign  _net_1227 = (in_do&_net_2);
   assign  _net_1228 = (in_do&_net_2);
   assign  _net_1229 = (in_do&_net_2);
   assign  _net_1230 = (in_do&_net_2);
   assign  _net_1231 = (in_do&_net_2);
   assign  _net_1232 = (in_do&_net_2);
   assign  _net_1233 = (in_do&_net_2);
   assign  _net_1234 = (in_do&_net_2);
   assign  _net_1235 = (in_do&_net_2);
   assign  _net_1236 = (in_do&_net_2);
   assign  _net_1237 = (in_do&_net_2);
   assign  _net_1238 = (in_do&_net_2);
   assign  _net_1239 = (in_do&_net_2);
   assign  _net_1240 = (in_do&_net_2);
   assign  _net_1241 = (in_do&_net_2);
   assign  _net_1242 = (in_do&_net_2);
   assign  _net_1243 = (in_do&_net_2);
   assign  _net_1244 = (in_do&_net_2);
   assign  _net_1245 = (in_do&_net_2);
   assign  _net_1246 = (in_do&_net_2);
   assign  _net_1247 = (in_do&_net_2);
   assign  _net_1248 = (in_do&_net_2);
   assign  _net_1249 = (in_do&_net_2);
   assign  _net_1250 = (in_do&_net_2);
   assign  _net_1251 = (in_do&_net_2);
   assign  _net_1252 = (in_do&_net_2);
   assign  _net_1253 = (in_do&_net_2);
   assign  _net_1254 = (in_do&_net_2);
   assign  _net_1255 = (in_do&_net_2);
   assign  _net_1256 = (in_do&_net_2);
   assign  _net_1257 = (in_do&_net_2);
   assign  _net_1258 = (in_do&_net_2);
   assign  _net_1259 = (in_do&_net_2);
   assign  _net_1260 = (in_do&_net_2);
   assign  _net_1261 = (in_do&_net_2);
   assign  _net_1262 = (in_do&_net_2);
   assign  _net_1263 = (in_do&_net_2);
   assign  _net_1264 = (in_do&_net_2);
   assign  _net_1265 = (in_do&_net_2);
   assign  _net_1266 = (in_do&_net_2);
   assign  _net_1267 = (in_do&_net_2);
   assign  _net_1268 = (in_do&_net_2);
   assign  _net_1269 = (in_do&_net_2);
   assign  _net_1270 = (in_do&_net_2);
   assign  _net_1271 = (in_do&_net_2);
   assign  _net_1272 = (in_do&_net_2);
   assign  _net_1273 = (in_do&_net_2);
   assign  _net_1274 = (in_do&_net_2);
   assign  _net_1275 = (in_do&_net_2);
   assign  _net_1276 = (in_do&_net_2);
   assign  _net_1277 = (in_do&_net_2);
   assign  _net_1278 = (in_do&_net_2);
   assign  _net_1279 = (in_do&_net_2);
   assign  _net_1280 = (in_do&_net_2);
   assign  _net_1281 = (in_do&_net_2);
   assign  _net_1282 = (in_do&_net_2);
   assign  _net_1283 = (in_do&_net_2);
   assign  _net_1284 = (in_do&_net_2);
   assign  _net_1285 = (in_do&_net_2);
   assign  _net_1286 = (in_do&_net_2);
   assign  _net_1287 = (in_do&_net_2);
   assign  _net_1288 = (in_do&_net_2);
   assign  _net_1289 = (in_do&_net_2);
   assign  _net_1290 = (in_do&_net_2);
   assign  _net_1291 = (in_do&_net_2);
   assign  _net_1292 = (in_do&_net_2);
   assign  _net_1293 = (in_do&_net_2);
   assign  _net_1294 = (in_do&_net_2);
   assign  _net_1295 = (in_do&_net_2);
   assign  _net_1296 = (in_do&_net_2);
   assign  _net_1297 = (in_do&_net_2);
   assign  _net_1298 = (in_do&_net_2);
   assign  _net_1299 = (in_do&_net_2);
   assign  _net_1300 = (in_do&_net_2);
   assign  _net_1301 = (in_do&_net_2);
   assign  _net_1302 = (in_do&_net_2);
   assign  _net_1303 = (in_do&_net_2);
   assign  _net_1304 = (in_do&_net_2);
   assign  _net_1305 = (in_do&_net_2);
   assign  _net_1306 = (in_do&_net_2);
   assign  _net_1307 = (in_do&_net_2);
   assign  _net_1308 = (in_do&_net_2);
   assign  _net_1309 = (in_do&_net_2);
   assign  _net_1310 = (in_do&_net_2);
   assign  _net_1311 = (in_do&_net_2);
   assign  _net_1312 = (in_do&_net_2);
   assign  _net_1313 = (in_do&_net_2);
   assign  _net_1314 = (in_do&_net_2);
   assign  _net_1315 = (in_do&_net_2);
   assign  _net_1316 = (in_do&_net_2);
   assign  _net_1317 = (in_do&_net_2);
   assign  _net_1318 = (in_do&_net_2);
   assign  _net_1319 = (in_do&_net_2);
   assign  _net_1320 = (in_do&_net_2);
   assign  _net_1321 = (in_do&_net_2);
   assign  _net_1322 = (in_do&_net_2);
   assign  _net_1323 = (in_do&_net_2);
   assign  _net_1324 = (in_do&_net_2);
   assign  _net_1325 = (in_do&_net_2);
   assign  _net_1326 = (in_do&_net_2);
   assign  _net_1327 = (in_do&_net_2);
   assign  _net_1328 = (in_do&_net_2);
   assign  _net_1329 = (in_do&_net_2);
   assign  _net_1330 = (in_do&_net_2);
   assign  _net_1331 = (in_do&_net_2);
   assign  _net_1332 = (in_do&_net_2);
   assign  _net_1333 = (in_do&_net_2);
   assign  _net_1334 = (in_do&_net_2);
   assign  _net_1335 = (in_do&_net_2);
   assign  _net_1336 = (in_do&_net_2);
   assign  _net_1337 = (in_do&_net_2);
   assign  _net_1338 = (in_do&_net_2);
   assign  _net_1339 = (in_do&_net_2);
   assign  _net_1340 = (in_do&_net_2);
   assign  _net_1341 = (in_do&_net_2);
   assign  _net_1342 = (in_do&_net_2);
   assign  _net_1343 = (in_do&_net_2);
   assign  _net_1344 = (in_do&_net_2);
   assign  _net_1345 = (in_do&_net_2);
   assign  _net_1346 = (in_do&_net_2);
   assign  _net_1347 = (in_do&_net_2);
   assign  _net_1348 = (in_do&_net_2);
   assign  _net_1349 = (in_do&_net_2);
   assign  _net_1350 = (in_do&_net_2);
   assign  _net_1351 = (in_do&_net_2);
   assign  _net_1352 = (in_do&_net_2);
   assign  _net_1353 = (in_do&_net_2);
   assign  _net_1354 = (in_do&_net_2);
   assign  _net_1355 = (in_do&_net_2);
   assign  _net_1356 = (in_do&_net_2);
   assign  _net_1357 = (in_do&_net_2);
   assign  _net_1358 = (in_do&_net_2);
   assign  _net_1359 = (in_do&_net_2);
   assign  _net_1360 = (in_do&_net_2);
   assign  _net_1361 = (in_do&_net_2);
   assign  _net_1362 = (in_do&_net_2);
   assign  _net_1363 = (in_do&_net_2);
   assign  _net_1364 = (in_do&_net_2);
   assign  _net_1365 = (in_do&_net_2);
   assign  _net_1366 = (in_do&_net_2);
   assign  _net_1367 = (in_do&_net_2);
   assign  _net_1368 = (in_do&_net_2);
   assign  _net_1369 = (in_do&_net_2);
   assign  _net_1370 = (in_do&_net_2);
   assign  _net_1371 = (in_do&_net_2);
   assign  _net_1372 = (in_do&_net_2);
   assign  _net_1373 = (in_do&_net_2);
   assign  _net_1374 = (in_do&_net_2);
   assign  _net_1375 = (in_do&_net_2);
   assign  _net_1376 = (in_do&_net_2);
   assign  _net_1377 = (in_do&_net_2);
   assign  _net_1378 = (in_do&_net_2);
   assign  _net_1379 = (in_do&_net_2);
   assign  _net_1380 = (in_do&_net_2);
   assign  _net_1381 = (in_do&_net_2);
   assign  _net_1382 = (in_do&_net_2);
   assign  _net_1383 = (in_do&_net_2);
   assign  _net_1384 = (in_do&_net_2);
   assign  _net_1385 = (in_do&_net_2);
   assign  _net_1386 = (in_do&_net_2);
   assign  _net_1387 = (in_do&_net_2);
   assign  _net_1388 = (in_do&_net_2);
   assign  _net_1389 = (in_do&_net_2);
   assign  _net_1390 = (in_do&_net_2);
   assign  _net_1391 = (in_do&_net_2);
   assign  _net_1392 = (in_do&_net_2);
   assign  _net_1393 = (in_do&_net_2);
   assign  _net_1394 = (in_do&_net_2);
   assign  _net_1395 = (in_do&_net_2);
   assign  _net_1396 = (in_do&_net_2);
   assign  _net_1397 = (in_do&_net_2);
   assign  _net_1398 = (in_do&_net_2);
   assign  _net_1399 = (in_do&_net_2);
   assign  _net_1400 = (in_do&_net_2);
   assign  _net_1401 = (in_do&_net_2);
   assign  _net_1402 = (in_do&_net_2);
   assign  _net_1403 = (in_do&_net_2);
   assign  _net_1404 = (in_do&_net_2);
   assign  _net_1405 = (in_do&_net_2);
   assign  _net_1406 = (in_do&_net_2);
   assign  _net_1407 = (in_do&_net_2);
   assign  _net_1408 = (in_do&_net_2);
   assign  _net_1409 = (in_do&_net_2);
   assign  _net_1410 = (in_do&_net_2);
   assign  _net_1411 = (in_do&_net_2);
   assign  _net_1412 = (in_do&_net_2);
   assign  _net_1413 = (in_do&_net_2);
   assign  _net_1414 = (in_do&_net_2);
   assign  _net_1415 = (in_do&_net_2);
   assign  _net_1416 = (in_do&_net_2);
   assign  _net_1417 = (in_do&_net_2);
   assign  _net_1418 = (in_do&_net_2);
   assign  _net_1419 = (in_do&_net_2);
   assign  _net_1420 = (in_do&_net_2);
   assign  _net_1421 = (in_do&_net_2);
   assign  _net_1422 = (in_do&_net_2);
   assign  _net_1423 = (in_do&_net_2);
   assign  _net_1424 = (in_do&_net_2);
   assign  _net_1425 = (in_do&_net_2);
   assign  _net_1426 = (in_do&_net_2);
   assign  _net_1427 = (in_do&_net_2);
   assign  _net_1428 = (in_do&_net_2);
   assign  _net_1429 = (in_do&_net_2);
   assign  _net_1430 = (in_do&_net_2);
   assign  _net_1431 = (in_do&_net_2);
   assign  _net_1432 = (in_do&_net_2);
   assign  _net_1433 = (in_do&_net_2);
   assign  _net_1434 = (in_do&_net_2);
   assign  _net_1435 = (in_do&_net_2);
   assign  _net_1436 = (in_do&_net_2);
   assign  _net_1437 = (in_do&_net_2);
   assign  _net_1438 = (in_do&_net_2);
   assign  _net_1439 = (in_do&_net_2);
   assign  _net_1440 = (in_do&_net_2);
   assign  _net_1441 = (in_do&_net_2);
   assign  _net_1442 = (in_do&_net_2);
   assign  _net_1443 = (in_do&_net_2);
   assign  _net_1444 = (in_do&_net_2);
   assign  _net_1445 = (in_do&_net_2);
   assign  _net_1446 = (in_do&_net_2);
   assign  _net_1447 = (in_do&_net_2);
   assign  _net_1448 = (in_do&_net_2);
   assign  _net_1449 = (in_do&_net_2);
   assign  _net_1450 = (in_do&_net_2);
   assign  _net_1451 = (in_do&_net_2);
   assign  _net_1452 = (in_do&_net_2);
   assign  _net_1453 = (in_do&_net_2);
   assign  _net_1454 = (in_do&_net_2);
   assign  _net_1455 = (in_do&_net_2);
   assign  _net_1456 = (in_do&_net_2);
   assign  _net_1457 = (in_do&_net_2);
   assign  _net_1458 = (in_do&_net_2);
   assign  _net_1459 = (in_do&_net_2);
   assign  _net_1460 = (in_do&_net_2);
   assign  _net_1461 = (in_do&_net_2);
   assign  _net_1462 = (in_do&_net_2);
   assign  _net_1463 = (in_do&_net_2);
   assign  _net_1464 = (in_do&_net_2);
   assign  _net_1465 = (in_do&_net_2);
   assign  _net_1466 = (in_do&_net_2);
   assign  _net_1467 = (in_do&_net_2);
   assign  _net_1468 = (in_do&_net_2);
   assign  _net_1469 = (in_do&_net_2);
   assign  _net_1470 = (in_do&_net_2);
   assign  _net_1471 = (in_do&_net_2);
   assign  _net_1472 = (in_do&_net_2);
   assign  _net_1473 = (in_do&_net_2);
   assign  _net_1474 = (in_do&_net_2);
   assign  _net_1475 = (in_do&_net_2);
   assign  _net_1476 = (in_do&_net_2);
   assign  _net_1477 = (in_do&_net_2);
   assign  _net_1478 = (in_do&_net_2);
   assign  _net_1479 = (in_do&_net_2);
   assign  _net_1480 = (in_do&_net_2);
   assign  _net_1481 = (in_do&_net_2);
   assign  _net_1482 = (in_do&_net_2);
   assign  _net_1483 = (in_do&_net_2);
   assign  _net_1484 = (in_do&_net_2);
   assign  _net_1485 = (in_do&_net_2);
   assign  _net_1486 = (in_do&_net_2);
   assign  _net_1487 = (in_do&_net_2);
   assign  _net_1488 = (in_do&_net_2);
   assign  _net_1489 = (in_do&_net_2);
   assign  _net_1490 = (in_do&_net_2);
   assign  _net_1491 = (in_do&_net_2);
   assign  _net_1492 = (in_do&_net_2);
   assign  _net_1493 = (in_do&_net_2);
   assign  _net_1494 = (in_do&_net_2);
   assign  _net_1495 = (in_do&_net_2);
   assign  _net_1496 = (in_do&_net_2);
   assign  _net_1497 = (in_do&_net_2);
   assign  _net_1498 = (in_do&_net_2);
   assign  _net_1499 = (in_do&_net_2);
   assign  _net_1500 = (in_do&_net_2);
   assign  _net_1501 = (in_do&_net_2);
   assign  _net_1502 = (in_do&_net_2);
   assign  _net_1503 = (in_do&_net_2);
   assign  _net_1504 = (in_do&_net_2);
   assign  _net_1505 = (in_do&_net_2);
   assign  _net_1506 = (in_do&_net_2);
   assign  _net_1507 = (in_do&_net_2);
   assign  _net_1508 = (in_do&_net_2);
   assign  _net_1509 = (in_do&_net_2);
   assign  _net_1510 = (in_do&_net_2);
   assign  _net_1511 = (in_do&_net_2);
   assign  _net_1512 = (in_do&_net_2);
   assign  _net_1513 = (in_do&_net_2);
   assign  _net_1514 = (in_do&_net_2);
   assign  _net_1515 = (in_do&_net_2);
   assign  _net_1516 = (in_do&_net_2);
   assign  _net_1517 = (in_do&_net_2);
   assign  _net_1518 = (in_do&_net_2);
   assign  _net_1519 = (in_do&_net_2);
   assign  _net_1520 = (in_do&_net_2);
   assign  _net_1521 = (in_do&_net_2);
   assign  _net_1522 = (in_do&_net_2);
   assign  _net_1523 = (in_do&_net_2);
   assign  _net_1524 = (in_do&_net_2);
   assign  _net_1525 = (in_do&_net_2);
   assign  _net_1526 = (in_do&_net_2);
   assign  _net_1527 = (in_do&_net_2);
   assign  _net_1528 = (in_do&_net_2);
   assign  _net_1529 = (in_do&_net_2);
   assign  _net_1530 = (in_do&_net_2);
   assign  _net_1531 = (in_do&_net_2);
   assign  _net_1532 = (in_do&_net_2);
   assign  _net_1533 = (in_do&_net_2);
   assign  _net_1534 = (in_do&_net_2);
   assign  _net_1535 = (in_do&_net_2);
   assign  _net_1536 = (in_do&_net_2);
   assign  _net_1537 = (in_do&_net_2);
   assign  _net_1538 = (in_do&_net_2);
   assign  _net_1539 = (in_do&_net_2);
   assign  _net_1540 = (in_do&_net_2);
   assign  _net_1541 = (in_do&_net_2);
   assign  _net_1542 = (in_do&_net_2);
   assign  _net_1543 = (in_do&_net_2);
   assign  _net_1544 = (in_do&_net_2);
   assign  _net_1545 = (in_do&_net_2);
   assign  _net_1546 = (in_do&_net_2);
   assign  _net_1547 = (in_do&_net_2);
   assign  _net_1548 = (in_do&_net_2);
   assign  _net_1549 = (in_do&_net_2);
   assign  _net_1550 = (in_do&_net_2);
   assign  _net_1551 = (in_do&_net_2);
   assign  _net_1552 = (in_do&_net_2);
   assign  _net_1553 = (in_do&_net_2);
   assign  _net_1554 = (in_do&_net_2);
   assign  _net_1555 = (in_do&_net_2);
   assign  _net_1556 = (in_do&_net_2);
   assign  _net_1557 = (in_do&_net_2);
   assign  _net_1558 = (in_do&_net_2);
   assign  _net_1559 = (in_do&_net_2);
   assign  _net_1560 = (in_do&_net_2);
   assign  _net_1561 = (in_do&_net_2);
   assign  _net_1562 = (in_do&_net_2);
   assign  _net_1563 = (in_do&_net_2);
   assign  _net_1564 = (in_do&_net_2);
   assign  _net_1565 = (in_do&_net_2);
   assign  _net_1566 = (in_do&_net_2);
   assign  _net_1567 = (in_do&_net_2);
   assign  _net_1568 = (in_do&_net_2);
   assign  _net_1569 = (in_do&_net_2);
   assign  _net_1570 = (in_do&_net_2);
   assign  _net_1571 = (in_do&_net_2);
   assign  _net_1572 = (in_do&_net_2);
   assign  _net_1573 = (in_do&_net_2);
   assign  _net_1574 = (in_do&_net_2);
   assign  _net_1575 = (in_do&_net_2);
   assign  _net_1576 = (in_do&_net_2);
   assign  _net_1577 = (in_do&_net_2);
   assign  _net_1578 = (in_do&_net_2);
   assign  _net_1579 = (in_do&_net_2);
   assign  _net_1580 = (in_do&_net_2);
   assign  _net_1581 = (in_do&_net_2);
   assign  _net_1582 = (in_do&_net_2);
   assign  _net_1583 = (in_do&_net_2);
   assign  _net_1584 = (in_do&_net_2);
   assign  _net_1585 = (in_do&_net_2);
   assign  _net_1586 = (in_do&_net_2);
   assign  _net_1587 = (in_do&_net_2);
   assign  _net_1588 = (in_do&_net_2);
   assign  _net_1589 = (in_do&_net_2);
   assign  _net_1590 = (in_do&_net_2);
   assign  _net_1591 = (in_do&_net_2);
   assign  _net_1592 = (in_do&_net_2);
   assign  _net_1593 = (in_do&_net_2);
   assign  _net_1594 = (in_do&_net_2);
   assign  _net_1595 = (in_do&_net_2);
   assign  _net_1596 = (in_do&_net_2);
   assign  _net_1597 = (in_do&_net_2);
   assign  _net_1598 = (in_do&_net_2);
   assign  _net_1599 = (in_do&_net_2);
   assign  _net_1600 = (in_do&_net_2);
   assign  _net_1601 = (in_do&_net_2);
   assign  _net_1602 = (in_do&_net_2);
   assign  _net_1603 = (in_do&_net_2);
   assign  _net_1604 = (in_do&_net_2);
   assign  _net_1605 = (in_do&_net_2);
   assign  _net_1606 = (in_do&_net_2);
   assign  _net_1607 = (in_do&_net_2);
   assign  _net_1608 = (in_do&_net_2);
   assign  _net_1609 = (in_do&_net_2);
   assign  _net_1610 = (in_do&_net_2);
   assign  _net_1611 = (in_do&_net_2);
   assign  _net_1612 = (in_do&_net_2);
   assign  _net_1613 = (in_do&_net_2);
   assign  _net_1614 = (in_do&_net_2);
   assign  _net_1615 = (in_do&_net_2);
   assign  _net_1616 = (in_do&_net_2);
   assign  _net_1617 = (in_do&_net_2);
   assign  _net_1618 = (in_do&_net_2);
   assign  _net_1619 = (in_do&_net_2);
   assign  _net_1620 = (in_do&_net_2);
   assign  _net_1621 = (in_do&_net_2);
   assign  _net_1622 = (in_do&_net_2);
   assign  _net_1623 = (in_do&_net_2);
   assign  _net_1624 = (in_do&_net_2);
   assign  _net_1625 = (in_do&_net_2);
   assign  _net_1626 = (in_do&_net_2);
   assign  _net_1627 = (in_do&_net_2);
   assign  _net_1628 = (in_do&_net_2);
   assign  _net_1629 = (in_do&_net_2);
   assign  _net_1630 = (in_do&_net_2);
   assign  _net_1631 = (in_do&_net_2);
   assign  _net_1632 = (in_do&_net_2);
   assign  _net_1633 = (in_do&_net_2);
   assign  _net_1634 = (in_do&_net_2);
   assign  _net_1635 = (in_do&_net_2);
   assign  _net_1636 = (in_do&_net_2);
   assign  _net_1637 = (in_do&_net_2);
   assign  _net_1638 = (in_do&_net_2);
   assign  _net_1639 = (in_do&_net_2);
   assign  _net_1640 = (in_do&_net_2);
   assign  _net_1641 = (in_do&_net_2);
   assign  _net_1642 = (in_do&_net_2);
   assign  _net_1643 = (in_do&_net_2);
   assign  _net_1644 = (in_do&_net_2);
   assign  _net_1645 = (in_do&_net_2);
   assign  _net_1646 = (in_do&_net_2);
   assign  _net_1647 = (in_do&_net_2);
   assign  _net_1648 = (in_do&_net_2);
   assign  _net_1649 = (in_do&_net_2);
   assign  _net_1650 = (in_do&_net_2);
   assign  _net_1651 = (in_do&_net_2);
   assign  _net_1652 = (in_do&_net_2);
   assign  _net_1653 = (in_do&_net_2);
   assign  _net_1654 = (in_do&_net_2);
   assign  _net_1655 = (in_do&_net_2);
   assign  _net_1656 = (in_do&_net_2);
   assign  _net_1657 = (in_do&_net_2);
   assign  _net_1658 = (in_do&_net_2);
   assign  _net_1659 = (in_do&_net_2);
   assign  _net_1660 = (in_do&_net_2);
   assign  _net_1661 = (in_do&_net_2);
   assign  _net_1662 = (in_do&_net_2);
   assign  _net_1663 = (in_do&_net_2);
   assign  _net_1664 = (in_do&_net_2);
   assign  _net_1665 = (in_do&_net_2);
   assign  _net_1666 = (in_do&_net_2);
   assign  _net_1667 = (in_do&_net_2);
   assign  _net_1668 = (in_do&_net_2);
   assign  _net_1669 = (in_do&_net_2);
   assign  _net_1670 = (in_do&_net_2);
   assign  _net_1671 = (in_do&_net_2);
   assign  _net_1672 = (in_do&_net_2);
   assign  _net_1673 = (in_do&_net_2);
   assign  _net_1674 = (in_do&_net_2);
   assign  _net_1675 = (in_do&_net_2);
   assign  _net_1676 = (in_do&_net_2);
   assign  _net_1677 = (in_do&_net_2);
   assign  _net_1678 = (in_do&_net_2);
   assign  _net_1679 = (in_do&_net_2);
   assign  _net_1680 = (in_do&_net_2);
   assign  _net_1681 = (in_do&_net_2);
   assign  _net_1682 = (in_do&_net_2);
   assign  _net_1683 = (in_do&_net_2);
   assign  _net_1684 = (in_do&_net_2);
   assign  _net_1685 = (in_do&_net_2);
   assign  _net_1686 = (in_do&_net_2);
   assign  _net_1687 = (in_do&_net_2);
   assign  _net_1688 = (in_do&_net_2);
   assign  _net_1689 = (in_do&_net_2);
   assign  _net_1690 = (in_do&_net_2);
   assign  _net_1691 = (in_do&_net_2);
   assign  _net_1692 = (in_do&_net_2);
   assign  _net_1693 = (in_do&_net_2);
   assign  _net_1694 = (in_do&_net_2);
   assign  _net_1695 = (in_do&_net_2);
   assign  _net_1696 = (in_do&_net_2);
   assign  _net_1697 = (in_do&_net_2);
   assign  _net_1698 = (in_do&_net_2);
   assign  _net_1699 = (in_do&_net_2);
   assign  _net_1700 = (in_do&_net_2);
   assign  _net_1701 = (in_do&_net_2);
   assign  _net_1702 = (in_do&_net_2);
   assign  _net_1703 = (in_do&_net_2);
   assign  _net_1704 = (in_do&_net_2);
   assign  _net_1705 = (in_do&_net_2);
   assign  _net_1706 = (in_do&_net_2);
   assign  _net_1707 = (in_do&_net_2);
   assign  _net_1708 = (in_do&_net_2);
   assign  _net_1709 = (in_do&_net_2);
   assign  _net_1710 = (in_do&_net_2);
   assign  _net_1711 = (in_do&_net_2);
   assign  _net_1712 = (in_do&_net_2);
   assign  _net_1713 = (in_do&_net_2);
   assign  _net_1714 = (in_do&_net_2);
   assign  _net_1715 = (in_do&_net_2);
   assign  _net_1716 = (in_do&_net_2);
   assign  _net_1717 = (in_do&_net_2);
   assign  _net_1718 = (in_do&_net_2);
   assign  _net_1719 = (in_do&_net_2);
   assign  _net_1720 = (in_do&_net_2);
   assign  _net_1721 = (in_do&_net_2);
   assign  _net_1722 = (in_do&_net_2);
   assign  _net_1723 = (in_do&_net_2);
   assign  _net_1724 = (in_do&_net_2);
   assign  _net_1725 = (in_do&_net_2);
   assign  _net_1726 = (in_do&_net_2);
   assign  _net_1727 = (in_do&_net_2);
   assign  _net_1728 = (in_do&_net_2);
   assign  _net_1729 = (in_do&_net_2);
   assign  _net_1730 = (in_do&_net_2);
   assign  _net_1731 = (in_do&_net_2);
   assign  _net_1732 = (in_do&_net_2);
   assign  _net_1733 = (in_do&_net_2);
   assign  _net_1734 = (in_do&_net_2);
   assign  _net_1735 = (in_do&_net_2);
   assign  _net_1736 = (in_do&_net_2);
   assign  _net_1737 = (in_do&_net_2);
   assign  _net_1738 = (in_do&_net_2);
   assign  _net_1739 = (in_do&_net_2);
   assign  _net_1740 = (in_do&_net_2);
   assign  _net_1741 = (in_do&_net_2);
   assign  _net_1742 = (in_do&_net_2);
   assign  _net_1743 = (in_do&_net_2);
   assign  _net_1744 = (in_do&_net_2);
   assign  _net_1745 = (in_do&_net_2);
   assign  _net_1746 = (in_do&_net_2);
   assign  _net_1747 = (in_do&_net_2);
   assign  _net_1748 = (in_do&_net_2);
   assign  _net_1749 = (in_do&_net_2);
   assign  _net_1750 = (in_do&_net_2);
   assign  _net_1751 = (in_do&_net_2);
   assign  _net_1752 = (in_do&_net_2);
   assign  _net_1753 = (in_do&_net_2);
   assign  _net_1754 = (in_do&_net_2);
   assign  _net_1755 = (in_do&_net_2);
   assign  _net_1756 = (in_do&_net_2);
   assign  _net_1757 = (in_do&_net_2);
   assign  _net_1758 = (in_do&_net_2);
   assign  _net_1759 = (in_do&_net_2);
   assign  _net_1760 = (in_do&_net_2);
   assign  _net_1761 = (in_do&_net_2);
   assign  _net_1762 = (in_do&_net_2);
   assign  _net_1763 = (in_do&_net_2);
   assign  _net_1764 = (in_do&_net_2);
   assign  _net_1765 = (in_do&_net_2);
   assign  _net_1766 = (in_do&_net_2);
   assign  _net_1767 = (in_do&_net_2);
   assign  _net_1768 = (in_do&_net_2);
   assign  _net_1769 = (in_do&_net_2);
   assign  _net_1770 = (in_do&_net_2);
   assign  _net_1771 = (in_do&_net_2);
   assign  _net_1772 = (in_do&_net_2);
   assign  _net_1773 = (in_do&_net_2);
   assign  _net_1774 = (in_do&_net_2);
   assign  _net_1775 = (in_do&_net_2);
   assign  _net_1776 = (in_do&_net_2);
   assign  _net_1777 = (in_do&_net_2);
   assign  _net_1778 = (in_do&_net_2);
   assign  _net_1779 = (in_do&_net_2);
   assign  _net_1780 = (in_do&_net_2);
   assign  _net_1781 = (in_do&_net_2);
   assign  _net_1782 = (in_do&_net_2);
   assign  _net_1783 = (in_do&_net_2);
   assign  _net_1784 = (in_do&_net_2);
   assign  _net_1785 = (in_do&_net_2);
   assign  _net_1786 = (in_do&_net_2);
   assign  _net_1787 = (in_do&_net_2);
   assign  _net_1788 = (in_do&_net_2);
   assign  _net_1789 = (in_do&_net_2);
   assign  _net_1790 = (in_do&_net_2);
   assign  _net_1791 = (in_do&_net_2);
   assign  _net_1792 = (in_do&_net_2);
   assign  _net_1793 = (in_do&_net_2);
   assign  _net_1794 = (in_do&_net_2);
   assign  _net_1795 = (in_do&_net_2);
   assign  _net_1796 = (in_do&_net_2);
   assign  _net_1797 = (in_do&_net_2);
   assign  _net_1798 = (in_do&_net_2);
   assign  _net_1799 = (in_do&_net_2);
   assign  _net_1800 = (in_do&_net_2);
   assign  _net_1801 = (in_do&_net_2);
   assign  _net_1802 = (in_do&_net_2);
   assign  _net_1803 = (in_do&_net_2);
   assign  _net_1804 = (in_do&_net_2);
   assign  _net_1805 = (in_do&_net_2);
   assign  _net_1806 = (in_do&_net_2);
   assign  _net_1807 = (in_do&_net_2);
   assign  _net_1808 = (in_do&_net_2);
   assign  _net_1809 = (in_do&_net_2);
   assign  _net_1810 = (in_do&_net_2);
   assign  _net_1811 = (in_do&_net_2);
   assign  _net_1812 = (in_do&_net_2);
   assign  _net_1813 = (in_do&_net_2);
   assign  _net_1814 = (in_do&_net_2);
   assign  _net_1815 = (in_do&_net_2);
   assign  _net_1816 = (in_do&_net_2);
   assign  _net_1817 = (in_do&_net_2);
   assign  _net_1818 = (in_do&_net_2);
   assign  _net_1819 = (in_do&_net_2);
   assign  _net_1820 = (in_do&_net_2);
   assign  _net_1821 = (in_do&_net_2);
   assign  _net_1822 = (in_do&_net_2);
   assign  _net_1823 = (in_do&_net_2);
   assign  _net_1824 = (in_do&_net_2);
   assign  _net_1825 = (in_do&_net_2);
   assign  _net_1826 = (in_do&_net_2);
   assign  _net_1827 = (in_do&_net_2);
   assign  _net_1828 = (in_do&_net_2);
   assign  _net_1829 = (in_do&_net_2);
   assign  _net_1830 = (in_do&_net_2);
   assign  _net_1831 = (in_do&_net_2);
   assign  _net_1832 = (in_do&_net_2);
   assign  _net_1833 = (in_do&_net_2);
   assign  _net_1834 = (in_do&_net_2);
   assign  _net_1835 = (in_do&_net_2);
   assign  _net_1836 = (in_do&_net_2);
   assign  _net_1837 = (in_do&_net_2);
   assign  _net_1838 = (in_do&_net_2);
   assign  _net_1839 = (in_do&_net_2);
   assign  _net_1840 = (in_do&_net_2);
   assign  _net_1841 = (in_do&_net_2);
   assign  _net_1842 = (in_do&_net_2);
   assign  _net_1843 = (in_do&_net_2);
   assign  _net_1844 = (in_do&_net_2);
   assign  _net_1845 = (in_do&_net_2);
   assign  _net_1846 = (in_do&_net_2);
   assign  _net_1847 = (in_do&_net_2);
   assign  _net_1848 = (in_do&_net_2);
   assign  _net_1849 = (in_do&_net_2);
   assign  _net_1850 = (in_do&_net_2);
   assign  _net_1851 = (in_do&_net_2);
   assign  _net_1852 = (in_do&_net_2);
   assign  _net_1853 = (in_do&_net_2);
   assign  _net_1854 = (in_do&_net_2);
   assign  _net_1855 = (in_do&_net_2);
   assign  _net_1856 = (in_do&_net_2);
   assign  _net_1857 = (in_do&_net_2);
   assign  _net_1858 = (in_do&_net_2);
   assign  _net_1859 = (in_do&_net_2);
   assign  _net_1860 = (in_do&_net_2);
   assign  _net_1861 = (in_do&_net_2);
   assign  _net_1862 = (in_do&_net_2);
   assign  _net_1863 = (in_do&_net_2);
   assign  _net_1864 = (in_do&_net_2);
   assign  _net_1865 = (in_do&_net_2);
   assign  _net_1866 = (in_do&_net_2);
   assign  _net_1867 = (in_do&_net_2);
   assign  _net_1868 = (in_do&_net_2);
   assign  _net_1869 = (in_do&_net_2);
   assign  _net_1870 = (in_do&_net_2);
   assign  _net_1871 = (in_do&_net_2);
   assign  _net_1872 = (in_do&_net_2);
   assign  _net_1873 = (in_do&_net_2);
   assign  _net_1874 = (in_do&_net_2);
   assign  _net_1875 = (in_do&_net_2);
   assign  _net_1876 = (in_do&_net_2);
   assign  _net_1877 = (in_do&_net_2);
   assign  _net_1878 = (in_do&_net_2);
   assign  _net_1879 = (in_do&_net_2);
   assign  _net_1880 = (in_do&_net_2);
   assign  _net_1881 = (in_do&_net_2);
   assign  _net_1882 = (in_do&_net_2);
   assign  _net_1883 = (in_do&_net_2);
   assign  _net_1884 = (in_do&_net_2);
   assign  _net_1885 = (in_do&_net_2);
   assign  _net_1886 = (in_do&_net_2);
   assign  _net_1887 = (in_do&_net_2);
   assign  _net_1888 = (in_do&_net_2);
   assign  _net_1889 = (in_do&_net_2);
   assign  _net_1890 = (in_do&_net_2);
   assign  _net_1891 = (in_do&_net_2);
   assign  _net_1892 = (in_do&_net_2);
   assign  _net_1893 = (in_do&_net_2);
   assign  _net_1894 = (in_do&_net_2);
   assign  _net_1895 = (in_do&_net_2);
   assign  _net_1896 = (in_do&_net_2);
   assign  _net_1897 = (in_do&_net_2);
   assign  _net_1898 = (in_do&_net_2);
   assign  _net_1899 = (in_do&_net_2);
   assign  _net_1900 = (in_do&_net_2);
   assign  _net_1901 = (in_do&_net_2);
   assign  _net_1902 = (in_do&_net_2);
   assign  _net_1903 = (in_do&_net_2);
   assign  _net_1904 = (in_do&_net_2);
   assign  _net_1905 = (in_do&_net_2);
   assign  _net_1906 = (in_do&_net_2);
   assign  _net_1907 = (in_do&_net_2);
   assign  _net_1908 = (in_do&_net_2);
   assign  _net_1909 = (in_do&_net_2);
   assign  _net_1910 = (in_do&_net_2);
   assign  _net_1911 = (in_do&_net_2);
   assign  _net_1912 = (in_do&_net_2);
   assign  _net_1913 = (in_do&_net_2);
   assign  _net_1914 = (in_do&_net_2);
   assign  _net_1915 = (in_do&_net_2);
   assign  _net_1916 = (in_do&_net_2);
   assign  _net_1917 = (in_do&_net_2);
   assign  _net_1918 = (in_do&_net_2);
   assign  _net_1919 = (in_do&_net_2);
   assign  _net_1920 = (in_do&_net_2);
   assign  _net_1921 = (in_do&_net_2);
   assign  _net_1922 = (in_do&_net_2);
   assign  _net_1923 = (in_do&_net_2);
   assign  _net_1924 = (in_do&_net_2);
   assign  _net_1925 = (in_do&_net_2);
   assign  _net_1926 = (in_do&_net_2);
   assign  _net_1927 = (in_do&_net_2);
   assign  _net_1928 = (in_do&_net_2);
   assign  _net_1929 = (in_do&_net_2);
   assign  _net_1930 = (in_do&_net_2);
   assign  _net_1931 = (in_do&_net_2);
   assign  _net_1932 = (in_do&_net_2);
   assign  _net_1933 = (in_do&_net_2);
   assign  _net_1934 = (in_do&_net_2);
   assign  _net_1935 = (in_do&_net_2);
   assign  _net_1936 = (in_do&_net_2);
   assign  _net_1937 = (in_do&_net_2);
   assign  _net_1938 = (in_do&_net_2);
   assign  _net_1939 = (in_do&_net_2);
   assign  _net_1940 = (in_do&_net_2);
   assign  _net_1941 = (in_do&_net_2);
   assign  _net_1942 = (in_do&_net_2);
   assign  _net_1943 = (in_do&_net_2);
   assign  _net_1944 = (in_do&_net_2);
   assign  _net_1945 = (in_do&_net_2);
   assign  _net_1946 = (in_do&_net_2);
   assign  _net_1947 = (in_do&_net_2);
   assign  _net_1948 = (in_do&_net_2);
   assign  _net_1949 = (in_do&_net_2);
   assign  _net_1950 = (in_do&_net_2);
   assign  _net_1951 = (in_do&_net_2);
   assign  _net_1952 = (in_do&_net_2);
   assign  _net_1953 = (in_do&_net_2);
   assign  _net_1954 = (in_do&_net_2);
   assign  _net_1955 = (in_do&_net_2);
   assign  _net_1956 = (in_do&_net_2);
   assign  _net_1957 = (in_do&_net_2);
   assign  _net_1958 = (in_do&_net_2);
   assign  _net_1959 = (in_do&_net_2);
   assign  _net_1960 = (in_do&_net_2);
   assign  _net_1961 = (in_do&_net_2);
   assign  _net_1962 = (in_do&_net_2);
   assign  _net_1963 = (in_do&_net_2);
   assign  _net_1964 = (in_do&_net_2);
   assign  _net_1965 = (in_do&_net_2);
   assign  _net_1966 = (in_do&_net_2);
   assign  _net_1967 = (in_do&_net_2);
   assign  _net_1968 = (in_do&_net_2);
   assign  _net_1969 = (in_do&_net_2);
   assign  _net_1970 = (in_do&_net_2);
   assign  _net_1971 = (in_do&_net_2);
   assign  _net_1972 = (in_do&_net_2);
   assign  _net_1973 = (in_do&_net_2);
   assign  _net_1974 = (in_do&_net_2);
   assign  _net_1975 = (in_do&_net_2);
   assign  _net_1976 = (in_do&_net_2);
   assign  _net_1977 = (in_do&_net_2);
   assign  _net_1978 = (in_do&_net_2);
   assign  _net_1979 = (in_do&_net_2);
   assign  _net_1980 = (in_do&_net_2);
   assign  _net_1981 = (in_do&_net_2);
   assign  _net_1982 = (in_do&_net_2);
   assign  _net_1983 = (in_do&_net_2);
   assign  _net_1984 = (in_do&_net_2);
   assign  _net_1985 = (in_do&_net_2);
   assign  _net_1986 = (in_do&_net_2);
   assign  _net_1987 = (in_do&_net_2);
   assign  _net_1988 = (in_do&_net_2);
   assign  _net_1989 = (in_do&_net_2);
   assign  _net_1990 = (in_do&_net_2);
   assign  _net_1991 = (in_do&_net_2);
   assign  _net_1992 = (in_do&_net_2);
   assign  _net_1993 = (in_do&_net_2);
   assign  _net_1994 = (in_do&_net_2);
   assign  _net_1995 = (in_do&_net_2);
   assign  _net_1996 = (in_do&_net_2);
   assign  _net_1997 = (in_do&_net_2);
   assign  _net_1998 = (in_do&_net_2);
   assign  _net_1999 = (in_do&_net_2);
   assign  _net_2000 = (in_do&_net_2);
   assign  _net_2001 = (in_do&_net_2);
   assign  _net_2002 = (in_do&_net_2);
   assign  _net_2003 = (in_do&_net_2);
   assign  _net_2004 = (in_do&_net_2);
   assign  _net_2005 = (in_do&_net_2);
   assign  _net_2006 = (in_do&_net_2);
   assign  _net_2007 = (in_do&_net_2);
   assign  _net_2008 = (in_do&_net_2);
   assign  _net_2009 = (in_do&_net_2);
   assign  _net_2010 = (in_do&_net_2);
   assign  _net_2011 = (in_do&_net_2);
   assign  _net_2012 = (in_do&_net_2);
   assign  _net_2013 = (in_do&_net_2);
   assign  _net_2014 = (in_do&_net_2);
   assign  _net_2015 = (in_do&_net_2);
   assign  _net_2016 = (in_do&_net_2);
   assign  _net_2017 = (in_do&_net_2);
   assign  _net_2018 = (in_do&_net_2);
   assign  _net_2019 = (in_do&_net_2);
   assign  _net_2020 = (in_do&_net_2);
   assign  _net_2021 = (in_do&_net_2);
   assign  _net_2022 = (in_do&_net_2);
   assign  _net_2023 = (in_do&_net_2);
   assign  _net_2024 = (in_do&_net_2);
   assign  _net_2025 = (in_do&_net_2);
   assign  _net_2026 = (in_do&_net_2);
   assign  _net_2027 = (in_do&_net_2);
   assign  _net_2028 = (in_do&_net_2);
   assign  _net_2029 = (in_do&_net_2);
   assign  _net_2030 = (in_do&_net_2);
   assign  _net_2031 = (in_do&_net_2);
   assign  _net_2032 = (in_do&_net_2);
   assign  _net_2033 = (in_do&_net_2);
   assign  _net_2034 = (in_do&_net_2);
   assign  _net_2035 = (in_do&_net_2);
   assign  _net_2036 = (in_do&_net_2);
   assign  _net_2037 = (in_do&_net_2);
   assign  _net_2038 = (in_do&_net_2);
   assign  _net_2039 = (in_do&_net_2);
   assign  _net_2040 = (in_do&_net_2);
   assign  _net_2041 = (in_do&_net_2);
   assign  _net_2042 = (in_do&_net_2);
   assign  _net_2043 = (in_do&_net_2);
   assign  _net_2044 = (in_do&_net_2);
   assign  _net_2045 = (in_do&_net_2);
   assign  _net_2046 = (in_do&_net_2);
   assign  _net_2047 = (in_do&_net_2);
   assign  _net_2048 = (in_do&_net_2);
   assign  _net_2049 = (in_do&_net_2);
   assign  _net_2050 = (in_do&_net_2);
   assign  _net_2051 = (in_do&_net_2);
   assign  _net_2052 = (in_do&_net_2);
   assign  _net_2053 = (in_do&_net_2);
   assign  _net_2054 = (in_do&_net_2);
   assign  _net_2055 = (in_do&_net_2);
   assign  _net_2056 = (in_do&_net_2);
   assign  _net_2057 = (in_do&_net_2);
   assign  _net_2058 = (in_do&_net_2);
   assign  _net_2059 = (in_do&_net_2);
   assign  _net_2060 = (in_do&_net_2);
   assign  _net_2061 = (in_do&_net_2);
   assign  _net_2062 = (in_do&_net_2);
   assign  _net_2063 = (in_do&_net_2);
   assign  _net_2064 = (in_do&_net_2);
   assign  _net_2065 = (in_do&_net_2);
   assign  _net_2066 = (in_do&_net_2);
   assign  _net_2067 = (in_do&_net_2);
   assign  _net_2068 = (in_do&_net_2);
   assign  _net_2069 = (in_do&_net_2);
   assign  _net_2070 = (in_do&_net_2);
   assign  _net_2071 = (in_do&_net_2);
   assign  _net_2072 = (in_do&_net_2);
   assign  _net_2073 = (in_do&_net_2);
   assign  _net_2074 = (in_do&_net_2);
   assign  _net_2075 = (in_do&_net_2);
   assign  _net_2076 = (in_do&_net_2);
   assign  _net_2077 = (in_do&_net_2);
   assign  _net_2078 = (in_do&_net_2);
   assign  _net_2079 = (in_do&_net_2);
   assign  _net_2080 = (in_do&_net_2);
   assign  _net_2081 = (in_do&_net_2);
   assign  _net_2082 = (in_do&_net_2);
   assign  _net_2083 = (in_do&_net_2);
   assign  _net_2084 = (in_do&_net_2);
   assign  _net_2085 = (in_do&_net_2);
   assign  _net_2086 = (in_do&_net_2);
   assign  _net_2087 = (in_do&_net_2);
   assign  _net_2088 = (in_do&_net_2);
   assign  _net_2089 = (in_do&_net_2);
   assign  _net_2090 = (in_do&_net_2);
   assign  _net_2091 = (in_do&_net_2);
   assign  _net_2092 = (in_do&_net_2);
   assign  _net_2093 = (in_do&_net_2);
   assign  _net_2094 = (in_do&_net_2);
   assign  _net_2095 = (in_do&_net_2);
   assign  _net_2096 = (in_do&_net_2);
   assign  _net_2097 = (in_do&_net_2);
   assign  _net_2098 = (in_do&_net_2);
   assign  _net_2099 = (in_do&_net_2);
   assign  _net_2100 = (in_do&_net_2);
   assign  _net_2101 = (in_do&_net_2);
   assign  _net_2102 = (in_do&_net_2);
   assign  _net_2103 = (in_do&_net_2);
   assign  _net_2104 = (in_do&_net_2);
   assign  _net_2105 = (in_do&_net_2);
   assign  _net_2106 = (in_do&_net_2);
   assign  _net_2107 = (in_do&_net_2);
   assign  _net_2108 = (in_do&_net_2);
   assign  _net_2109 = (in_do&_net_2);
   assign  _net_2110 = (in_do&_net_2);
   assign  _net_2111 = (in_do&_net_2);
   assign  _net_2112 = (in_do&_net_2);
   assign  _net_2113 = (in_do&_net_2);
   assign  _net_2114 = (in_do&_net_2);
   assign  _net_2115 = (in_do&_net_2);
   assign  _net_2116 = (in_do&_net_2);
   assign  _net_2117 = (in_do&_net_2);
   assign  _net_2118 = (in_do&_net_2);
   assign  _net_2119 = (in_do&_net_2);
   assign  _net_2120 = (in_do&_net_2);
   assign  _net_2121 = (in_do&_net_2);
   assign  _net_2122 = (in_do&_net_2);
   assign  _net_2123 = (in_do&_net_2);
   assign  _net_2124 = (in_do&_net_2);
   assign  _net_2125 = (in_do&_net_2);
   assign  _net_2126 = (in_do&_net_2);
   assign  _net_2127 = (in_do&_net_2);
   assign  _net_2128 = (in_do&_net_2);
   assign  _net_2129 = (in_do&_net_2);
   assign  _net_2130 = (in_do&_net_2);
   assign  _net_2131 = (in_do&_net_2);
   assign  _net_2132 = (in_do&_net_2);
   assign  _net_2133 = (in_do&_net_2);
   assign  _net_2134 = (in_do&_net_2);
   assign  _net_2135 = (in_do&_net_2);
   assign  _net_2136 = (in_do&_net_2);
   assign  _net_2137 = (in_do&_net_2);
   assign  _net_2138 = (in_do&_net_2);
   assign  _net_2139 = (in_do&_net_2);
   assign  _net_2140 = (in_do&_net_2);
   assign  _net_2141 = (in_do&_net_2);
   assign  _net_2142 = (in_do&_net_2);
   assign  _net_2143 = (in_do&_net_2);
   assign  _net_2144 = (in_do&_net_2);
   assign  _net_2145 = (in_do&_net_2);
   assign  _net_2146 = (in_do&_net_2);
   assign  _net_2147 = (in_do&_net_2);
   assign  _net_2148 = (in_do&_net_2);
   assign  _net_2149 = (in_do&_net_2);
   assign  _net_2150 = (in_do&_net_2);
   assign  _net_2151 = (in_do&_net_2);
   assign  _net_2152 = (in_do&_net_2);
   assign  _net_2153 = (in_do&_net_2);
   assign  _net_2154 = (in_do&_net_2);
   assign  _net_2155 = (in_do&_net_2);
   assign  _net_2156 = (in_do&_net_2);
   assign  _net_2157 = (in_do&_net_2);
   assign  _net_2158 = (in_do&_net_2);
   assign  _net_2159 = (in_do&_net_2);
   assign  _net_2160 = (in_do&_net_2);
   assign  _net_2161 = (in_do&_net_2);
   assign  _net_2162 = (in_do&_net_2);
   assign  _net_2163 = (in_do&_net_2);
   assign  _net_2164 = (in_do&_net_2);
   assign  _net_2165 = (in_do&_net_2);
   assign  _net_2166 = (in_do&_net_2);
   assign  _net_2167 = (in_do&_net_2);
   assign  _net_2168 = (in_do&_net_2);
   assign  _net_2169 = (in_do&_net_2);
   assign  _net_2170 = (in_do&_net_2);
   assign  _net_2171 = (in_do&_net_2);
   assign  _net_2172 = (in_do&_net_2);
   assign  _net_2173 = (in_do&_net_2);
   assign  _net_2174 = (in_do&_net_2);
   assign  _net_2175 = (in_do&_net_2);
   assign  _net_2176 = (in_do&_net_2);
   assign  _net_2177 = (in_do&_net_2);
   assign  _net_2178 = (in_do&_net_2);
   assign  _net_2179 = (in_do&_net_2);
   assign  _net_2180 = (in_do&_net_2);
   assign  _net_2181 = (in_do&_net_2);
   assign  _net_2182 = (in_do&_net_2);
   assign  _net_2183 = (in_do&_net_2);
   assign  _net_2184 = (in_do&_net_2);
   assign  _net_2185 = (in_do&_net_2);
   assign  _net_2186 = (in_do&_net_2);
   assign  _net_2187 = (in_do&_net_2);
   assign  _net_2188 = (in_do&_net_2);
   assign  _net_2189 = (in_do&_net_2);
   assign  _net_2190 = (in_do&_net_2);
   assign  _net_2191 = (in_do&_net_2);
   assign  _net_2192 = (in_do&_net_2);
   assign  _net_2193 = (in_do&_net_2);
   assign  _net_2194 = (in_do&_net_2);
   assign  _net_2195 = (in_do&_net_2);
   assign  _net_2196 = (in_do&_net_2);
   assign  _net_2197 = (in_do&_net_2);
   assign  _net_2198 = (in_do&_net_2);
   assign  _net_2199 = (in_do&_net_2);
   assign  _net_2200 = (in_do&_net_2);
   assign  _net_2201 = (in_do&_net_2);
   assign  _net_2202 = (in_do&_net_2);
   assign  _net_2203 = (in_do&_net_2);
   assign  _net_2204 = (in_do&_net_2);
   assign  _net_2205 = (in_do&_net_2);
   assign  _net_2206 = (in_do&_net_2);
   assign  _net_2207 = (in_do&_net_2);
   assign  _net_2208 = (in_do&_net_2);
   assign  _net_2209 = (in_do&_net_2);
   assign  _net_2210 = (in_do&_net_2);
   assign  _net_2211 = (in_do&_net_2);
   assign  _net_2212 = (in_do&_net_2);
   assign  _net_2213 = (in_do&_net_2);
   assign  _net_2214 = (in_do&_net_2);
   assign  _net_2215 = (in_do&_net_2);
   assign  _net_2216 = (in_do&_net_2);
   assign  _net_2217 = (in_do&_net_2);
   assign  _net_2218 = (in_do&_net_2);
   assign  _net_2219 = (in_do&_net_2);
   assign  _net_2220 = (in_do&_net_2);
   assign  _net_2221 = (in_do&_net_2);
   assign  _net_2222 = (in_do&_net_2);
   assign  _net_2223 = (in_do&_net_2);
   assign  _net_2224 = (in_do&_net_2);
   assign  _net_2225 = (in_do&_net_2);
   assign  _net_2226 = (in_do&_net_2);
   assign  _net_2227 = (in_do&_net_2);
   assign  _net_2228 = (in_do&_net_2);
   assign  _net_2229 = (in_do&_net_2);
   assign  _net_2230 = (in_do&_net_2);
   assign  _net_2231 = (in_do&_net_2);
   assign  _net_2232 = (in_do&_net_2);
   assign  _net_2233 = (in_do&_net_2);
   assign  _net_2234 = (in_do&_net_2);
   assign  _net_2235 = (in_do&_net_2);
   assign  _net_2236 = (in_do&_net_2);
   assign  _net_2237 = (in_do&_net_2);
   assign  _net_2238 = (in_do&_net_2);
   assign  _net_2239 = (in_do&_net_2);
   assign  _net_2240 = (in_do&_net_2);
   assign  _net_2241 = (in_do&_net_2);
   assign  _net_2242 = (in_do&_net_2);
   assign  _net_2243 = (in_do&_net_2);
   assign  _net_2244 = (in_do&_net_2);
   assign  _net_2245 = (in_do&_net_2);
   assign  _net_2246 = (in_do&_net_2);
   assign  _net_2247 = (in_do&_net_2);
   assign  _net_2248 = (in_do&_net_2);
   assign  _net_2249 = (in_do&_net_2);
   assign  _net_2250 = (in_do&_net_2);
   assign  _net_2251 = (in_do&_net_2);
   assign  _net_2252 = (in_do&_net_2);
   assign  _net_2253 = (in_do&_net_2);
   assign  _net_2254 = (in_do&_net_2);
   assign  _net_2255 = (in_do&_net_2);
   assign  _net_2256 = (in_do&_net_2);
   assign  _net_2257 = (in_do&_net_2);
   assign  _net_2258 = (in_do&_net_2);
   assign  _net_2259 = (in_do&_net_2);
   assign  _net_2260 = (in_do&_net_2);
   assign  _net_2261 = (in_do&_net_2);
   assign  _net_2262 = (in_do&_net_2);
   assign  _net_2263 = (in_do&_net_2);
   assign  _net_2264 = (in_do&_net_2);
   assign  _net_2265 = (in_do&_net_2);
   assign  _net_2266 = (in_do&_net_2);
   assign  _net_2267 = (in_do&_net_2);
   assign  _net_2268 = (in_do&_net_2);
   assign  _net_2269 = (in_do&_net_2);
   assign  _net_2270 = (in_do&_net_2);
   assign  _net_2271 = (in_do&_net_2);
   assign  _net_2272 = (in_do&_net_2);
   assign  _net_2273 = (in_do&_net_2);
   assign  _net_2274 = (in_do&_net_2);
   assign  _net_2275 = (in_do&_net_2);
   assign  _net_2276 = (in_do&_net_2);
   assign  _net_2277 = (in_do&_net_2);
   assign  _net_2278 = (in_do&_net_2);
   assign  _net_2279 = (in_do&_net_2);
   assign  _net_2280 = (in_do&_net_2);
   assign  _net_2281 = (in_do&_net_2);
   assign  _net_2282 = (in_do&_net_2);
   assign  _net_2283 = (in_do&_net_2);
   assign  _net_2284 = (in_do&_net_2);
   assign  _net_2285 = (in_do&_net_2);
   assign  _net_2286 = (in_do&_net_2);
   assign  _net_2287 = (in_do&_net_2);
   assign  _net_2288 = (in_do&_net_2);
   assign  _net_2289 = (in_do&_net_2);
   assign  _net_2290 = (in_do&_net_2);
   assign  _net_2291 = (in_do&_net_2);
   assign  _net_2292 = (in_do&_net_2);
   assign  _net_2293 = (in_do&_net_2);
   assign  _net_2294 = (in_do&_net_2);
   assign  _net_2295 = (in_do&_net_2);
   assign  _net_2296 = (in_do&_net_2);
   assign  _net_2297 = (in_do&_net_2);
   assign  _net_2298 = (in_do&_net_2);
   assign  _net_2299 = (in_do&_net_2);
   assign  _net_2300 = (in_do&_net_2);
   assign  _net_2301 = (in_do&_net_2);
   assign  _net_2302 = (in_do&_net_2);
   assign  _net_2303 = (in_do&_net_2);
   assign  _net_2304 = (in_do&_net_2);
   assign  _net_2305 = (in_do&_net_2);
   assign  _net_2306 = (in_do&_net_2);
   assign  _net_2307 = (in_do&_net_2);
   assign  _net_2308 = (in_do&_net_2);
   assign  _net_2309 = (in_do&_net_2);
   assign  _net_2310 = (in_do&_net_2);
   assign  _net_2311 = (in_do&_net_2);
   assign  _net_2312 = (in_do&_net_2);
   assign  _net_2313 = (in_do&_net_2);
   assign  _net_2314 = (in_do&_net_2);
   assign  _net_2315 = (in_do&_net_2);
   assign  _net_2316 = (in_do&_net_2);
   assign  _net_2317 = (in_do&_net_2);
   assign  _net_2318 = (in_do&_net_2);
   assign  _net_2319 = (in_do&_net_2);
   assign  _net_2320 = (in_do&_net_2);
   assign  _net_2321 = (in_do&_net_2);
   assign  _net_2322 = (in_do&_net_2);
   assign  _net_2323 = (in_do&_net_2);
   assign  _net_2324 = (in_do&_net_2);
   assign  _net_2325 = (in_do&_net_2);
   assign  _net_2326 = (in_do&_net_2);
   assign  _net_2327 = (in_do&_net_2);
   assign  _net_2328 = (in_do&_net_2);
   assign  _net_2329 = (in_do&_net_2);
   assign  _net_2330 = (in_do&_net_2);
   assign  _net_2331 = (in_do&_net_2);
   assign  _net_2332 = (in_do&_net_2);
   assign  _net_2333 = (in_do&_net_2);
   assign  _net_2334 = (in_do&_net_2);
   assign  _net_2335 = (in_do&_net_2);
   assign  _net_2336 = (in_do&_net_2);
   assign  _net_2337 = (in_do&_net_2);
   assign  _net_2338 = (in_do&_net_2);
   assign  _net_2339 = (in_do&_net_2);
   assign  _net_2340 = (in_do&_net_2);
   assign  _net_2341 = (in_do&_net_2);
   assign  _net_2342 = (in_do&_net_2);
   assign  _net_2343 = (in_do&_net_2);
   assign  _net_2344 = (in_do&_net_2);
   assign  _net_2345 = (in_do&_net_2);
   assign  _net_2346 = (in_do&_net_2);
   assign  _net_2347 = (in_do&_net_2);
   assign  _net_2348 = (in_do&_net_2);
   assign  _net_2349 = (in_do&_net_2);
   assign  _net_2350 = (in_do&_net_2);
   assign  _net_2351 = (in_do&_net_2);
   assign  _net_2352 = (in_do&_net_2);
   assign  _net_2353 = (in_do&_net_2);
   assign  _net_2354 = (in_do&_net_2);
   assign  _net_2355 = (in_do&_net_2);
   assign  _net_2356 = (in_do&_net_2);
   assign  _net_2357 = (in_do&_net_2);
   assign  _net_2358 = (in_do&_net_2);
   assign  _net_2359 = (in_do&_net_2);
   assign  _net_2360 = (in_do&_net_2);
   assign  _net_2361 = (in_do&_net_2);
   assign  _net_2362 = (in_do&_net_2);
   assign  _net_2363 = (in_do&_net_2);
   assign  _net_2364 = (in_do&_net_2);
   assign  _net_2365 = (in_do&_net_2);
   assign  _net_2366 = (in_do&_net_2);
   assign  _net_2367 = (in_do&_net_2);
   assign  _net_2368 = (in_do&_net_2);
   assign  _net_2369 = (in_do&_net_2);
   assign  _net_2370 = (in_do&_net_2);
   assign  _net_2371 = (in_do&_net_2);
   assign  _net_2372 = (in_do&_net_2);
   assign  _net_2373 = (in_do&_net_2);
   assign  _net_2374 = (in_do&_net_2);
   assign  _net_2375 = (in_do&_net_2);
   assign  _net_2376 = (in_do&_net_2);
   assign  _net_2377 = (in_do&_net_2);
   assign  _net_2378 = (in_do&_net_2);
   assign  _net_2379 = (in_do&_net_2);
   assign  _net_2380 = (in_do&_net_2);
   assign  _net_2381 = (in_do&_net_2);
   assign  _net_2382 = (in_do&_net_2);
   assign  _net_2383 = (in_do&_net_2);
   assign  _net_2384 = (in_do&_net_2);
   assign  _net_2385 = (in_do&_net_2);
   assign  _net_2386 = (in_do&_net_2);
   assign  _net_2387 = (in_do&_net_2);
   assign  _net_2388 = (in_do&_net_2);
   assign  _net_2389 = (in_do&_net_2);
   assign  _net_2390 = (in_do&_net_2);
   assign  _net_2391 = (in_do&_net_2);
   assign  _net_2392 = (in_do&_net_2);
   assign  _net_2393 = (in_do&_net_2);
   assign  _net_2394 = (in_do&_net_2);
   assign  _net_2395 = (in_do&_net_2);
   assign  _net_2396 = (in_do&_net_2);
   assign  _net_2397 = (in_do&_net_2);
   assign  _net_2398 = (in_do&_net_2);
   assign  _net_2399 = (in_do&_net_2);
   assign  _net_2400 = (in_do&_net_2);
   assign  _net_2401 = (in_do&_net_2);
   assign  _net_2402 = (in_do&_net_2);
   assign  _net_2403 = (in_do&_net_2);
   assign  _net_2404 = (in_do&_net_2);
   assign  _net_2405 = (in_do&_net_2);
   assign  _net_2406 = (in_do&_net_2);
   assign  _net_2407 = (in_do&_net_2);
   assign  _net_2408 = (in_do&_net_2);
   assign  _net_2409 = (in_do&_net_2);
   assign  _net_2410 = (in_do&_net_2);
   assign  _net_2411 = (in_do&_net_2);
   assign  _net_2412 = (in_do&_net_2);
   assign  _net_2413 = (in_do&_net_2);
   assign  _net_2414 = (in_do&_net_2);
   assign  _net_2415 = (in_do&_net_2);
   assign  _net_2416 = (in_do&_net_2);
   assign  _net_2417 = (in_do&_net_2);
   assign  _net_2418 = (in_do&_net_2);
   assign  _net_2419 = (in_do&_net_2);
   assign  _net_2420 = (in_do&_net_2);
   assign  _net_2421 = (in_do&_net_2);
   assign  _net_2422 = (in_do&_net_2);
   assign  _net_2423 = (in_do&_net_2);
   assign  _net_2424 = (in_do&_net_2);
   assign  _net_2425 = (in_do&_net_2);
   assign  _net_2426 = (in_do&_net_2);
   assign  _net_2427 = (in_do&_net_2);
   assign  _net_2428 = (in_do&_net_2);
   assign  _net_2429 = (in_do&_net_2);
   assign  _net_2430 = (in_do&_net_2);
   assign  _net_2431 = (in_do&_net_2);
   assign  _net_2432 = (in_do&_net_2);
   assign  _net_2433 = (in_do&_net_2);
   assign  _net_2434 = (in_do&_net_2);
   assign  _net_2435 = (in_do&_net_2);
   assign  _net_2436 = (in_do&_net_2);
   assign  _net_2437 = (in_do&_net_2);
   assign  _net_2438 = (in_do&_net_2);
   assign  _net_2439 = (in_do&_net_2);
   assign  _net_2440 = (in_do&_net_2);
   assign  _net_2441 = (in_do&_net_2);
   assign  _net_2442 = (in_do&_net_2);
   assign  _net_2443 = (in_do&_net_2);
   assign  _net_2444 = (in_do&_net_2);
   assign  _net_2445 = (in_do&_net_2);
   assign  _net_2446 = (in_do&_net_2);
   assign  _net_2447 = (in_do&_net_2);
   assign  _net_2448 = (in_do&_net_2);
   assign  _net_2449 = (in_do&_net_2);
   assign  _net_2450 = (in_do&_net_2);
   assign  _net_2451 = (in_do&_net_2);
   assign  _net_2452 = (in_do&_net_2);
   assign  _net_2453 = (in_do&_net_2);
   assign  _net_2454 = (in_do&_net_2);
   assign  _net_2455 = (in_do&_net_2);
   assign  _net_2456 = (in_do&_net_2);
   assign  _net_2457 = (in_do&_net_2);
   assign  _net_2458 = (in_do&_net_2);
   assign  _net_2459 = (in_do&_net_2);
   assign  _net_2460 = (in_do&_net_2);
   assign  _net_2461 = (in_do&_net_2);
   assign  _net_2462 = (in_do&_net_2);
   assign  _net_2463 = (in_do&_net_2);
   assign  _net_2464 = (in_do&_net_2);
   assign  _net_2465 = (in_do&_net_2);
   assign  _net_2466 = (in_do&_net_2);
   assign  _net_2467 = (in_do&_net_2);
   assign  _net_2468 = (in_do&_net_2);
   assign  _net_2469 = (in_do&_net_2);
   assign  _net_2470 = (in_do&_net_2);
   assign  _net_2471 = (in_do&_net_2);
   assign  _net_2472 = (in_do&_net_2);
   assign  _net_2473 = (in_do&_net_2);
   assign  _net_2474 = (in_do&_net_2);
   assign  _net_2475 = (in_do&_net_2);
   assign  _net_2476 = (in_do&_net_2);
   assign  _net_2477 = (in_do&_net_2);
   assign  _net_2478 = (in_do&_net_2);
   assign  _net_2479 = (in_do&_net_2);
   assign  _net_2480 = (in_do&_net_2);
   assign  _net_2481 = (in_do&_net_2);
   assign  _net_2482 = (in_do&_net_2);
   assign  _net_2483 = (in_do&_net_2);
   assign  _net_2484 = (in_do&_net_2);
   assign  _net_2485 = (in_do&_net_2);
   assign  _net_2486 = (in_do&_net_2);
   assign  _net_2487 = (in_do&_net_2);
   assign  _net_2488 = (in_do&_net_2);
   assign  _net_2489 = (in_do&_net_2);
   assign  _net_2490 = (in_do&_net_2);
   assign  _net_2491 = (in_do&_net_2);
   assign  _net_2492 = (in_do&_net_2);
   assign  _net_2493 = (in_do&_net_2);
   assign  _net_2494 = (in_do&_net_2);
   assign  _net_2495 = (in_do&_net_2);
   assign  _net_2496 = (in_do&_net_2);
   assign  _net_2497 = (in_do&_net_2);
   assign  _net_2498 = (in_do&_net_2);
   assign  _net_2499 = (in_do&_net_2);
   assign  _net_2500 = (in_do&_net_2);
   assign  _net_2501 = (in_do&_net_2);
   assign  _net_2502 = (in_do&_net_2);
   assign  _net_2503 = (in_do&_net_2);
   assign  _net_2504 = (in_do&_net_2);
   assign  _net_2505 = (in_do&_net_2);
   assign  _net_2506 = (in_do&_net_2);
   assign  _net_2507 = (in_do&_net_2);
   assign  _net_2508 = (in_do&_net_2);
   assign  _net_2509 = (in_do&_net_2);
   assign  _net_2510 = (in_do&_net_2);
   assign  _net_2511 = (in_do&_net_2);
   assign  _net_2512 = (in_do&_net_2);
   assign  _net_2513 = (in_do&_net_2);
   assign  _net_2514 = (in_do&_net_2);
   assign  _net_2515 = (in_do&_net_2);
   assign  _net_2516 = (in_do&_net_2);
   assign  _net_2517 = (in_do&_net_2);
   assign  _net_2518 = (in_do&_net_2);
   assign  _net_2519 = (in_do&_net_2);
   assign  _net_2520 = (in_do&_net_2);
   assign  _net_2521 = (in_do&_net_2);
   assign  _net_2522 = (in_do&_net_2);
   assign  _net_2523 = (in_do&_net_2);
   assign  _net_2524 = (in_do&_net_2);
   assign  _net_2525 = (in_do&_net_2);
   assign  _net_2526 = (in_do&_net_2);
   assign  _net_2527 = (in_do&_net_2);
   assign  _net_2528 = (in_do&_net_2);
   assign  _net_2529 = (in_do&_net_2);
   assign  _net_2530 = (in_do&_net_2);
   assign  _net_2531 = (in_do&_net_2);
   assign  _net_2532 = (in_do&_net_2);
   assign  _net_2533 = (in_do&_net_2);
   assign  _net_2534 = (in_do&_net_2);
   assign  _net_2535 = (in_do&_net_2);
   assign  _net_2536 = (in_do&_net_2);
   assign  _net_2537 = (in_do&_net_2);
   assign  _net_2538 = (in_do&_net_2);
   assign  _net_2539 = (in_do&_net_2);
   assign  _net_2540 = (in_do&_net_2);
   assign  _net_2541 = (in_do&_net_2);
   assign  _net_2542 = (in_do&_net_2);
   assign  _net_2543 = (in_do&_net_2);
   assign  _net_2544 = (in_do&_net_2);
   assign  _net_2545 = (in_do&_net_2);
   assign  _net_2546 = (in_do&_net_2);
   assign  _net_2547 = (in_do&_net_2);
   assign  _net_2548 = (in_do&_net_2);
   assign  _net_2549 = (in_do&_net_2);
   assign  _net_2550 = (in_do&_net_2);
   assign  _net_2551 = (in_do&_net_2);
   assign  _net_2552 = (in_do&_net_2);
   assign  _net_2553 = (in_do&_net_2);
   assign  _net_2554 = (in_do&_net_2);
   assign  _net_2555 = (in_do&_net_2);
   assign  _net_2556 = (in_do&_net_2);
   assign  _net_2557 = (in_do&_net_2);
   assign  _net_2558 = (in_do&_net_2);
   assign  _net_2559 = (in_do&_net_2);
   assign  _net_2560 = (in_do&_net_2);
   assign  _net_2561 = (in_do&_net_2);
   assign  _net_2562 = (in_do&_net_2);
   assign  _net_2563 = (in_do&_net_2);
   assign  _net_2564 = (in_do&_net_2);
   assign  _net_2565 = (in_do&_net_2);
   assign  _net_2566 = (in_do&_net_2);
   assign  _net_2567 = (in_do&_net_2);
   assign  _net_2568 = (in_do&_net_2);
   assign  _net_2569 = (in_do&_net_2);
   assign  _net_2570 = (in_do&_net_2);
   assign  _net_2571 = (in_do&_net_2);
   assign  _net_2572 = (in_do&_net_2);
   assign  _net_2573 = (in_do&_net_2);
   assign  _net_2574 = (in_do&_net_2);
   assign  _net_2575 = (in_do&_net_2);
   assign  _net_2576 = (in_do&_net_2);
   assign  _net_2577 = (in_do&_net_2);
   assign  _net_2578 = (in_do&_net_2);
   assign  _net_2579 = (in_do&_net_2);
   assign  _net_2580 = (in_do&_net_2);
   assign  _net_2581 = (in_do&_net_2);
   assign  _net_2582 = (in_do&_net_2);
   assign  _net_2583 = (in_do&_net_2);
   assign  _net_2584 = (in_do&_net_2);
   assign  _net_2585 = (in_do&_net_2);
   assign  _net_2586 = (in_do&_net_2);
   assign  _net_2587 = (in_do&_net_2);
   assign  _net_2588 = (in_do&_net_2);
   assign  _net_2589 = (in_do&_net_2);
   assign  _net_2590 = (in_do&_net_2);
   assign  _net_2591 = (in_do&_net_2);
   assign  _net_2592 = (in_do&_net_2);
   assign  _net_2593 = (in_do&_net_2);
   assign  _net_2594 = (in_do&_net_2);
   assign  _net_2595 = (in_do&_net_2);
   assign  _net_2596 = (in_do&_net_2);
   assign  _net_2597 = (in_do&_net_2);
   assign  _net_2598 = (in_do&_net_2);
   assign  _net_2599 = (in_do&_net_2);
   assign  _net_2600 = (in_do&_net_2);
   assign  _net_2601 = (in_do&_net_2);
   assign  _net_2602 = (in_do&_net_2);
   assign  _net_2603 = (in_do&_net_2);
   assign  _net_2604 = (in_do&_net_2);
   assign  _net_2605 = (in_do&_net_2);
   assign  _net_2606 = (in_do&_net_2);
   assign  _net_2607 = (in_do&_net_2);
   assign  _net_2608 = (in_do&_net_2);
   assign  _net_2609 = (in_do&_net_2);
   assign  _net_2610 = (in_do&_net_2);
   assign  _net_2611 = (in_do&_net_2);
   assign  _net_2612 = (in_do&_net_2);
   assign  _net_2613 = (in_do&_net_2);
   assign  _net_2614 = (in_do&_net_2);
   assign  _net_2615 = (in_do&_net_2);
   assign  _net_2616 = (in_do&_net_2);
   assign  _net_2617 = (in_do&_net_2);
   assign  _net_2618 = (in_do&_net_2);
   assign  _net_2619 = (in_do&_net_2);
   assign  _net_2620 = (in_do&_net_2);
   assign  _net_2621 = (in_do&_net_2);
   assign  _net_2622 = (in_do&_net_2);
   assign  _net_2623 = (in_do&_net_2);
   assign  _net_2624 = (in_do&_net_2);
   assign  _net_2625 = (in_do&_net_2);
   assign  _net_2626 = (in_do&_net_2);
   assign  _net_2627 = (in_do&_net_2);
   assign  _net_2628 = (in_do&_net_2);
   assign  _net_2629 = (in_do&_net_2);
   assign  _net_2630 = (in_do&_net_2);
   assign  _net_2631 = (in_do&_net_2);
   assign  _net_2632 = (in_do&_net_2);
   assign  _net_2633 = (in_do&_net_2);
   assign  _net_2634 = (in_do&_net_2);
   assign  _net_2635 = (in_do&_net_2);
   assign  _net_2636 = (in_do&_net_2);
   assign  _net_2637 = (in_do&_net_2);
   assign  _net_2638 = (in_do&_net_2);
   assign  _net_2639 = (in_do&_net_2);
   assign  _net_2640 = (in_do&_net_2);
   assign  _net_2641 = (in_do&_net_2);
   assign  _net_2642 = (in_do&_net_2);
   assign  _net_2643 = (in_do&_net_2);
   assign  _net_2644 = (in_do&_net_2);
   assign  _net_2645 = (in_do&_net_2);
   assign  _net_2646 = (in_do&_net_2);
   assign  _net_2647 = (in_do&_net_2);
   assign  _net_2648 = (in_do&_net_2);
   assign  _net_2649 = (in_do&_net_2);
   assign  _net_2650 = (in_do&_net_2);
   assign  _net_2651 = (in_do&_net_2);
   assign  _net_2652 = (in_do&_net_2);
   assign  _net_2653 = (in_do&_net_2);
   assign  _net_2654 = (in_do&_net_2);
   assign  _net_2655 = (in_do&_net_2);
   assign  _net_2656 = (in_do&_net_2);
   assign  _net_2657 = (in_do&_net_2);
   assign  _net_2658 = (in_do&_net_2);
   assign  _net_2659 = (in_do&_net_2);
   assign  _net_2660 = (in_do&_net_2);
   assign  _net_2661 = (in_do&_net_2);
   assign  _net_2662 = (in_do&_net_2);
   assign  _net_2663 = (in_do&_net_2);
   assign  _net_2664 = (in_do&_net_2);
   assign  _net_2665 = (in_do&_net_2);
   assign  _net_2666 = (in_do&_net_2);
   assign  _net_2667 = (in_do&_net_2);
   assign  _net_2668 = (in_do&_net_2);
   assign  _net_2669 = (in_do&_net_2);
   assign  _net_2670 = (in_do&_net_2);
   assign  _net_2671 = (in_do&_net_2);
   assign  _net_2672 = (in_do&_net_2);
   assign  _net_2673 = (in_do&_net_2);
   assign  _net_2674 = (in_do&_net_2);
   assign  _net_2675 = (in_do&_net_2);
   assign  _net_2676 = (in_do&_net_2);
   assign  _net_2677 = (in_do&_net_2);
   assign  _net_2678 = (in_do&_net_2);
   assign  _net_2679 = (in_do&_net_2);
   assign  _net_2680 = (in_do&_net_2);
   assign  _net_2681 = (in_do&_net_2);
   assign  _net_2682 = (in_do&_net_2);
   assign  _net_2683 = (in_do&_net_2);
   assign  _net_2684 = (in_do&_net_2);
   assign  _net_2685 = (in_do&_net_2);
   assign  _net_2686 = (in_do&_net_2);
   assign  _net_2687 = (in_do&_net_2);
   assign  _net_2688 = (in_do&_net_2);
   assign  _net_2689 = (in_do&_net_2);
   assign  _net_2690 = (in_do&_net_2);
   assign  _net_2691 = (in_do&_net_2);
   assign  _net_2692 = (in_do&_net_2);
   assign  _net_2693 = (in_do&_net_2);
   assign  _net_2694 = (in_do&_net_2);
   assign  _net_2695 = (in_do&_net_2);
   assign  _net_2696 = (in_do&_net_2);
   assign  _net_2697 = (in_do&_net_2);
   assign  _net_2698 = (in_do&_net_2);
   assign  _net_2699 = (in_do&_net_2);
   assign  _net_2700 = (in_do&_net_2);
   assign  _net_2701 = (in_do&_net_2);
   assign  _net_2702 = (in_do&_net_2);
   assign  _net_2703 = (in_do&_net_2);
   assign  _net_2704 = (in_do&_net_2);
   assign  _net_2705 = (in_do&_net_2);
   assign  _net_2706 = (in_do&_net_2);
   assign  _net_2707 = (in_do&_net_2);
   assign  _net_2708 = (in_do&_net_2);
   assign  _net_2709 = (in_do&_net_2);
   assign  _net_2710 = (in_do&_net_2);
   assign  _net_2711 = (in_do&_net_2);
   assign  _net_2712 = (in_do&_net_2);
   assign  _net_2713 = (in_do&_net_2);
   assign  _net_2714 = (in_do&_net_2);
   assign  _net_2715 = (in_do&_net_2);
   assign  _net_2716 = (in_do&_net_2);
   assign  _net_2717 = (in_do&_net_2);
   assign  _net_2718 = (in_do&_net_2);
   assign  _net_2719 = (in_do&_net_2);
   assign  _net_2720 = (in_do&_net_2);
   assign  _net_2721 = (in_do&_net_2);
   assign  _net_2722 = (in_do&_net_2);
   assign  _net_2723 = (in_do&_net_2);
   assign  _net_2724 = (in_do&_net_2);
   assign  _net_2725 = (in_do&_net_2);
   assign  _net_2726 = (in_do&_net_2);
   assign  _net_2727 = (in_do&_net_2);
   assign  _net_2728 = (in_do&_net_2);
   assign  _net_2729 = (in_do&_net_2);
   assign  _net_2730 = (in_do&_net_2);
   assign  _net_2731 = (in_do&_net_2);
   assign  _net_2732 = (in_do&_net_2);
   assign  _net_2733 = (in_do&_net_2);
   assign  _net_2734 = (in_do&_net_2);
   assign  _net_2735 = (in_do&_net_2);
   assign  _net_2736 = (in_do&_net_2);
   assign  _net_2737 = (in_do&_net_2);
   assign  _net_2738 = (in_do&_net_2);
   assign  _net_2739 = (in_do&_net_2);
   assign  _net_2740 = (in_do&_net_2);
   assign  _net_2741 = (in_do&_net_2);
   assign  _net_2742 = (in_do&_net_2);
   assign  _net_2743 = (in_do&_net_2);
   assign  _net_2744 = (in_do&_net_2);
   assign  _net_2745 = (in_do&_net_2);
   assign  _net_2746 = (in_do&_net_2);
   assign  _net_2747 = (in_do&_net_2);
   assign  _net_2748 = (in_do&_net_2);
   assign  _net_2749 = (in_do&_net_2);
   assign  _net_2750 = (in_do&_net_2);
   assign  _net_2751 = (in_do&_net_2);
   assign  _net_2752 = (in_do&_net_2);
   assign  _net_2753 = (in_do&_net_2);
   assign  _net_2754 = (in_do&_net_2);
   assign  _net_2755 = (in_do&_net_2);
   assign  _net_2756 = (in_do&_net_2);
   assign  _net_2757 = (in_do&_net_2);
   assign  _net_2758 = (in_do&_net_2);
   assign  _net_2759 = (in_do&_net_2);
   assign  _net_2760 = (in_do&_net_2);
   assign  _net_2761 = (in_do&_net_2);
   assign  _net_2762 = (in_do&_net_2);
   assign  _net_2763 = (in_do&_net_2);
   assign  _net_2764 = (in_do&_net_2);
   assign  _net_2765 = (in_do&_net_2);
   assign  _net_2766 = (in_do&_net_2);
   assign  _net_2767 = (in_do&_net_2);
   assign  _net_2768 = (in_do&_net_2);
   assign  _net_2769 = (in_do&_net_2);
   assign  _net_2770 = (in_do&_net_2);
   assign  _net_2771 = (in_do&_net_2);
   assign  _net_2772 = (in_do&_net_2);
   assign  _net_2773 = (in_do&_net_2);
   assign  _net_2774 = (in_do&_net_2);
   assign  _net_2775 = (in_do&_net_2);
   assign  _net_2776 = (in_do&_net_2);
   assign  _net_2777 = (in_do&_net_2);
   assign  _net_2778 = (in_do&_net_2);
   assign  _net_2779 = (in_do&_net_2);
   assign  _net_2780 = (in_do&_net_2);
   assign  _net_2781 = (in_do&_net_2);
   assign  _net_2782 = (in_do&_net_2);
   assign  _net_2783 = (in_do&_net_2);
   assign  _net_2784 = (in_do&_net_2);
   assign  _net_2785 = (in_do&_net_2);
   assign  _net_2786 = (in_do&_net_2);
   assign  _net_2787 = (in_do&_net_2);
   assign  _net_2788 = (in_do&_net_2);
   assign  _net_2789 = (in_do&_net_2);
   assign  _net_2790 = (in_do&_net_2);
   assign  _net_2791 = (in_do&_net_2);
   assign  _net_2792 = (in_do&_net_2);
   assign  _net_2793 = (in_do&_net_2);
   assign  _net_2794 = (in_do&_net_2);
   assign  _net_2795 = (in_do&_net_2);
   assign  _net_2796 = (in_do&_net_2);
   assign  _net_2797 = (in_do&_net_2);
   assign  _net_2798 = (in_do&_net_2);
   assign  _net_2799 = (in_do&_net_2);
   assign  _net_2800 = (in_do&_net_2);
   assign  _net_2801 = (in_do&_net_2);
   assign  _net_2802 = (in_do&_net_2);
   assign  _net_2803 = (in_do&_net_2);
   assign  _net_2804 = (in_do&_net_2);
   assign  _net_2805 = (in_do&_net_2);
   assign  _net_2806 = (in_do&_net_2);
   assign  _net_2807 = (in_do&_net_2);
   assign  _net_2808 = (in_do&_net_2);
   assign  _net_2809 = (in_do&_net_2);
   assign  _net_2810 = (in_do&_net_2);
   assign  _net_2811 = (in_do&_net_2);
   assign  _net_2812 = (in_do&_net_2);
   assign  _net_2813 = (in_do&_net_2);
   assign  _net_2814 = (in_do&_net_2);
   assign  _net_2815 = (in_do&_net_2);
   assign  _net_2816 = (in_do&_net_2);
   assign  _net_2817 = (in_do&_net_2);
   assign  _net_2818 = (in_do&_net_2);
   assign  _net_2819 = (in_do&_net_2);
   assign  _net_2820 = (in_do&_net_2);
   assign  _net_2821 = (in_do&_net_2);
   assign  _net_2822 = (in_do&_net_2);
   assign  _net_2823 = (in_do&_net_2);
   assign  _net_2824 = (in_do&_net_2);
   assign  _net_2825 = (in_do&_net_2);
   assign  _net_2826 = (in_do&_net_2);
   assign  _net_2827 = (in_do&_net_2);
   assign  _net_2828 = (in_do&_net_2);
   assign  _net_2829 = (in_do&_net_2);
   assign  _net_2830 = (in_do&_net_2);
   assign  _net_2831 = (in_do&_net_2);
   assign  _net_2832 = (in_do&_net_2);
   assign  _net_2833 = (in_do&_net_2);
   assign  _net_2834 = (in_do&_net_2);
   assign  _net_2835 = (in_do&_net_2);
   assign  _net_2836 = (in_do&_net_2);
   assign  _net_2837 = (in_do&_net_2);
   assign  _net_2838 = (in_do&_net_2);
   assign  _net_2839 = (in_do&_net_2);
   assign  _net_2840 = (in_do&_net_2);
   assign  _net_2841 = (in_do&_net_2);
   assign  _net_2842 = (in_do&_net_2);
   assign  _net_2843 = (in_do&_net_2);
   assign  _net_2844 = (in_do&_net_2);
   assign  _net_2845 = (in_do&_net_2);
   assign  _net_2846 = (in_do&_net_2);
   assign  _net_2847 = (in_do&_net_2);
   assign  _net_2848 = (in_do&_net_2);
   assign  _net_2849 = (in_do&_net_2);
   assign  _net_2850 = (in_do&_net_2);
   assign  _net_2851 = (in_do&_net_2);
   assign  _net_2852 = (in_do&_net_2);
   assign  _net_2853 = (in_do&_net_2);
   assign  _net_2854 = (in_do&_net_2);
   assign  _net_2855 = (in_do&_net_2);
   assign  _net_2856 = (in_do&_net_2);
   assign  _net_2857 = (in_do&_net_2);
   assign  _net_2858 = (in_do&_net_2);
   assign  _net_2859 = (in_do&_net_2);
   assign  _net_2860 = (in_do&_net_2);
   assign  _net_2861 = (in_do&_net_2);
   assign  _net_2862 = (in_do&_net_2);
   assign  _net_2863 = (in_do&_net_2);
   assign  _net_2864 = (in_do&_net_2);
   assign  _net_2865 = (in_do&_net_2);
   assign  _net_2866 = (in_do&_net_2);
   assign  _net_2867 = (in_do&_net_2);
   assign  _net_2868 = (in_do&_net_2);
   assign  _net_2869 = (in_do&_net_2);
   assign  _net_2870 = (in_do&_net_2);
   assign  _net_2871 = (in_do&_net_2);
   assign  _net_2872 = (in_do&_net_2);
   assign  _net_2873 = (in_do&_net_2);
   assign  _net_2874 = (in_do&_net_2);
   assign  _net_2875 = (in_do&_net_2);
   assign  _net_2876 = (in_do&_net_2);
   assign  _net_2877 = (in_do&_net_2);
   assign  _net_2878 = (in_do&_net_2);
   assign  _net_2879 = (in_do&_net_2);
   assign  _net_2880 = (in_do&_net_2);
   assign  _net_2881 = (in_do&_net_2);
   assign  _net_2882 = (in_do&_net_2);
   assign  _net_2883 = (in_do&_net_2);
   assign  _net_2884 = (in_do&_net_2);
   assign  _net_2885 = (in_do&_net_2);
   assign  _net_2886 = (in_do&_net_2);
   assign  _net_2887 = (in_do&_net_2);
   assign  _net_2888 = (in_do&_net_2);
   assign  _net_2889 = (in_do&_net_2);
   assign  _net_2890 = (in_do&_net_2);
   assign  _net_2891 = (in_do&_net_2);
   assign  _net_2892 = (in_do&_net_2);
   assign  _net_2893 = (in_do&_net_2);
   assign  _net_2894 = (in_do&_net_2);
   assign  _net_2895 = (in_do&_net_2);
   assign  _net_2896 = (in_do&_net_2);
   assign  _net_2897 = (in_do&_net_2);
   assign  _net_2898 = (in_do&_net_2);
   assign  _net_2899 = (in_do&_net_2);
   assign  _net_2900 = (in_do&_net_2);
   assign  _net_2901 = (in_do&_net_2);
   assign  _net_2902 = (in_do&_net_2);
   assign  _net_2903 = (in_do&_net_2);
   assign  _net_2904 = (in_do&_net_2);
   assign  _net_2905 = (in_do&_net_2);
   assign  _net_2906 = (in_do&_net_2);
   assign  _net_2907 = (in_do&_net_2);
   assign  _net_2908 = (in_do&_net_2);
   assign  _net_2909 = (in_do&_net_2);
   assign  _net_2910 = (in_do&_net_2);
   assign  _net_2911 = (in_do&_net_2);
   assign  _net_2912 = (in_do&_net_2);
   assign  _net_2913 = (in_do&_net_2);
   assign  _net_2914 = (in_do&_net_2);
   assign  _net_2915 = (in_do&_net_2);
   assign  _net_2916 = (in_do&_net_2);
   assign  _net_2917 = (in_do&_net_2);
   assign  _net_2918 = (in_do&_net_2);
   assign  _net_2919 = (in_do&_net_2);
   assign  _net_2920 = (in_do&_net_2);
   assign  _net_2921 = (in_do&_net_2);
   assign  _net_2922 = (in_do&_net_2);
   assign  _net_2923 = (in_do&_net_2);
   assign  _net_2924 = (in_do&_net_2);
   assign  _net_2925 = (in_do&_net_2);
   assign  _net_2926 = (in_do&_net_2);
   assign  _net_2927 = (in_do&_net_2);
   assign  _net_2928 = (in_do&_net_2);
   assign  _net_2929 = (in_do&_net_2);
   assign  _net_2930 = (in_do&_net_2);
   assign  _net_2931 = (in_do&_net_2);
   assign  _net_2932 = (in_do&_net_2);
   assign  _net_2933 = (in_do&_net_2);
   assign  _net_2934 = (in_do&_net_2);
   assign  _net_2935 = (in_do&_net_2);
   assign  _net_2936 = (in_do&_net_2);
   assign  _net_2937 = (in_do&_net_2);
   assign  _net_2938 = (in_do&_net_2);
   assign  _net_2939 = (in_do&_net_2);
   assign  _net_2940 = (in_do&_net_2);
   assign  _net_2941 = (in_do&_net_2);
   assign  _net_2942 = (in_do&_net_2);
   assign  _net_2943 = (in_do&_net_2);
   assign  _net_2944 = (in_do&_net_2);
   assign  _net_2945 = (in_do&_net_2);
   assign  _net_2946 = (in_do&_net_2);
   assign  _net_2947 = (in_do&_net_2);
   assign  _net_2948 = (in_do&_net_2);
   assign  _net_2949 = (in_do&_net_2);
   assign  _net_2950 = (in_do&_net_2);
   assign  _net_2951 = (in_do&_net_2);
   assign  _net_2952 = (in_do&_net_2);
   assign  _net_2953 = (in_do&_net_2);
   assign  _net_2954 = (in_do&_net_2);
   assign  _net_2955 = (in_do&_net_2);
   assign  _net_2956 = (in_do&_net_2);
   assign  _net_2957 = (in_do&_net_2);
   assign  _net_2958 = (in_do&_net_2);
   assign  _net_2959 = (in_do&_net_2);
   assign  _net_2960 = (in_do&_net_2);
   assign  _net_2961 = (in_do&_net_2);
   assign  _net_2962 = (in_do&_net_2);
   assign  _net_2963 = (in_do&_net_2);
   assign  _net_2964 = (in_do&_net_2);
   assign  _net_2965 = (in_do&_net_2);
   assign  _net_2966 = (in_do&_net_2);
   assign  _net_2967 = (in_do&_net_2);
   assign  _net_2968 = (in_do&_net_2);
   assign  _net_2969 = (in_do&_net_2);
   assign  _net_2970 = (in_do&_net_2);
   assign  _net_2971 = (in_do&_net_2);
   assign  _net_2972 = (in_do&_net_2);
   assign  _net_2973 = (in_do&_net_2);
   assign  _net_2974 = (in_do&_net_2);
   assign  _net_2975 = (in_do&_net_2);
   assign  _net_2976 = (in_do&_net_2);
   assign  _net_2977 = (in_do&_net_2);
   assign  _net_2978 = (in_do&_net_2);
   assign  _net_2979 = (in_do&_net_2);
   assign  _net_2980 = (in_do&_net_2);
   assign  _net_2981 = (in_do&_net_2);
   assign  _net_2982 = (in_do&_net_2);
   assign  _net_2983 = (in_do&_net_2);
   assign  _net_2984 = (in_do&_net_2);
   assign  _net_2985 = (in_do&_net_2);
   assign  _net_2986 = (in_do&_net_2);
   assign  _net_2987 = (in_do&_net_2);
   assign  _net_2988 = (in_do&_net_2);
   assign  _net_2989 = (in_do&_net_2);
   assign  _net_2990 = (in_do&_net_2);
   assign  _net_2991 = (in_do&_net_2);
   assign  _net_2992 = (in_do&_net_2);
   assign  _net_2993 = (in_do&_net_2);
   assign  _net_2994 = (in_do&_net_2);
   assign  _net_2995 = (in_do&_net_2);
   assign  _net_2996 = (in_do&_net_2);
   assign  _net_2997 = (in_do&_net_2);
   assign  _net_2998 = (in_do&_net_2);
   assign  _net_2999 = (in_do&_net_2);
   assign  _net_3000 = (in_do&_net_2);
   assign  _net_3001 = (in_do&_net_2);
   assign  _net_3002 = (in_do&_net_2);
   assign  _net_3003 = (in_do&_net_2);
   assign  _net_3004 = (in_do&_net_2);
   assign  _net_3005 = (in_do&_net_2);
   assign  _net_3006 = (in_do&_net_2);
   assign  _net_3007 = (in_do&_net_2);
   assign  _net_3008 = (in_do&_net_2);
   assign  _net_3009 = (in_do&_net_2);
   assign  _net_3010 = (in_do&_net_2);
   assign  _net_3011 = (in_do&_net_2);
   assign  _net_3012 = (in_do&_net_2);
   assign  _net_3013 = (in_do&_net_2);
   assign  _net_3014 = (in_do&_net_2);
   assign  _net_3015 = (in_do&_net_2);
   assign  _net_3016 = (in_do&_net_2);
   assign  _net_3017 = (in_do&_net_2);
   assign  _net_3018 = (in_do&_net_2);
   assign  _net_3019 = (in_do&_net_2);
   assign  _net_3020 = (in_do&_net_2);
   assign  _net_3021 = (in_do&_net_2);
   assign  _net_3022 = (in_do&_net_2);
   assign  _net_3023 = (in_do&_net_2);
   assign  _net_3024 = (in_do&_net_2);
   assign  _net_3025 = (in_do&_net_2);
   assign  _net_3026 = (in_do&_net_2);
   assign  _net_3027 = (in_do&_net_2);
   assign  _net_3028 = (in_do&_net_2);
   assign  _net_3029 = (in_do&_net_2);
   assign  _net_3030 = (in_do&_net_2);
   assign  _net_3031 = (in_do&_net_2);
   assign  _net_3032 = (in_do&_net_2);
   assign  _net_3033 = (in_do&_net_2);
   assign  _net_3034 = (in_do&_net_2);
   assign  _net_3035 = (in_do&_net_2);
   assign  _net_3036 = (in_do&_net_2);
   assign  _net_3037 = (in_do&_net_2);
   assign  _net_3038 = (in_do&_net_2);
   assign  _net_3039 = (in_do&_net_2);
   assign  _net_3040 = (in_do&_net_2);
   assign  _net_3041 = (in_do&_net_2);
   assign  _net_3042 = (in_do&_net_2);
   assign  _net_3043 = (in_do&_net_2);
   assign  _net_3044 = (in_do&_net_2);
   assign  _net_3045 = (in_do&_net_2);
   assign  _net_3046 = (in_do&_net_2);
   assign  _net_3047 = (in_do&_net_2);
   assign  _net_3048 = (in_do&_net_2);
   assign  _net_3049 = (in_do&_net_2);
   assign  _net_3050 = (in_do&_net_2);
   assign  _net_3051 = (in_do&_net_2);
   assign  _net_3052 = (in_do&_net_2);
   assign  _net_3053 = (in_do&_net_2);
   assign  _net_3054 = (in_do&_net_2);
   assign  _net_3055 = (in_do&_net_2);
   assign  _net_3056 = (in_do&_net_2);
   assign  _net_3057 = (in_do&_net_2);
   assign  _net_3058 = (in_do&_net_2);
   assign  _net_3059 = (in_do&_net_2);
   assign  _net_3060 = (in_do&_net_2);
   assign  _net_3061 = (in_do&_net_2);
   assign  _net_3062 = (in_do&_net_2);
   assign  _net_3063 = (in_do&_net_2);
   assign  _net_3064 = (in_do&_net_2);
   assign  _net_3065 = (in_do&_net_2);
   assign  _net_3066 = (in_do&_net_2);
   assign  _net_3067 = (in_do&_net_2);
   assign  _net_3068 = (in_do&_net_2);
   assign  _net_3069 = (in_do&_net_2);
   assign  _net_3070 = (in_do&_net_2);
   assign  _net_3071 = (in_do&_net_2);
   assign  _net_3072 = (in_do&_net_2);
   assign  _net_3073 = (in_do&_net_2);
   assign  _net_3074 = (in_do&_net_2);
   assign  _net_3075 = (in_do&_net_2);
   assign  _net_3076 = (in_do&_net_2);
   assign  _net_3077 = (in_do&_net_2);
   assign  _net_3078 = (in_do&_net_2);
   assign  _net_3079 = (in_do&_net_2);
   assign  _net_3080 = (in_do&_net_2);
   assign  _net_3081 = (in_do&_net_2);
   assign  _net_3082 = (in_do&_net_2);
   assign  _net_3083 = (in_do&_net_2);
   assign  _net_3084 = (in_do&_net_2);
   assign  _net_3085 = (in_do&_net_2);
   assign  _net_3086 = (in_do&_net_2);
   assign  _net_3087 = (in_do&_net_2);
   assign  _net_3088 = (in_do&_net_2);
   assign  _net_3089 = (in_do&_net_2);
   assign  _net_3090 = (in_do&_net_2);
   assign  _net_3091 = (in_do&_net_2);
   assign  _net_3092 = (in_do&_net_2);
   assign  _net_3093 = (in_do&_net_2);
   assign  _net_3094 = (in_do&_net_2);
   assign  _net_3095 = (in_do&_net_2);
   assign  _net_3096 = (in_do&_net_2);
   assign  _net_3097 = (in_do&_net_2);
   assign  _net_3098 = (in_do&_net_2);
   assign  _net_3099 = (in_do&_net_2);
   assign  _net_3100 = (in_do&_net_2);
   assign  _net_3101 = (in_do&_net_2);
   assign  _net_3102 = (in_do&_net_2);
   assign  _net_3103 = (in_do&_net_2);
   assign  _net_3104 = (in_do&_net_2);
   assign  _net_3105 = (in_do&_net_2);
   assign  _net_3106 = (in_do&_net_2);
   assign  _net_3107 = (in_do&_net_2);
   assign  _net_3108 = (in_do&_net_2);
   assign  _net_3109 = (in_do&_net_2);
   assign  _net_3110 = (in_do&_net_2);
   assign  _net_3111 = (in_do&_net_2);
   assign  _net_3112 = (in_do&_net_2);
   assign  _net_3113 = (in_do&_net_2);
   assign  _net_3114 = (in_do&_net_2);
   assign  _net_3115 = (in_do&_net_2);
   assign  _net_3116 = (in_do&_net_2);
   assign  _net_3117 = (in_do&_net_2);
   assign  _net_3118 = (in_do&_net_2);
   assign  _net_3119 = (in_do&_net_2);
   assign  _net_3120 = (in_do&_net_2);
   assign  _net_3121 = (in_do&_net_2);
   assign  _net_3122 = (in_do&_net_2);
   assign  _net_3123 = (in_do&_net_2);
   assign  _net_3124 = (in_do&_net_2);
   assign  _net_3125 = (in_do&_net_2);
   assign  _net_3126 = (in_do&_net_2);
   assign  _net_3127 = (in_do&_net_2);
   assign  _net_3128 = (in_do&_net_2);
   assign  _net_3129 = (in_do&_net_2);
   assign  _net_3130 = (in_do&_net_2);
   assign  _net_3131 = (in_do&_net_2);
   assign  _net_3132 = (in_do&_net_2);
   assign  _net_3133 = (in_do&_net_2);
   assign  _net_3134 = (in_do&_net_2);
   assign  _net_3135 = (in_do&_net_2);
   assign  _net_3136 = (in_do&_net_2);
   assign  _net_3137 = (in_do&_net_2);
   assign  _net_3138 = (in_do&_net_2);
   assign  _net_3139 = (in_do&_net_2);
   assign  _net_3140 = (in_do&_net_2);
   assign  _net_3141 = (in_do&_net_2);
   assign  _net_3142 = (in_do&_net_2);
   assign  _net_3143 = (in_do&_net_2);
   assign  _net_3144 = (in_do&_net_2);
   assign  _net_3145 = (in_do&_net_2);
   assign  _net_3146 = (in_do&_net_2);
   assign  _net_3147 = (in_do&_net_2);
   assign  _net_3148 = (in_do&_net_2);
   assign  _net_3149 = (in_do&_net_2);
   assign  _net_3150 = (in_do&_net_2);
   assign  _net_3151 = (in_do&_net_2);
   assign  _net_3152 = (in_do&_net_2);
   assign  _net_3153 = (in_do&_net_2);
   assign  _net_3154 = (in_do&_net_2);
   assign  _net_3155 = (in_do&_net_2);
   assign  _net_3156 = (in_do&_net_2);
   assign  _net_3157 = (in_do&_net_2);
   assign  _net_3158 = (in_do&_net_2);
   assign  _net_3159 = (in_do&_net_2);
   assign  _net_3160 = (in_do&_net_2);
   assign  _net_3161 = (in_do&_net_2);
   assign  _net_3162 = (in_do&_net_2);
   assign  _net_3163 = (in_do&_net_2);
   assign  _net_3164 = (in_do&_net_2);
   assign  _net_3165 = (in_do&_net_2);
   assign  _net_3166 = (in_do&_net_2);
   assign  _net_3167 = (in_do&_net_2);
   assign  _net_3168 = (in_do&_net_2);
   assign  _net_3169 = (in_do&_net_2);
   assign  _net_3170 = (in_do&_net_2);
   assign  _net_3171 = (in_do&_net_2);
   assign  _net_3172 = (in_do&_net_2);
   assign  _net_3173 = (in_do&_net_2);
   assign  _net_3174 = (in_do&_net_2);
   assign  _net_3175 = (in_do&_net_2);
   assign  _net_3176 = (in_do&_net_2);
   assign  _net_3177 = (in_do&_net_2);
   assign  _net_3178 = (in_do&_net_2);
   assign  _net_3179 = (in_do&_net_2);
   assign  _net_3180 = (in_do&_net_2);
   assign  _net_3181 = (in_do&_net_2);
   assign  _net_3182 = (in_do&_net_2);
   assign  _net_3183 = (in_do&_net_2);
   assign  _net_3184 = (in_do&_net_2);
   assign  _net_3185 = (in_do&_net_2);
   assign  _net_3186 = (in_do&_net_2);
   assign  _net_3187 = (in_do&_net_2);
   assign  _net_3188 = (in_do&_net_2);
   assign  _net_3189 = (in_do&_net_2);
   assign  _net_3190 = (in_do&_net_2);
   assign  _net_3191 = (in_do&_net_2);
   assign  _net_3192 = (in_do&_net_2);
   assign  _net_3193 = (in_do&_net_2);
   assign  _net_3194 = (in_do&_net_2);
   assign  _net_3195 = (in_do&_net_2);
   assign  _net_3196 = (in_do&_net_2);
   assign  _net_3197 = (in_do&_net_2);
   assign  _net_3198 = (in_do&_net_2);
   assign  _net_3199 = (in_do&_net_2);
   assign  _net_3200 = (in_do&_net_2);
   assign  _net_3201 = (in_do&_net_2);
   assign  _net_3202 = (in_do&_net_2);
   assign  _net_3203 = (in_do&_net_2);
   assign  _net_3204 = (in_do&_net_2);
   assign  _net_3205 = (in_do&_net_2);
   assign  _net_3206 = (in_do&_net_2);
   assign  _net_3207 = (in_do&_net_2);
   assign  _net_3208 = (in_do&_net_2);
   assign  _net_3209 = (in_do&_net_2);
   assign  _net_3210 = (in_do&_net_2);
   assign  _net_3211 = (in_do&_net_2);
   assign  _net_3212 = (in_do&_net_2);
   assign  _net_3213 = (in_do&_net_2);
   assign  _net_3214 = (in_do&_net_2);
   assign  _net_3215 = (in_do&_net_2);
   assign  _net_3216 = (in_do&_net_2);
   assign  _net_3217 = (in_do&_net_2);
   assign  _net_3218 = (in_do&_net_2);
   assign  _net_3219 = (in_do&_net_2);
   assign  _net_3220 = (in_do&_net_2);
   assign  _net_3221 = (in_do&_net_2);
   assign  _net_3222 = (in_do&_net_2);
   assign  _net_3223 = (in_do&_net_2);
   assign  _net_3224 = (in_do&_net_2);
   assign  _net_3225 = (in_do&_net_2);
   assign  _net_3226 = (in_do&_net_2);
   assign  _net_3227 = (in_do&_net_2);
   assign  _net_3228 = (in_do&_net_2);
   assign  _net_3229 = (in_do&_net_2);
   assign  _net_3230 = (in_do&_net_2);
   assign  _net_3231 = (in_do&_net_2);
   assign  _net_3232 = (in_do&_net_2);
   assign  _net_3233 = (in_do&_net_2);
   assign  _net_3234 = (in_do&_net_2);
   assign  _net_3235 = (in_do&_net_2);
   assign  _net_3236 = (in_do&_net_2);
   assign  _net_3237 = (in_do&_net_2);
   assign  _net_3238 = (in_do&_net_2);
   assign  _net_3239 = (in_do&_net_2);
   assign  _net_3240 = (in_do&_net_2);
   assign  _net_3241 = (in_do&_net_2);
   assign  _net_3242 = (in_do&_net_2);
   assign  _net_3243 = (in_do&_net_2);
   assign  _net_3244 = (in_do&_net_2);
   assign  _net_3245 = (in_do&_net_2);
   assign  _net_3246 = (in_do&_net_2);
   assign  _net_3247 = (in_do&_net_2);
   assign  _net_3248 = (in_do&_net_2);
   assign  _net_3249 = (in_do&_net_2);
   assign  _net_3250 = (in_do&_net_2);
   assign  _net_3251 = (in_do&_net_2);
   assign  _net_3252 = (in_do&_net_2);
   assign  _net_3253 = (in_do&_net_2);
   assign  _net_3254 = (in_do&_net_2);
   assign  _net_3255 = (in_do&_net_2);
   assign  _net_3256 = (in_do&_net_2);
   assign  _net_3257 = (in_do&_net_2);
   assign  _net_3258 = (in_do&_net_2);
   assign  _net_3259 = (in_do&_net_2);
   assign  _net_3260 = (in_do&_net_2);
   assign  _net_3261 = (in_do&_net_2);
   assign  _net_3262 = (in_do&_net_2);
   assign  _net_3263 = (in_do&_net_2);
   assign  _net_3264 = (in_do&_net_2);
   assign  _net_3265 = (in_do&_net_2);
   assign  _net_3266 = (in_do&_net_2);
   assign  _net_3267 = (in_do&_net_2);
   assign  _net_3268 = (in_do&_net_2);
   assign  _net_3269 = (in_do&_net_2);
   assign  _net_3270 = (in_do&_net_2);
   assign  _net_3271 = (in_do&_net_2);
   assign  _net_3272 = (in_do&_net_2);
   assign  _net_3273 = (in_do&_net_2);
   assign  _net_3274 = (in_do&_net_2);
   assign  _net_3275 = (in_do&_net_2);
   assign  _net_3276 = (in_do&_net_2);
   assign  _net_3277 = (in_do&_net_2);
   assign  _net_3278 = (in_do&_net_2);
   assign  _net_3279 = (in_do&_net_2);
   assign  _net_3280 = (in_do&_net_2);
   assign  _net_3281 = (in_do&_net_2);
   assign  _net_3282 = (in_do&_net_2);
   assign  _net_3283 = (in_do&_net_2);
   assign  _net_3284 = (in_do&_net_2);
   assign  _net_3285 = (in_do&_net_2);
   assign  _net_3286 = (in_do&_net_2);
   assign  _net_3287 = (in_do&_net_2);
   assign  _net_3288 = (in_do&_net_2);
   assign  _net_3289 = (in_do&_net_2);
   assign  _net_3290 = (in_do&_net_2);
   assign  _net_3291 = (in_do&_net_2);
   assign  _net_3292 = (in_do&_net_2);
   assign  _net_3293 = (in_do&_net_2);
   assign  _net_3294 = (in_do&_net_2);
   assign  _net_3295 = (in_do&_net_2);
   assign  _net_3296 = (in_do&_net_2);
   assign  _net_3297 = (in_do&_net_2);
   assign  _net_3298 = (in_do&_net_2);
   assign  _net_3299 = (in_do&_net_2);
   assign  _net_3300 = (in_do&_net_2);
   assign  _net_3301 = (in_do&_net_2);
   assign  _net_3302 = (in_do&_net_2);
   assign  _net_3303 = (in_do&_net_2);
   assign  _net_3304 = (in_do&_net_2);
   assign  _net_3305 = (in_do&_net_2);
   assign  _net_3306 = (in_do&_net_2);
   assign  _net_3307 = (in_do&_net_2);
   assign  _net_3308 = (in_do&_net_2);
   assign  _net_3309 = (in_do&_net_2);
   assign  _net_3310 = (in_do&_net_2);
   assign  _net_3311 = (in_do&_net_2);
   assign  _net_3312 = (in_do&_net_2);
   assign  _net_3313 = (in_do&_net_2);
   assign  _net_3314 = (in_do&_net_2);
   assign  _net_3315 = (in_do&_net_2);
   assign  _net_3316 = (in_do&_net_2);
   assign  _net_3317 = (in_do&_net_2);
   assign  _net_3318 = (in_do&_net_2);
   assign  _net_3319 = (in_do&_net_2);
   assign  _net_3320 = (in_do&_net_2);
   assign  _net_3321 = (in_do&_net_2);
   assign  _net_3322 = (in_do&_net_2);
   assign  _net_3323 = (in_do&_net_2);
   assign  _net_3324 = (in_do&_net_2);
   assign  _net_3325 = (in_do&_net_2);
   assign  _net_3326 = (in_do&_net_2);
   assign  _net_3327 = (in_do&_net_2);
   assign  _net_3328 = (in_do&_net_2);
   assign  _net_3329 = (in_do&_net_2);
   assign  _net_3330 = (in_do&_net_2);
   assign  _net_3331 = (in_do&_net_2);
   assign  _net_3332 = (in_do&_net_2);
   assign  _net_3333 = (in_do&_net_2);
   assign  _net_3334 = (in_do&_net_2);
   assign  _net_3335 = (in_do&_net_2);
   assign  _net_3336 = (in_do&_net_2);
   assign  _net_3337 = (in_do&_net_2);
   assign  _net_3338 = (in_do&_net_2);
   assign  _net_3339 = (in_do&_net_2);
   assign  _net_3340 = (in_do&_net_2);
   assign  _net_3341 = (in_do&_net_2);
   assign  _net_3342 = (in_do&_net_2);
   assign  _net_3343 = (in_do&_net_2);
   assign  _net_3344 = (in_do&_net_2);
   assign  _net_3345 = (in_do&_net_2);
   assign  _net_3346 = (in_do&_net_2);
   assign  _net_3347 = (in_do&_net_2);
   assign  _net_3348 = (in_do&_net_2);
   assign  _net_3349 = (in_do&_net_2);
   assign  _net_3350 = (in_do&_net_2);
   assign  _net_3351 = (in_do&_net_2);
   assign  _net_3352 = (in_do&_net_2);
   assign  _net_3353 = (in_do&_net_2);
   assign  _net_3354 = (in_do&_net_2);
   assign  _net_3355 = (in_do&_net_2);
   assign  _net_3356 = (in_do&_net_2);
   assign  _net_3357 = (in_do&_net_2);
   assign  _net_3358 = (in_do&_net_2);
   assign  _net_3359 = (in_do&_net_2);
   assign  _net_3360 = (in_do&_net_2);
   assign  _net_3361 = (in_do&_net_2);
   assign  _net_3362 = (in_do&_net_2);
   assign  _net_3363 = (in_do&_net_2);
   assign  _net_3364 = (in_do&_net_2);
   assign  _net_3365 = (in_do&_net_2);
   assign  _net_3366 = (in_do&_net_2);
   assign  _net_3367 = (in_do&_net_2);
   assign  _net_3368 = (in_do&_net_2);
   assign  _net_3369 = (in_do&_net_2);
   assign  _net_3370 = (in_do&_net_2);
   assign  _net_3371 = (in_do&_net_2);
   assign  _net_3372 = (in_do&_net_2);
   assign  _net_3373 = (in_do&_net_2);
   assign  _net_3374 = (in_do&_net_2);
   assign  _net_3375 = (in_do&_net_2);
   assign  _net_3376 = (in_do&_net_2);
   assign  _net_3377 = (in_do&_net_2);
   assign  _net_3378 = (in_do&_net_2);
   assign  _net_3379 = (in_do&_net_2);
   assign  _net_3380 = (in_do&_net_2);
   assign  _net_3381 = (in_do&_net_2);
   assign  _net_3382 = (in_do&_net_2);
   assign  _net_3383 = (in_do&_net_2);
   assign  _net_3384 = (in_do&_net_2);
   assign  _net_3385 = (in_do&_net_2);
   assign  _net_3386 = (in_do&_net_2);
   assign  _net_3387 = (in_do&_net_2);
   assign  _net_3388 = (in_do&_net_2);
   assign  _net_3389 = (in_do&_net_2);
   assign  _net_3390 = (in_do&_net_2);
   assign  _net_3391 = (in_do&_net_2);
   assign  _net_3392 = (in_do&_net_2);
   assign  _net_3393 = (in_do&_net_2);
   assign  _net_3394 = (in_do&_net_2);
   assign  _net_3395 = (in_do&_net_2);
   assign  _net_3396 = (in_do&_net_2);
   assign  _net_3397 = (in_do&_net_2);
   assign  _net_3398 = (in_do&_net_2);
   assign  _net_3399 = (in_do&_net_2);
   assign  _net_3400 = (in_do&_net_2);
   assign  _net_3401 = (in_do&_net_2);
   assign  _net_3402 = (in_do&_net_2);
   assign  _net_3403 = (in_do&_net_2);
   assign  _net_3404 = (in_do&_net_2);
   assign  _net_3405 = (in_do&_net_2);
   assign  _net_3406 = (in_do&_net_2);
   assign  _net_3407 = (in_do&_net_2);
   assign  _net_3408 = (in_do&_net_2);
   assign  _net_3409 = (in_do&_net_2);
   assign  _net_3410 = (in_do&_net_2);
   assign  _net_3411 = (in_do&_net_2);
   assign  _net_3412 = (in_do&_net_2);
   assign  _net_3413 = (in_do&_net_2);
   assign  _net_3414 = (in_do&_net_2);
   assign  _net_3415 = (in_do&_net_2);
   assign  _net_3416 = (in_do&_net_2);
   assign  _net_3417 = (in_do&_net_2);
   assign  _net_3418 = (in_do&_net_2);
   assign  _net_3419 = (in_do&_net_2);
   assign  _net_3420 = (in_do&_net_2);
   assign  _net_3421 = (in_do&_net_2);
   assign  _net_3422 = (in_do&_net_2);
   assign  _net_3423 = (in_do&_net_2);
   assign  _net_3424 = (in_do&_net_2);
   assign  _net_3425 = (in_do&_net_2);
   assign  _net_3426 = (in_do&_net_2);
   assign  _net_3427 = (in_do&_net_2);
   assign  _net_3428 = (in_do&_net_2);
   assign  _net_3429 = (in_do&_net_2);
   assign  _net_3430 = (in_do&_net_2);
   assign  _net_3431 = (in_do&_net_2);
   assign  _net_3432 = (in_do&_net_2);
   assign  _net_3433 = (in_do&_net_2);
   assign  _net_3434 = (in_do&_net_2);
   assign  _net_3435 = (in_do&_net_2);
   assign  _net_3436 = (in_do&_net_2);
   assign  _net_3437 = (in_do&_net_2);
   assign  _net_3438 = (in_do&_net_2);
   assign  _net_3439 = (in_do&_net_2);
   assign  _net_3440 = (in_do&_net_2);
   assign  _net_3441 = (in_do&_net_2);
   assign  _net_3442 = (in_do&_net_2);
   assign  _net_3443 = (in_do&_net_2);
   assign  _net_3444 = (in_do&_net_2);
   assign  _net_3445 = (in_do&_net_2);
   assign  _net_3446 = (in_do&_net_2);
   assign  _net_3447 = (in_do&_net_2);
   assign  _net_3448 = (in_do&_net_2);
   assign  _net_3449 = (in_do&_net_2);
   assign  _net_3450 = (in_do&_net_2);
   assign  _net_3451 = (in_do&_net_2);
   assign  _net_3452 = (in_do&_net_2);
   assign  _net_3453 = (in_do&_net_2);
   assign  _net_3454 = (in_do&_net_2);
   assign  _net_3455 = (in_do&_net_2);
   assign  _net_3456 = (in_do&_net_2);
   assign  _net_3457 = (in_do&_net_2);
   assign  _net_3458 = (in_do&_net_2);
   assign  _net_3459 = (in_do&_net_2);
   assign  _net_3460 = (in_do&_net_2);
   assign  _net_3461 = (in_do&_net_2);
   assign  _net_3462 = (in_do&_net_2);
   assign  _net_3463 = (in_do&_net_2);
   assign  _net_3464 = (in_do&_net_2);
   assign  _net_3465 = (in_do&_net_2);
   assign  _net_3466 = (in_do&_net_2);
   assign  _net_3467 = (in_do&_net_2);
   assign  _net_3468 = (in_do&_net_2);
   assign  _net_3469 = (in_do&_net_2);
   assign  _net_3470 = (in_do&_net_2);
   assign  _net_3471 = (in_do&_net_2);
   assign  _net_3472 = (in_do&_net_2);
   assign  _net_3473 = (in_do&_net_2);
   assign  _net_3474 = (in_do&_net_2);
   assign  _net_3475 = (in_do&_net_2);
   assign  _net_3476 = (in_do&_net_2);
   assign  _net_3477 = (in_do&_net_2);
   assign  _net_3478 = (in_do&_net_2);
   assign  _net_3479 = (in_do&_net_2);
   assign  _net_3480 = (in_do&_net_2);
   assign  _net_3481 = (in_do&_net_2);
   assign  _net_3482 = (in_do&_net_2);
   assign  _net_3483 = (in_do&_net_2);
   assign  _net_3484 = (in_do&_net_2);
   assign  _net_3485 = (in_do&_net_2);
   assign  _net_3486 = (in_do&_net_2);
   assign  _net_3487 = (in_do&_net_2);
   assign  _net_3488 = (in_do&_net_2);
   assign  _net_3489 = (in_do&_net_2);
   assign  _net_3490 = (in_do&_net_2);
   assign  _net_3491 = (in_do&_net_2);
   assign  _net_3492 = (in_do&_net_2);
   assign  _net_3493 = (in_do&_net_2);
   assign  _net_3494 = (in_do&_net_2);
   assign  _net_3495 = (in_do&_net_2);
   assign  _net_3496 = (in_do&_net_2);
   assign  _net_3497 = (in_do&_net_2);
   assign  _net_3498 = (in_do&_net_2);
   assign  _net_3499 = (in_do&_net_2);
   assign  _net_3500 = (in_do&_net_2);
   assign  _net_3501 = (in_do&_net_2);
   assign  _net_3502 = (in_do&_net_2);
   assign  _net_3503 = (in_do&_net_2);
   assign  _net_3504 = (in_do&_net_2);
   assign  _net_3505 = (in_do&_net_2);
   assign  _net_3506 = (in_do&_net_2);
   assign  _net_3507 = (in_do&_net_2);
   assign  _net_3508 = (in_do&_net_2);
   assign  _net_3509 = (in_do&_net_2);
   assign  _net_3510 = (in_do&_net_2);
   assign  _net_3511 = (in_do&_net_2);
   assign  _net_3512 = (in_do&_net_2);
   assign  _net_3513 = (in_do&_net_2);
   assign  _net_3514 = (in_do&_net_2);
   assign  _net_3515 = (in_do&_net_2);
   assign  _net_3516 = (in_do&_net_2);
   assign  _net_3517 = (in_do&_net_2);
   assign  _net_3518 = (in_do&_net_2);
   assign  _net_3519 = (in_do&_net_2);
   assign  _net_3520 = (in_do&_net_2);
   assign  _net_3521 = (in_do&_net_2);
   assign  _net_3522 = (in_do&_net_2);
   assign  _net_3523 = (in_do&_net_2);
   assign  _net_3524 = (in_do&_net_2);
   assign  _net_3525 = (in_do&_net_2);
   assign  _net_3526 = (in_do&_net_2);
   assign  _net_3527 = (in_do&_net_2);
   assign  _net_3528 = (in_do&_net_2);
   assign  _net_3529 = (in_do&_net_2);
   assign  _net_3530 = (in_do&_net_2);
   assign  _net_3531 = (in_do&_net_2);
   assign  _net_3532 = (in_do&_net_2);
   assign  _net_3533 = (in_do&_net_2);
   assign  _net_3534 = (in_do&_net_2);
   assign  _net_3535 = (in_do&_net_2);
   assign  _net_3536 = (in_do&_net_2);
   assign  _net_3537 = (in_do&_net_2);
   assign  _net_3538 = (in_do&_net_2);
   assign  _net_3539 = (in_do&_net_2);
   assign  _net_3540 = (in_do&_net_2);
   assign  _net_3541 = (in_do&_net_2);
   assign  _net_3542 = (in_do&_net_2);
   assign  _net_3543 = (in_do&_net_2);
   assign  _net_3544 = (in_do&_net_2);
   assign  _net_3545 = (in_do&_net_2);
   assign  _net_3546 = (in_do&_net_2);
   assign  _net_3547 = (in_do&_net_2);
   assign  _net_3548 = (in_do&_net_2);
   assign  _net_3549 = (in_do&_net_2);
   assign  _net_3550 = (in_do&_net_2);
   assign  _net_3551 = (in_do&_net_2);
   assign  _net_3552 = (in_do&_net_2);
   assign  _net_3553 = (in_do&_net_2);
   assign  _net_3554 = (in_do&_net_2);
   assign  _net_3555 = (in_do&_net_2);
   assign  _net_3556 = (in_do&_net_2);
   assign  _net_3557 = (in_do&_net_2);
   assign  _net_3558 = (in_do&_net_2);
   assign  _net_3559 = (in_do&_net_2);
   assign  _net_3560 = (in_do&_net_2);
   assign  _net_3561 = (in_do&_net_2);
   assign  _net_3562 = (in_do&_net_2);
   assign  _net_3563 = (in_do&_net_2);
   assign  _net_3564 = (in_do&_net_2);
   assign  _net_3565 = (in_do&_net_2);
   assign  _net_3566 = (in_do&_net_2);
   assign  _net_3567 = (in_do&_net_2);
   assign  _net_3568 = (in_do&_net_2);
   assign  _net_3569 = (in_do&_net_2);
   assign  _net_3570 = (in_do&_net_2);
   assign  _net_3571 = (in_do&_net_2);
   assign  _net_3572 = (in_do&_net_2);
   assign  _net_3573 = (in_do&_net_2);
   assign  _net_3574 = (in_do&_net_2);
   assign  _net_3575 = (in_do&_net_2);
   assign  _net_3576 = (in_do&_net_2);
   assign  _net_3577 = (in_do&_net_2);
   assign  _net_3578 = (in_do&_net_2);
   assign  _net_3579 = (in_do&_net_2);
   assign  _net_3580 = (in_do&_net_2);
   assign  _net_3581 = (in_do&_net_2);
   assign  _net_3582 = (in_do&_net_2);
   assign  _net_3583 = (in_do&_net_2);
   assign  _net_3584 = (in_do&_net_2);
   assign  _net_3585 = (in_do&_net_2);
   assign  _net_3586 = (in_do&_net_2);
   assign  _net_3587 = (in_do&_net_2);
   assign  _net_3588 = (in_do&_net_2);
   assign  _net_3589 = (in_do&_net_2);
   assign  _net_3590 = (in_do&_net_2);
   assign  _net_3591 = (in_do&_net_2);
   assign  _net_3592 = (in_do&_net_2);
   assign  _net_3593 = (in_do&_net_2);
   assign  _net_3594 = (in_do&_net_2);
   assign  _net_3595 = (in_do&_net_2);
   assign  _net_3596 = (in_do&_net_2);
   assign  _net_3597 = (in_do&_net_2);
   assign  _net_3598 = (in_do&_net_2);
   assign  _net_3599 = (in_do&_net_2);
   assign  _net_3600 = (in_do&_net_2);
   assign  _net_3601 = (in_do&_net_2);
   assign  _net_3602 = (in_do&_net_2);
   assign  _net_3603 = (in_do&_net_2);
   assign  _net_3604 = (in_do&_net_2);
   assign  _net_3605 = (in_do&_net_2);
   assign  _net_3606 = (in_do&_net_2);
   assign  _net_3607 = (in_do&_net_2);
   assign  _net_3608 = (in_do&_net_2);
   assign  _net_3609 = (in_do&_net_2);
   assign  _net_3610 = (in_do&_net_2);
   assign  _net_3611 = (in_do&_net_2);
   assign  _net_3612 = (in_do&_net_2);
   assign  _net_3613 = (in_do&_net_2);
   assign  _net_3614 = (in_do&_net_2);
   assign  _net_3615 = (in_do&_net_2);
   assign  _net_3616 = (in_do&_net_2);
   assign  _net_3617 = (in_do&_net_2);
   assign  _net_3618 = (in_do&_net_2);
   assign  _net_3619 = (in_do&_net_2);
   assign  _net_3620 = (in_do&_net_2);
   assign  _net_3621 = (in_do&_net_2);
   assign  _net_3622 = (in_do&_net_2);
   assign  _net_3623 = (in_do&_net_2);
   assign  _net_3624 = (in_do&_net_2);
   assign  _net_3625 = (in_do&_net_2);
   assign  _net_3626 = (in_do&_net_2);
   assign  _net_3627 = (in_do&_net_2);
   assign  _net_3628 = (in_do&_net_2);
   assign  _net_3629 = (in_do&_net_2);
   assign  _net_3630 = (in_do&_net_2);
   assign  _net_3631 = (in_do&_net_2);
   assign  _net_3632 = (in_do&_net_2);
   assign  _net_3633 = (in_do&_net_2);
   assign  _net_3634 = (in_do&_net_2);
   assign  _net_3635 = (in_do&_net_2);
   assign  _net_3636 = (in_do&_net_2);
   assign  _net_3637 = (in_do&_net_2);
   assign  _net_3638 = (in_do&_net_2);
   assign  _net_3639 = (in_do&_net_2);
   assign  _net_3640 = (in_do&_net_2);
   assign  _net_3641 = (in_do&_net_2);
   assign  _net_3642 = (in_do&_net_2);
   assign  _net_3643 = (in_do&_net_2);
   assign  _net_3644 = (in_do&_net_2);
   assign  _net_3645 = (in_do&_net_2);
   assign  _net_3646 = (in_do&_net_2);
   assign  _net_3647 = (in_do&_net_2);
   assign  _net_3648 = (in_do&_net_2);
   assign  _net_3649 = (in_do&_net_2);
   assign  _net_3650 = (in_do&_net_2);
   assign  _net_3651 = (in_do&_net_2);
   assign  _net_3652 = (in_do&_net_2);
   assign  _net_3653 = (in_do&_net_2);
   assign  _net_3654 = (in_do&_net_2);
   assign  _net_3655 = (in_do&_net_2);
   assign  _net_3656 = (in_do&_net_2);
   assign  _net_3657 = (in_do&_net_2);
   assign  _net_3658 = (in_do&_net_2);
   assign  _net_3659 = (in_do&_net_2);
   assign  _net_3660 = (in_do&_net_2);
   assign  _net_3661 = (in_do&_net_2);
   assign  _net_3662 = (in_do&_net_2);
   assign  _net_3663 = (in_do&_net_2);
   assign  _net_3664 = (in_do&_net_2);
   assign  _net_3665 = (in_do&_net_2);
   assign  _net_3666 = (in_do&_net_2);
   assign  _net_3667 = (in_do&_net_2);
   assign  _net_3668 = (in_do&_net_2);
   assign  _net_3669 = (in_do&_net_2);
   assign  _net_3670 = (in_do&_net_2);
   assign  _net_3671 = (in_do&_net_2);
   assign  _net_3672 = (in_do&_net_2);
   assign  _net_3673 = (in_do&_net_2);
   assign  _net_3674 = (in_do&_net_2);
   assign  _net_3675 = (in_do&_net_2);
   assign  _net_3676 = (in_do&_net_2);
   assign  _net_3677 = (in_do&_net_2);
   assign  _net_3678 = (in_do&_net_2);
   assign  _net_3679 = (in_do&_net_2);
   assign  _net_3680 = (in_do&_net_2);
   assign  _net_3681 = (in_do&_net_2);
   assign  _net_3682 = (in_do&_net_2);
   assign  _net_3683 = (in_do&_net_2);
   assign  _net_3684 = (in_do&_net_2);
   assign  _net_3685 = (in_do&_net_2);
   assign  _net_3686 = (in_do&_net_2);
   assign  _net_3687 = (in_do&_net_2);
   assign  _net_3688 = (in_do&_net_2);
   assign  _net_3689 = (in_do&_net_2);
   assign  _net_3690 = (in_do&_net_2);
   assign  _net_3691 = (in_do&_net_2);
   assign  _net_3692 = (in_do&_net_2);
   assign  _net_3693 = (in_do&_net_2);
   assign  _net_3694 = (in_do&_net_2);
   assign  _net_3695 = (in_do&_net_2);
   assign  _net_3696 = (in_do&_net_2);
   assign  _net_3697 = (in_do&_net_2);
   assign  _net_3698 = (in_do&_net_2);
   assign  _net_3699 = (in_do&_net_2);
   assign  _net_3700 = (in_do&_net_2);
   assign  _net_3701 = (in_do&_net_2);
   assign  _net_3702 = (in_do&_net_2);
   assign  _net_3703 = (in_do&_net_2);
   assign  _net_3704 = (in_do&_net_2);
   assign  _net_3705 = (in_do&_net_2);
   assign  _net_3706 = (in_do&_net_2);
   assign  _net_3707 = (in_do&_net_2);
   assign  _net_3708 = (in_do&_net_2);
   assign  _net_3709 = (in_do&_net_2);
   assign  _net_3710 = (in_do&_net_2);
   assign  _net_3711 = (in_do&_net_2);
   assign  _net_3712 = (in_do&_net_2);
   assign  _net_3713 = (in_do&_net_2);
   assign  _net_3714 = (in_do&_net_2);
   assign  _net_3715 = (in_do&_net_2);
   assign  _net_3716 = (in_do&_net_2);
   assign  _net_3717 = (in_do&_net_2);
   assign  _net_3718 = (in_do&_net_2);
   assign  _net_3719 = (in_do&_net_2);
   assign  _net_3720 = (in_do&_net_2);
   assign  _net_3721 = (in_do&_net_2);
   assign  _net_3722 = (in_do&_net_2);
   assign  _net_3723 = (in_do&_net_2);
   assign  _net_3724 = (in_do&_net_2);
   assign  _net_3725 = (in_do&_net_2);
   assign  _net_3726 = (in_do&_net_2);
   assign  _net_3727 = (in_do&_net_2);
   assign  _net_3728 = (in_do&_net_2);
   assign  _net_3729 = (in_do&_net_2);
   assign  _net_3730 = (in_do&_net_2);
   assign  _net_3731 = (in_do&_net_2);
   assign  _net_3732 = (in_do&_net_2);
   assign  _net_3733 = (in_do&_net_2);
   assign  _net_3734 = (in_do&_net_2);
   assign  _net_3735 = (in_do&_net_2);
   assign  _net_3736 = (in_do&_net_2);
   assign  _net_3737 = (in_do&_net_2);
   assign  _net_3738 = (in_do&_net_2);
   assign  _net_3739 = (in_do&_net_2);
   assign  _net_3740 = (in_do&_net_2);
   assign  _net_3741 = (in_do&_net_2);
   assign  _net_3742 = (in_do&_net_2);
   assign  _net_3743 = (in_do&_net_2);
   assign  _net_3744 = (in_do&_net_2);
   assign  _net_3745 = (in_do&_net_2);
   assign  _net_3746 = (in_do&_net_2);
   assign  _net_3747 = (in_do&_net_2);
   assign  _net_3748 = (in_do&_net_2);
   assign  _net_3749 = (in_do&_net_2);
   assign  _net_3750 = (in_do&_net_2);
   assign  _net_3751 = (in_do&_net_2);
   assign  _net_3752 = (in_do&_net_2);
   assign  _net_3753 = (in_do&_net_2);
   assign  _net_3754 = (in_do&_net_2);
   assign  _net_3755 = (in_do&_net_2);
   assign  _net_3756 = (in_do&_net_2);
   assign  _net_3757 = (in_do&_net_2);
   assign  _net_3758 = (in_do&_net_2);
   assign  _net_3759 = (in_do&_net_2);
   assign  _net_3760 = (in_do&_net_2);
   assign  _net_3761 = (in_do&_net_2);
   assign  _net_3762 = (in_do&_net_2);
   assign  _net_3763 = (in_do&_net_2);
   assign  _net_3764 = (in_do&_net_2);
   assign  _net_3765 = (in_do&_net_2);
   assign  _net_3766 = (in_do&_net_2);
   assign  _net_3767 = (in_do&_net_2);
   assign  _net_3768 = (in_do&_net_2);
   assign  _net_3769 = (in_do&_net_2);
   assign  _net_3770 = (in_do&_net_2);
   assign  _net_3771 = (in_do&_net_2);
   assign  _net_3772 = (in_do&_net_2);
   assign  _net_3773 = (in_do&_net_2);
   assign  _net_3774 = (in_do&_net_2);
   assign  _net_3775 = (in_do&_net_2);
   assign  _net_3776 = (in_do&_net_2);
   assign  _net_3777 = (in_do&_net_2);
   assign  _net_3778 = (in_do&_net_2);
   assign  _net_3779 = (in_do&_net_2);
   assign  _net_3780 = (in_do&_net_2);
   assign  _net_3781 = (in_do&_net_2);
   assign  _net_3782 = (in_do&_net_2);
   assign  _net_3783 = (in_do&_net_2);
   assign  _net_3784 = (in_do&_net_2);
   assign  _net_3785 = (in_do&_net_2);
   assign  _net_3786 = (in_do&_net_2);
   assign  _net_3787 = (in_do&_net_2);
   assign  _net_3788 = (in_do&_net_2);
   assign  _net_3789 = (in_do&_net_2);
   assign  _net_3790 = (in_do&_net_2);
   assign  _net_3791 = (in_do&_net_2);
   assign  _net_3792 = (in_do&_net_2);
   assign  _net_3793 = (in_do&_net_2);
   assign  _net_3794 = (in_do&_net_2);
   assign  _net_3795 = (in_do&_net_2);
   assign  _net_3796 = (in_do&_net_2);
   assign  _net_3797 = (in_do&_net_2);
   assign  _net_3798 = (in_do&_net_2);
   assign  _net_3799 = (in_do&_net_2);
   assign  _net_3800 = (in_do&_net_2);
   assign  _net_3801 = (in_do&_net_2);
   assign  _net_3802 = (in_do&_net_2);
   assign  _net_3803 = (in_do&_net_2);
   assign  _net_3804 = (in_do&_net_2);
   assign  _net_3805 = (in_do&_net_2);
   assign  _net_3806 = (in_do&_net_2);
   assign  _net_3807 = (in_do&_net_2);
   assign  _net_3808 = (in_do&_net_2);
   assign  _net_3809 = (in_do&_net_2);
   assign  _net_3810 = (in_do&_net_2);
   assign  _net_3811 = (in_do&_net_2);
   assign  _net_3812 = (in_do&_net_2);
   assign  _net_3813 = (in_do&_net_2);
   assign  _net_3814 = (in_do&_net_2);
   assign  _net_3815 = (in_do&_net_2);
   assign  _net_3816 = (in_do&_net_2);
   assign  _net_3817 = (in_do&_net_2);
   assign  _net_3818 = (in_do&_net_2);
   assign  _net_3819 = (in_do&_net_2);
   assign  _net_3820 = (in_do&_net_2);
   assign  _net_3821 = (in_do&_net_2);
   assign  _net_3822 = (in_do&_net_2);
   assign  _net_3823 = (in_do&_net_2);
   assign  _net_3824 = (in_do&_net_2);
   assign  _net_3825 = (in_do&_net_2);
   assign  _net_3826 = (in_do&_net_2);
   assign  _net_3827 = (in_do&_net_2);
   assign  _net_3828 = (in_do&_net_2);
   assign  _net_3829 = (in_do&_net_2);
   assign  _net_3830 = (in_do&_net_2);
   assign  _net_3831 = (in_do&_net_2);
   assign  _net_3832 = (in_do&_net_2);
   assign  _net_3833 = (in_do&_net_2);
   assign  _net_3834 = (in_do&_net_2);
   assign  _net_3835 = (in_do&_net_2);
   assign  _net_3836 = (in_do&_net_2);
   assign  _net_3837 = (in_do&_net_2);
   assign  _net_3838 = (in_do&_net_2);
   assign  _net_3839 = (in_do&_net_2);
   assign  _net_3840 = (in_do&_net_2);
   assign  _net_3841 = (in_do&_net_2);
   assign  _net_3842 = (in_do&_net_2);
   assign  _net_3843 = (in_do&_net_2);
   assign  _net_3844 = (in_do&_net_2);
   assign  _net_3845 = (in_do&_net_2);
   assign  _net_3846 = (in_do&_net_2);
   assign  _net_3847 = (in_do&_net_2);
   assign  _net_3848 = (in_do&_net_2);
   assign  _net_3849 = (in_do&_net_2);
   assign  _net_3850 = (in_do&_net_2);
   assign  _net_3851 = (in_do&_net_2);
   assign  _net_3852 = (in_do&_net_2);
   assign  _net_3853 = (in_do&_net_2);
   assign  _net_3854 = (in_do&_net_2);
   assign  _net_3855 = (in_do&_net_2);
   assign  _net_3856 = (in_do&_net_2);
   assign  _net_3857 = (in_do&_net_2);
   assign  _net_3858 = (in_do&_net_2);
   assign  _net_3859 = (in_do&_net_2);
   assign  _net_3860 = (in_do&_net_2);
   assign  _net_3861 = (in_do&_net_2);
   assign  _net_3862 = (in_do&_net_2);
   assign  _net_3863 = (in_do&_net_2);
   assign  _net_3864 = (in_do&_net_2);
   assign  _net_3865 = (in_do&_net_2);
   assign  _net_3866 = (in_do&_net_2);
   assign  _net_3867 = (in_do&_net_2);
   assign  _net_3868 = (in_do&_net_2);
   assign  _net_3869 = (in_do&_net_2);
   assign  _net_3870 = (in_do&_net_2);
   assign  _net_3871 = (in_do&_net_2);
   assign  _net_3872 = (in_do&_net_2);
   assign  _net_3873 = (in_do&_net_2);
   assign  _net_3874 = (in_do&_net_2);
   assign  _net_3875 = (in_do&_net_2);
   assign  _net_3876 = (in_do&_net_2);
   assign  _net_3877 = (in_do&_net_2);
   assign  _net_3878 = (in_do&_net_2);
   assign  _net_3879 = (in_do&_net_2);
   assign  _net_3880 = (in_do&_net_2);
   assign  _net_3881 = (in_do&_net_2);
   assign  _net_3882 = (in_do&_net_2);
   assign  _net_3883 = (in_do&_net_2);
   assign  _net_3884 = (in_do&_net_2);
   assign  _net_3885 = (in_do&_net_2);
   assign  _net_3886 = (in_do&_net_2);
   assign  _net_3887 = (in_do&_net_2);
   assign  _net_3888 = (in_do&_net_2);
   assign  _net_3889 = (in_do&_net_2);
   assign  _net_3890 = (in_do&_net_2);
   assign  _net_3891 = (in_do&_net_2);
   assign  _net_3892 = (in_do&_net_2);
   assign  _net_3893 = (in_do&_net_2);
   assign  _net_3894 = (in_do&_net_2);
   assign  _net_3895 = (in_do&_net_2);
   assign  _net_3896 = (in_do&_net_2);
   assign  _net_3897 = (in_do&_net_2);
   assign  _net_3898 = (in_do&_net_2);
   assign  _net_3899 = (in_do&_net_2);
   assign  _net_3900 = (in_do&_net_2);
   assign  _net_3901 = (in_do&_net_2);
   assign  _net_3902 = (in_do&_net_2);
   assign  _net_3903 = (in_do&_net_2);
   assign  _net_3904 = (in_do&_net_2);
   assign  _net_3905 = (in_do&_net_2);
   assign  _net_3906 = (in_do&_net_2);
   assign  _net_3907 = (in_do&_net_2);
   assign  _net_3908 = (in_do&_net_2);
   assign  _net_3909 = (in_do&_net_2);
   assign  _net_3910 = (in_do&_net_2);
   assign  _net_3911 = (in_do&_net_2);
   assign  _net_3912 = (in_do&_net_2);
   assign  _net_3913 = (in_do&_net_2);
   assign  _net_3914 = (in_do&_net_2);
   assign  _net_3915 = (in_do&_net_2);
   assign  _net_3916 = (in_do&_net_2);
   assign  _net_3917 = (in_do&_net_2);
   assign  _net_3918 = (in_do&_net_2);
   assign  _net_3919 = (in_do&_net_2);
   assign  _net_3920 = (in_do&_net_2);
   assign  _net_3921 = (in_do&_net_2);
   assign  _net_3922 = (in_do&_net_2);
   assign  _net_3923 = (in_do&_net_2);
   assign  _net_3924 = (in_do&_net_2);
   assign  _net_3925 = (in_do&_net_2);
   assign  _net_3926 = (in_do&_net_2);
   assign  _net_3927 = (in_do&_net_2);
   assign  _net_3928 = (in_do&_net_2);
   assign  _net_3929 = (in_do&_net_2);
   assign  _net_3930 = (in_do&_net_2);
   assign  _net_3931 = (in_do&_net_2);
   assign  _net_3932 = (in_do&_net_2);
   assign  _net_3933 = (in_do&_net_2);
   assign  _net_3934 = (in_do&_net_2);
   assign  _net_3935 = (in_do&_net_2);
   assign  _net_3936 = (in_do&_net_2);
   assign  _net_3937 = (in_do&_net_2);
   assign  _net_3938 = (in_do&_net_2);
   assign  _net_3939 = (in_do&_net_2);
   assign  _net_3940 = (in_do&_net_2);
   assign  _net_3941 = (in_do&_net_2);
   assign  _net_3942 = (in_do&_net_2);
   assign  _net_3943 = (in_do&_net_2);
   assign  _net_3944 = (in_do&_net_2);
   assign  _net_3945 = (in_do&_net_2);
   assign  _net_3946 = (in_do&_net_2);
   assign  _net_3947 = (in_do&_net_2);
   assign  _net_3948 = (in_do&_net_2);
   assign  _net_3949 = (in_do&_net_2);
   assign  _net_3950 = (in_do&_net_2);
   assign  _net_3951 = (in_do&_net_2);
   assign  _net_3952 = (in_do&_net_2);
   assign  _net_3953 = (in_do&_net_2);
   assign  _net_3954 = (in_do&_net_2);
   assign  _net_3955 = (in_do&_net_2);
   assign  _net_3956 = (in_do&_net_2);
   assign  _net_3957 = (in_do&_net_2);
   assign  _net_3958 = (in_do&_net_2);
   assign  _net_3959 = (in_do&_net_2);
   assign  _net_3960 = (in_do&_net_2);
   assign  _net_3961 = (in_do&_net_2);
   assign  _net_3962 = (in_do&_net_2);
   assign  _net_3963 = (in_do&_net_2);
   assign  _net_3964 = (in_do&_net_2);
   assign  _net_3965 = (in_do&_net_2);
   assign  _net_3966 = (in_do&_net_2);
   assign  _net_3967 = (in_do&_net_2);
   assign  _net_3968 = (in_do&_net_2);
   assign  _net_3969 = (in_do&_net_2);
   assign  _net_3970 = (in_do&_net_2);
   assign  _net_3971 = (in_do&_net_2);
   assign  _net_3972 = (in_do&_net_2);
   assign  _net_3973 = (in_do&_net_2);
   assign  _net_3974 = (in_do&_net_2);
   assign  _net_3975 = (in_do&_net_2);
   assign  _net_3976 = (in_do&_net_2);
   assign  _net_3977 = (in_do&_net_2);
   assign  _net_3978 = (in_do&_net_2);
   assign  _net_3979 = (in_do&_net_2);
   assign  _net_3980 = (in_do&_net_2);
   assign  _net_3981 = (in_do&_net_2);
   assign  _net_3982 = (in_do&_net_2);
   assign  _net_3983 = (in_do&_net_2);
   assign  _net_3984 = (in_do&_net_2);
   assign  _net_3985 = (in_do&_net_2);
   assign  _net_3986 = (in_do&_net_2);
   assign  _net_3987 = (in_do&_net_2);
   assign  _net_3988 = (in_do&_net_2);
   assign  _net_3989 = (in_do&_net_2);
   assign  _net_3990 = (in_do&_net_2);
   assign  _net_3991 = (in_do&_net_2);
   assign  _net_3992 = (in_do&_net_2);
   assign  _net_3993 = (in_do&_net_2);
   assign  _net_3994 = (sig==1'b0);
   assign  _net_3995 = (in_do&_net_3994);
   assign  _net_3996 = (in_do&_net_3994);
   assign  _net_3997 = (in_do&_net_3994);
   assign  _net_3998 = (in_do&_net_3994);
   assign  _net_3999 = (in_do&_net_3994);
   assign  _net_4000 = (in_do&_net_3994);
   assign  _net_4001 = (in_do&_net_3994);
   assign  _net_4002 = (in_do&_net_3994);
   assign  _net_4003 = (in_do&_net_3994);
   assign  _net_4004 = (in_do&_net_3994);
   assign  _net_4005 = (in_do&_net_3994);
   assign  _net_4006 = (in_do&_net_3994);
   assign  _net_4007 = (in_do&_net_3994);
   assign  _net_4008 = (in_do&_net_3994);
   assign  _net_4009 = (in_do&_net_3994);
   assign  _net_4010 = (in_do&_net_3994);
   assign  _net_4011 = (in_do&_net_3994);
   assign  _net_4012 = (in_do&_net_3994);
   assign  _net_4013 = (in_do&_net_3994);
   assign  _net_4014 = (in_do&_net_3994);
   assign  _net_4015 = (in_do&_net_3994);
   assign  _net_4016 = (in_do&_net_3994);
   assign  _net_4017 = (in_do&_net_3994);
   assign  _net_4018 = (in_do&_net_3994);
   assign  _net_4019 = (in_do&_net_3994);
   assign  _net_4020 = (in_do&_net_3994);
   assign  _net_4021 = (in_do&_net_3994);
   assign  _net_4022 = (in_do&_net_3994);
   assign  _net_4023 = (in_do&_net_3994);
   assign  _net_4024 = (in_do&_net_3994);
   assign  _net_4025 = (in_do&_net_3994);
   assign  _net_4026 = (in_do&_net_3994);
   assign  _net_4027 = (in_do&_net_3994);
   assign  _net_4028 = (in_do&_net_3994);
   assign  _net_4029 = (in_do&_net_3994);
   assign  _net_4030 = (in_do&_net_3994);
   assign  _net_4031 = (in_do&_net_3994);
   assign  _net_4032 = (in_do&_net_3994);
   assign  _net_4033 = (in_do&_net_3994);
   assign  _net_4034 = (in_do&_net_3994);
   assign  _net_4035 = (in_do&_net_3994);
   assign  _net_4036 = (in_do&_net_3994);
   assign  _net_4037 = (in_do&_net_3994);
   assign  _net_4038 = (in_do&_net_3994);
   assign  _net_4039 = (in_do&_net_3994);
   assign  _net_4040 = (in_do&_net_3994);
   assign  _net_4041 = (in_do&_net_3994);
   assign  _net_4042 = (in_do&_net_3994);
   assign  _net_4043 = (in_do&_net_3994);
   assign  _net_4044 = (in_do&_net_3994);
   assign  _net_4045 = (in_do&_net_3994);
   assign  _net_4046 = (in_do&_net_3994);
   assign  _net_4047 = (in_do&_net_3994);
   assign  _net_4048 = (in_do&_net_3994);
   assign  _net_4049 = (in_do&_net_3994);
   assign  _net_4050 = (in_do&_net_3994);
   assign  _net_4051 = (in_do&_net_3994);
   assign  _net_4052 = (in_do&_net_3994);
   assign  _net_4053 = (in_do&_net_3994);
   assign  _net_4054 = (in_do&_net_3994);
   assign  _net_4055 = (in_do&_net_3994);
   assign  _net_4056 = (in_do&_net_3994);
   assign  _net_4057 = (in_do&_net_3994);
   assign  _net_4058 = (in_do&_net_3994);
   assign  _net_4059 = (in_do&_net_3994);
   assign  _net_4060 = (in_do&_net_3994);
   assign  _net_4061 = (in_do&_net_3994);
   assign  _net_4062 = (in_do&_net_3994);
   assign  _net_4063 = (in_do&_net_3994);
   assign  _net_4064 = (in_do&_net_3994);
   assign  _net_4065 = (in_do&_net_3994);
   assign  _net_4066 = (in_do&_net_3994);
   assign  _net_4067 = (in_do&_net_3994);
   assign  _net_4068 = (in_do&_net_3994);
   assign  _net_4069 = (in_do&_net_3994);
   assign  _net_4070 = (in_do&_net_3994);
   assign  _net_4071 = (in_do&_net_3994);
   assign  _net_4072 = (in_do&_net_3994);
   assign  _net_4073 = (in_do&_net_3994);
   assign  _net_4074 = (in_do&_net_3994);
   assign  _net_4075 = (in_do&_net_3994);
   assign  _net_4076 = (in_do&_net_3994);
   assign  _net_4077 = (in_do&_net_3994);
   assign  _net_4078 = (in_do&_net_3994);
   assign  _net_4079 = (in_do&_net_3994);
   assign  _net_4080 = (in_do&_net_3994);
   assign  _net_4081 = (in_do&_net_3994);
   assign  _net_4082 = (in_do&_net_3994);
   assign  _net_4083 = (in_do&_net_3994);
   assign  _net_4084 = (in_do&_net_3994);
   assign  _net_4085 = (in_do&_net_3994);
   assign  _net_4086 = (in_do&_net_3994);
   assign  _net_4087 = (in_do&_net_3994);
   assign  _net_4088 = (in_do&_net_3994);
   assign  _net_4089 = (in_do&_net_3994);
   assign  _net_4090 = (in_do&_net_3994);
   assign  _net_4091 = (in_do&_net_3994);
   assign  _net_4092 = (in_do&_net_3994);
   assign  _net_4093 = (in_do&_net_3994);
   assign  _net_4094 = (in_do&_net_3994);
   assign  _net_4095 = (in_do&_net_3994);
   assign  _net_4096 = (in_do&_net_3994);
   assign  _net_4097 = (in_do&_net_3994);
   assign  _net_4098 = (in_do&_net_3994);
   assign  _net_4099 = (in_do&_net_3994);
   assign  _net_4100 = (in_do&_net_3994);
   assign  _net_4101 = (in_do&_net_3994);
   assign  _net_4102 = (in_do&_net_3994);
   assign  _net_4103 = (in_do&_net_3994);
   assign  _net_4104 = (in_do&_net_3994);
   assign  _net_4105 = (in_do&_net_3994);
   assign  _net_4106 = (in_do&_net_3994);
   assign  _net_4107 = (in_do&_net_3994);
   assign  _net_4108 = (in_do&_net_3994);
   assign  _net_4109 = (in_do&_net_3994);
   assign  _net_4110 = (in_do&_net_3994);
   assign  _net_4111 = (in_do&_net_3994);
   assign  _net_4112 = (in_do&_net_3994);
   assign  _net_4113 = (in_do&_net_3994);
   assign  _net_4114 = (in_do&_net_3994);
   assign  _net_4115 = (in_do&_net_3994);
   assign  _net_4116 = (in_do&_net_3994);
   assign  _net_4117 = (in_do&_net_3994);
   assign  _net_4118 = (in_do&_net_3994);
   assign  _net_4119 = (in_do&_net_3994);
   assign  _net_4120 = (in_do&_net_3994);
   assign  _net_4121 = (in_do&_net_3994);
   assign  _net_4122 = (in_do&_net_3994);
   assign  _net_4123 = (in_do&_net_3994);
   assign  _net_4124 = (in_do&_net_3994);
   assign  _net_4125 = (in_do&_net_3994);
   assign  _net_4126 = (in_do&_net_3994);
   assign  _net_4127 = (in_do&_net_3994);
   assign  _net_4128 = (in_do&_net_3994);
   assign  _net_4129 = (in_do&_net_3994);
   assign  _net_4130 = (in_do&_net_3994);
   assign  _net_4131 = (in_do&_net_3994);
   assign  _net_4132 = (in_do&_net_3994);
   assign  _net_4133 = (in_do&_net_3994);
   assign  _net_4134 = (in_do&_net_3994);
   assign  _net_4135 = (in_do&_net_3994);
   assign  _net_4136 = (in_do&_net_3994);
   assign  _net_4137 = (in_do&_net_3994);
   assign  _net_4138 = (in_do&_net_3994);
   assign  _net_4139 = (in_do&_net_3994);
   assign  _net_4140 = (in_do&_net_3994);
   assign  _net_4141 = (in_do&_net_3994);
   assign  _net_4142 = (in_do&_net_3994);
   assign  _net_4143 = (in_do&_net_3994);
   assign  _net_4144 = (in_do&_net_3994);
   assign  _net_4145 = (in_do&_net_3994);
   assign  _net_4146 = (in_do&_net_3994);
   assign  _net_4147 = (in_do&_net_3994);
   assign  _net_4148 = (in_do&_net_3994);
   assign  _net_4149 = (in_do&_net_3994);
   assign  _net_4150 = (in_do&_net_3994);
   assign  _net_4151 = (in_do&_net_3994);
   assign  _net_4152 = (in_do&_net_3994);
   assign  _net_4153 = (in_do&_net_3994);
   assign  _net_4154 = (in_do&_net_3994);
   assign  _net_4155 = (in_do&_net_3994);
   assign  _net_4156 = (in_do&_net_3994);
   assign  _net_4157 = (in_do&_net_3994);
   assign  _net_4158 = (in_do&_net_3994);
   assign  _net_4159 = (in_do&_net_3994);
   assign  _net_4160 = (in_do&_net_3994);
   assign  _net_4161 = (in_do&_net_3994);
   assign  _net_4162 = (in_do&_net_3994);
   assign  _net_4163 = (in_do&_net_3994);
   assign  _net_4164 = (in_do&_net_3994);
   assign  _net_4165 = (in_do&_net_3994);
   assign  _net_4166 = (in_do&_net_3994);
   assign  _net_4167 = (in_do&_net_3994);
   assign  _net_4168 = (in_do&_net_3994);
   assign  _net_4169 = (in_do&_net_3994);
   assign  _net_4170 = (in_do&_net_3994);
   assign  _net_4171 = (in_do&_net_3994);
   assign  _net_4172 = (in_do&_net_3994);
   assign  _net_4173 = (in_do&_net_3994);
   assign  _net_4174 = (in_do&_net_3994);
   assign  _net_4175 = (in_do&_net_3994);
   assign  _net_4176 = (in_do&_net_3994);
   assign  _net_4177 = (in_do&_net_3994);
   assign  _net_4178 = (in_do&_net_3994);
   assign  _net_4179 = (in_do&_net_3994);
   assign  _net_4180 = (in_do&_net_3994);
   assign  _net_4181 = (in_do&_net_3994);
   assign  _net_4182 = (in_do&_net_3994);
   assign  _net_4183 = (in_do&_net_3994);
   assign  _net_4184 = (in_do&_net_3994);
   assign  _net_4185 = (in_do&_net_3994);
   assign  _net_4186 = (in_do&_net_3994);
   assign  _net_4187 = (in_do&_net_3994);
   assign  _net_4188 = (in_do&_net_3994);
   assign  _net_4189 = (in_do&_net_3994);
   assign  _net_4190 = (in_do&_net_3994);
   assign  _net_4191 = (in_do&_net_3994);
   assign  _net_4192 = (in_do&_net_3994);
   assign  _net_4193 = (in_do&_net_3994);
   assign  _net_4194 = (in_do&_net_3994);
   assign  _net_4195 = (in_do&_net_3994);
   assign  _net_4196 = (in_do&_net_3994);
   assign  _net_4197 = (in_do&_net_3994);
   assign  _net_4198 = (in_do&_net_3994);
   assign  _net_4199 = (in_do&_net_3994);
   assign  _net_4200 = (in_do&_net_3994);
   assign  _net_4201 = (in_do&_net_3994);
   assign  _net_4202 = (in_do&_net_3994);
   assign  _net_4203 = (in_do&_net_3994);
   assign  _net_4204 = (in_do&_net_3994);
   assign  _net_4205 = (in_do&_net_3994);
   assign  _net_4206 = (in_do&_net_3994);
   assign  _net_4207 = (in_do&_net_3994);
   assign  _net_4208 = (in_do&_net_3994);
   assign  _net_4209 = (in_do&_net_3994);
   assign  _net_4210 = (in_do&_net_3994);
   assign  _net_4211 = (in_do&_net_3994);
   assign  _net_4212 = (in_do&_net_3994);
   assign  _net_4213 = (in_do&_net_3994);
   assign  _net_4214 = (in_do&_net_3994);
   assign  _net_4215 = (in_do&_net_3994);
   assign  _net_4216 = (in_do&_net_3994);
   assign  _net_4217 = (in_do&_net_3994);
   assign  _net_4218 = (in_do&_net_3994);
   assign  _net_4219 = (in_do&_net_3994);
   assign  _net_4220 = (in_do&_net_3994);
   assign  _net_4221 = (in_do&_net_3994);
   assign  _net_4222 = (in_do&_net_3994);
   assign  _net_4223 = (in_do&_net_3994);
   assign  _net_4224 = (in_do&_net_3994);
   assign  _net_4225 = (in_do&_net_3994);
   assign  _net_4226 = (in_do&_net_3994);
   assign  _net_4227 = (in_do&_net_3994);
   assign  _net_4228 = (in_do&_net_3994);
   assign  _net_4229 = (in_do&_net_3994);
   assign  _net_4230 = (in_do&_net_3994);
   assign  _net_4231 = (in_do&_net_3994);
   assign  _net_4232 = (in_do&_net_3994);
   assign  _net_4233 = (in_do&_net_3994);
   assign  _net_4234 = (in_do&_net_3994);
   assign  _net_4235 = (in_do&_net_3994);
   assign  _net_4236 = (in_do&_net_3994);
   assign  _net_4237 = (in_do&_net_3994);
   assign  _net_4238 = (in_do&_net_3994);
   assign  _net_4239 = (in_do&_net_3994);
   assign  _net_4240 = (in_do&_net_3994);
   assign  _net_4241 = (in_do&_net_3994);
   assign  _net_4242 = (in_do&_net_3994);
   assign  _net_4243 = (in_do&_net_3994);
   assign  _net_4244 = (in_do&_net_3994);
   assign  _net_4245 = (in_do&_net_3994);
   assign  _net_4246 = (in_do&_net_3994);
   assign  _net_4247 = (in_do&_net_3994);
   assign  _net_4248 = (in_do&_net_3994);
   assign  _net_4249 = (in_do&_net_3994);
   assign  _net_4250 = (in_do&_net_3994);
   assign  _net_4251 = (in_do&_net_3994);
   assign  _net_4252 = (in_do&_net_3994);
   assign  _net_4253 = (in_do&_net_3994);
   assign  _net_4254 = (in_do&_net_3994);
   assign  _net_4255 = (in_do&_net_3994);
   assign  _net_4256 = (in_do&_net_3994);
   assign  _net_4257 = (in_do&_net_3994);
   assign  _net_4258 = (in_do&_net_3994);
   assign  _net_4259 = (in_do&_net_3994);
   assign  _net_4260 = (in_do&_net_3994);
   assign  _net_4261 = (in_do&_net_3994);
   assign  _net_4262 = (in_do&_net_3994);
   assign  _net_4263 = (in_do&_net_3994);
   assign  _net_4264 = (in_do&_net_3994);
   assign  _net_4265 = (in_do&_net_3994);
   assign  _net_4266 = (in_do&_net_3994);
   assign  _net_4267 = (in_do&_net_3994);
   assign  _net_4268 = (in_do&_net_3994);
   assign  _net_4269 = (in_do&_net_3994);
   assign  _net_4270 = (in_do&_net_3994);
   assign  _net_4271 = (in_do&_net_3994);
   assign  _net_4272 = (in_do&_net_3994);
   assign  _net_4273 = (in_do&_net_3994);
   assign  _net_4274 = (in_do&_net_3994);
   assign  _net_4275 = (in_do&_net_3994);
   assign  _net_4276 = (in_do&_net_3994);
   assign  _net_4277 = (in_do&_net_3994);
   assign  _net_4278 = (in_do&_net_3994);
   assign  _net_4279 = (in_do&_net_3994);
   assign  _net_4280 = (in_do&_net_3994);
   assign  _net_4281 = (in_do&_net_3994);
   assign  _net_4282 = (in_do&_net_3994);
   assign  _net_4283 = (in_do&_net_3994);
   assign  _net_4284 = (in_do&_net_3994);
   assign  _net_4285 = (in_do&_net_3994);
   assign  _net_4286 = (in_do&_net_3994);
   assign  _net_4287 = (in_do&_net_3994);
   assign  _net_4288 = (in_do&_net_3994);
   assign  _net_4289 = (in_do&_net_3994);
   assign  _net_4290 = (in_do&_net_3994);
   assign  _net_4291 = (in_do&_net_3994);
   assign  _net_4292 = (in_do&_net_3994);
   assign  _net_4293 = (in_do&_net_3994);
   assign  _net_4294 = (in_do&_net_3994);
   assign  _net_4295 = (in_do&_net_3994);
   assign  _net_4296 = (in_do&_net_3994);
   assign  _net_4297 = (in_do&_net_3994);
   assign  _net_4298 = (in_do&_net_3994);
   assign  _net_4299 = (in_do&_net_3994);
   assign  _net_4300 = (in_do&_net_3994);
   assign  _net_4301 = (in_do&_net_3994);
   assign  _net_4302 = (in_do&_net_3994);
   assign  _net_4303 = (in_do&_net_3994);
   assign  _net_4304 = (in_do&_net_3994);
   assign  _net_4305 = (in_do&_net_3994);
   assign  _net_4306 = (in_do&_net_3994);
   assign  _net_4307 = (in_do&_net_3994);
   assign  _net_4308 = (in_do&_net_3994);
   assign  _net_4309 = (in_do&_net_3994);
   assign  _net_4310 = (in_do&_net_3994);
   assign  _net_4311 = (in_do&_net_3994);
   assign  _net_4312 = (in_do&_net_3994);
   assign  _net_4313 = (in_do&_net_3994);
   assign  _net_4314 = (in_do&_net_3994);
   assign  _net_4315 = (in_do&_net_3994);
   assign  _net_4316 = (in_do&_net_3994);
   assign  _net_4317 = (in_do&_net_3994);
   assign  _net_4318 = (in_do&_net_3994);
   assign  _net_4319 = (in_do&_net_3994);
   assign  _net_4320 = (in_do&_net_3994);
   assign  _net_4321 = (in_do&_net_3994);
   assign  _net_4322 = (in_do&_net_3994);
   assign  _net_4323 = (in_do&_net_3994);
   assign  _net_4324 = (in_do&_net_3994);
   assign  _net_4325 = (in_do&_net_3994);
   assign  _net_4326 = (in_do&_net_3994);
   assign  _net_4327 = (in_do&_net_3994);
   assign  _net_4328 = (in_do&_net_3994);
   assign  _net_4329 = (in_do&_net_3994);
   assign  _net_4330 = (in_do&_net_3994);
   assign  _net_4331 = (in_do&_net_3994);
   assign  _net_4332 = (in_do&_net_3994);
   assign  _net_4333 = (in_do&_net_3994);
   assign  _net_4334 = (in_do&_net_3994);
   assign  _net_4335 = (in_do&_net_3994);
   assign  _net_4336 = (in_do&_net_3994);
   assign  _net_4337 = (in_do&_net_3994);
   assign  _net_4338 = (in_do&_net_3994);
   assign  _net_4339 = (in_do&_net_3994);
   assign  _net_4340 = (in_do&_net_3994);
   assign  _net_4341 = (in_do&_net_3994);
   assign  _net_4342 = (in_do&_net_3994);
   assign  _net_4343 = (in_do&_net_3994);
   assign  _net_4344 = (in_do&_net_3994);
   assign  _net_4345 = (in_do&_net_3994);
   assign  _net_4346 = (in_do&_net_3994);
   assign  _net_4347 = (in_do&_net_3994);
   assign  _net_4348 = (in_do&_net_3994);
   assign  _net_4349 = (in_do&_net_3994);
   assign  _net_4350 = (in_do&_net_3994);
   assign  _net_4351 = (in_do&_net_3994);
   assign  _net_4352 = (in_do&_net_3994);
   assign  _net_4353 = (in_do&_net_3994);
   assign  _net_4354 = (in_do&_net_3994);
   assign  _net_4355 = (in_do&_net_3994);
   assign  _net_4356 = (in_do&_net_3994);
   assign  _net_4357 = (in_do&_net_3994);
   assign  _net_4358 = (in_do&_net_3994);
   assign  _net_4359 = (in_do&_net_3994);
   assign  _net_4360 = (in_do&_net_3994);
   assign  _net_4361 = (in_do&_net_3994);
   assign  _net_4362 = (in_do&_net_3994);
   assign  _net_4363 = (in_do&_net_3994);
   assign  _net_4364 = (in_do&_net_3994);
   assign  _net_4365 = (in_do&_net_3994);
   assign  _net_4366 = (in_do&_net_3994);
   assign  _net_4367 = (in_do&_net_3994);
   assign  _net_4368 = (in_do&_net_3994);
   assign  _net_4369 = (in_do&_net_3994);
   assign  _net_4370 = (in_do&_net_3994);
   assign  _net_4371 = (in_do&_net_3994);
   assign  _net_4372 = (in_do&_net_3994);
   assign  _net_4373 = (in_do&_net_3994);
   assign  _net_4374 = (in_do&_net_3994);
   assign  _net_4375 = (in_do&_net_3994);
   assign  _net_4376 = (in_do&_net_3994);
   assign  _net_4377 = (in_do&_net_3994);
   assign  _net_4378 = (in_do&_net_3994);
   assign  _net_4379 = (in_do&_net_3994);
   assign  _net_4380 = (in_do&_net_3994);
   assign  _net_4381 = (in_do&_net_3994);
   assign  _net_4382 = (in_do&_net_3994);
   assign  _net_4383 = (in_do&_net_3994);
   assign  _net_4384 = (in_do&_net_3994);
   assign  _net_4385 = (in_do&_net_3994);
   assign  _net_4386 = (in_do&_net_3994);
   assign  _net_4387 = (in_do&_net_3994);
   assign  _net_4388 = (in_do&_net_3994);
   assign  _net_4389 = (in_do&_net_3994);
   assign  _net_4390 = (in_do&_net_3994);
   assign  _net_4391 = (in_do&_net_3994);
   assign  _net_4392 = (in_do&_net_3994);
   assign  _net_4393 = (in_do&_net_3994);
   assign  _net_4394 = (in_do&_net_3994);
   assign  _net_4395 = (in_do&_net_3994);
   assign  _net_4396 = (in_do&_net_3994);
   assign  _net_4397 = (in_do&_net_3994);
   assign  _net_4398 = (in_do&_net_3994);
   assign  _net_4399 = (in_do&_net_3994);
   assign  _net_4400 = (in_do&_net_3994);
   assign  _net_4401 = (in_do&_net_3994);
   assign  _net_4402 = (in_do&_net_3994);
   assign  _net_4403 = (in_do&_net_3994);
   assign  _net_4404 = (in_do&_net_3994);
   assign  _net_4405 = (in_do&_net_3994);
   assign  _net_4406 = (in_do&_net_3994);
   assign  _net_4407 = (in_do&_net_3994);
   assign  _net_4408 = (in_do&_net_3994);
   assign  _net_4409 = (in_do&_net_3994);
   assign  _net_4410 = (in_do&_net_3994);
   assign  _net_4411 = (in_do&_net_3994);
   assign  _net_4412 = (in_do&_net_3994);
   assign  _net_4413 = (in_do&_net_3994);
   assign  _net_4414 = (in_do&_net_3994);
   assign  _net_4415 = (in_do&_net_3994);
   assign  _net_4416 = (in_do&_net_3994);
   assign  _net_4417 = (in_do&_net_3994);
   assign  _net_4418 = (in_do&_net_3994);
   assign  _net_4419 = (in_do&_net_3994);
   assign  _net_4420 = (in_do&_net_3994);
   assign  _net_4421 = (in_do&_net_3994);
   assign  _net_4422 = (in_do&_net_3994);
   assign  _net_4423 = (in_do&_net_3994);
   assign  _net_4424 = (in_do&_net_3994);
   assign  _net_4425 = (in_do&_net_3994);
   assign  _net_4426 = (in_do&_net_3994);
   assign  _net_4427 = (in_do&_net_3994);
   assign  _net_4428 = (in_do&_net_3994);
   assign  _net_4429 = (in_do&_net_3994);
   assign  _net_4430 = (in_do&_net_3994);
   assign  _net_4431 = (in_do&_net_3994);
   assign  _net_4432 = (in_do&_net_3994);
   assign  _net_4433 = (in_do&_net_3994);
   assign  _net_4434 = (in_do&_net_3994);
   assign  _net_4435 = (in_do&_net_3994);
   assign  _net_4436 = (in_do&_net_3994);
   assign  _net_4437 = (in_do&_net_3994);
   assign  _net_4438 = (in_do&_net_3994);
   assign  _net_4439 = (in_do&_net_3994);
   assign  _net_4440 = (in_do&_net_3994);
   assign  _net_4441 = (in_do&_net_3994);
   assign  _net_4442 = (in_do&_net_3994);
   assign  _net_4443 = (in_do&_net_3994);
   assign  _net_4444 = (in_do&_net_3994);
   assign  _net_4445 = (in_do&_net_3994);
   assign  _net_4446 = (in_do&_net_3994);
   assign  _net_4447 = (in_do&_net_3994);
   assign  _net_4448 = (in_do&_net_3994);
   assign  _net_4449 = (in_do&_net_3994);
   assign  _net_4450 = (in_do&_net_3994);
   assign  _net_4451 = (in_do&_net_3994);
   assign  _net_4452 = (in_do&_net_3994);
   assign  _net_4453 = (in_do&_net_3994);
   assign  _net_4454 = (in_do&_net_3994);
   assign  _net_4455 = (in_do&_net_3994);
   assign  _net_4456 = (in_do&_net_3994);
   assign  _net_4457 = (in_do&_net_3994);
   assign  _net_4458 = (in_do&_net_3994);
   assign  _net_4459 = (in_do&_net_3994);
   assign  _net_4460 = (in_do&_net_3994);
   assign  _net_4461 = (in_do&_net_3994);
   assign  _net_4462 = (in_do&_net_3994);
   assign  _net_4463 = (in_do&_net_3994);
   assign  _net_4464 = (in_do&_net_3994);
   assign  _net_4465 = (in_do&_net_3994);
   assign  _net_4466 = (in_do&_net_3994);
   assign  _net_4467 = (in_do&_net_3994);
   assign  _net_4468 = (in_do&_net_3994);
   assign  _net_4469 = (in_do&_net_3994);
   assign  _net_4470 = (in_do&_net_3994);
   assign  _net_4471 = (in_do&_net_3994);
   assign  _net_4472 = (in_do&_net_3994);
   assign  _net_4473 = (in_do&_net_3994);
   assign  _net_4474 = (in_do&_net_3994);
   assign  _net_4475 = (in_do&_net_3994);
   assign  _net_4476 = (in_do&_net_3994);
   assign  _net_4477 = (in_do&_net_3994);
   assign  _net_4478 = (in_do&_net_3994);
   assign  _net_4479 = (in_do&_net_3994);
   assign  _net_4480 = (in_do&_net_3994);
   assign  _net_4481 = (in_do&_net_3994);
   assign  _net_4482 = (in_do&_net_3994);
   assign  _net_4483 = (in_do&_net_3994);
   assign  _net_4484 = (in_do&_net_3994);
   assign  _net_4485 = (in_do&_net_3994);
   assign  _net_4486 = (in_do&_net_3994);
   assign  _net_4487 = (in_do&_net_3994);
   assign  _net_4488 = (in_do&_net_3994);
   assign  _net_4489 = (in_do&_net_3994);
   assign  _net_4490 = (in_do&_net_3994);
   assign  _net_4491 = (in_do&_net_3994);
   assign  _net_4492 = (in_do&_net_3994);
   assign  _net_4493 = (in_do&_net_3994);
   assign  _net_4494 = (in_do&_net_3994);
   assign  _net_4495 = (in_do&_net_3994);
   assign  _net_4496 = (in_do&_net_3994);
   assign  _net_4497 = (in_do&_net_3994);
   assign  _net_4498 = (in_do&_net_3994);
   assign  _net_4499 = (in_do&_net_3994);
   assign  _net_4500 = (in_do&_net_3994);
   assign  _net_4501 = (in_do&_net_3994);
   assign  _net_4502 = (in_do&_net_3994);
   assign  _net_4503 = (in_do&_net_3994);
   assign  _net_4504 = (in_do&_net_3994);
   assign  _net_4505 = (in_do&_net_3994);
   assign  _net_4506 = (in_do&_net_3994);
   assign  _net_4507 = (in_do&_net_3994);
   assign  _net_4508 = (in_do&_net_3994);
   assign  _net_4509 = (in_do&_net_3994);
   assign  _net_4510 = (in_do&_net_3994);
   assign  _net_4511 = (in_do&_net_3994);
   assign  _net_4512 = (in_do&_net_3994);
   assign  _net_4513 = (in_do&_net_3994);
   assign  _net_4514 = (in_do&_net_3994);
   assign  _net_4515 = (in_do&_net_3994);
   assign  _net_4516 = (in_do&_net_3994);
   assign  _net_4517 = (in_do&_net_3994);
   assign  _net_4518 = (in_do&_net_3994);
   assign  _net_4519 = (in_do&_net_3994);
   assign  _net_4520 = (in_do&_net_3994);
   assign  _net_4521 = (in_do&_net_3994);
   assign  _net_4522 = (in_do&_net_3994);
   assign  _net_4523 = (in_do&_net_3994);
   assign  _net_4524 = (in_do&_net_3994);
   assign  _net_4525 = (in_do&_net_3994);
   assign  _net_4526 = (in_do&_net_3994);
   assign  _net_4527 = (in_do&_net_3994);
   assign  _net_4528 = (in_do&_net_3994);
   assign  _net_4529 = (in_do&_net_3994);
   assign  _net_4530 = (in_do&_net_3994);
   assign  _net_4531 = (in_do&_net_3994);
   assign  _net_4532 = (in_do&_net_3994);
   assign  _net_4533 = (in_do&_net_3994);
   assign  _net_4534 = (in_do&_net_3994);
   assign  _net_4535 = (in_do&_net_3994);
   assign  _net_4536 = (in_do&_net_3994);
   assign  _net_4537 = (in_do&_net_3994);
   assign  _net_4538 = (in_do&_net_3994);
   assign  _net_4539 = (in_do&_net_3994);
   assign  _net_4540 = (in_do&_net_3994);
   assign  _net_4541 = (in_do&_net_3994);
   assign  _net_4542 = (in_do&_net_3994);
   assign  _net_4543 = (in_do&_net_3994);
   assign  _net_4544 = (in_do&_net_3994);
   assign  _net_4545 = (in_do&_net_3994);
   assign  _net_4546 = (in_do&_net_3994);
   assign  _net_4547 = (in_do&_net_3994);
   assign  _net_4548 = (in_do&_net_3994);
   assign  _net_4549 = (in_do&_net_3994);
   assign  _net_4550 = (in_do&_net_3994);
   assign  _net_4551 = (in_do&_net_3994);
   assign  _net_4552 = (in_do&_net_3994);
   assign  _net_4553 = (in_do&_net_3994);
   assign  _net_4554 = (in_do&_net_3994);
   assign  _net_4555 = (in_do&_net_3994);
   assign  _net_4556 = (in_do&_net_3994);
   assign  _net_4557 = (in_do&_net_3994);
   assign  _net_4558 = (in_do&_net_3994);
   assign  _net_4559 = (in_do&_net_3994);
   assign  _net_4560 = (in_do&_net_3994);
   assign  _net_4561 = (in_do&_net_3994);
   assign  _net_4562 = (in_do&_net_3994);
   assign  _net_4563 = (in_do&_net_3994);
   assign  _net_4564 = (in_do&_net_3994);
   assign  _net_4565 = (in_do&_net_3994);
   assign  _net_4566 = (in_do&_net_3994);
   assign  _net_4567 = (in_do&_net_3994);
   assign  _net_4568 = (in_do&_net_3994);
   assign  _net_4569 = (in_do&_net_3994);
   assign  _net_4570 = (in_do&_net_3994);
   assign  _net_4571 = (in_do&_net_3994);
   assign  _net_4572 = (in_do&_net_3994);
   assign  _net_4573 = (in_do&_net_3994);
   assign  _net_4574 = (in_do&_net_3994);
   assign  _net_4575 = (in_do&_net_3994);
   assign  _net_4576 = (in_do&_net_3994);
   assign  _net_4577 = (in_do&_net_3994);
   assign  _net_4578 = (in_do&_net_3994);
   assign  _net_4579 = (in_do&_net_3994);
   assign  _net_4580 = (in_do&_net_3994);
   assign  _net_4581 = (in_do&_net_3994);
   assign  _net_4582 = (in_do&_net_3994);
   assign  _net_4583 = (in_do&_net_3994);
   assign  _net_4584 = (in_do&_net_3994);
   assign  _net_4585 = (in_do&_net_3994);
   assign  _net_4586 = (in_do&_net_3994);
   assign  _net_4587 = (in_do&_net_3994);
   assign  _net_4588 = (in_do&_net_3994);
   assign  _net_4589 = (in_do&_net_3994);
   assign  _net_4590 = (in_do&_net_3994);
   assign  _net_4591 = (in_do&_net_3994);
   assign  _net_4592 = (in_do&_net_3994);
   assign  _net_4593 = (in_do&_net_3994);
   assign  _net_4594 = (in_do&_net_3994);
   assign  _net_4595 = (in_do&_net_3994);
   assign  _net_4596 = (in_do&_net_3994);
   assign  _net_4597 = (in_do&_net_3994);
   assign  _net_4598 = (in_do&_net_3994);
   assign  _net_4599 = (in_do&_net_3994);
   assign  _net_4600 = (in_do&_net_3994);
   assign  _net_4601 = (in_do&_net_3994);
   assign  _net_4602 = (in_do&_net_3994);
   assign  _net_4603 = (in_do&_net_3994);
   assign  _net_4604 = (in_do&_net_3994);
   assign  _net_4605 = (in_do&_net_3994);
   assign  _net_4606 = (in_do&_net_3994);
   assign  _net_4607 = (in_do&_net_3994);
   assign  _net_4608 = (in_do&_net_3994);
   assign  _net_4609 = (in_do&_net_3994);
   assign  _net_4610 = (in_do&_net_3994);
   assign  _net_4611 = (in_do&_net_3994);
   assign  _net_4612 = (in_do&_net_3994);
   assign  _net_4613 = (in_do&_net_3994);
   assign  _net_4614 = (in_do&_net_3994);
   assign  _net_4615 = (in_do&_net_3994);
   assign  _net_4616 = (in_do&_net_3994);
   assign  _net_4617 = (in_do&_net_3994);
   assign  _net_4618 = (in_do&_net_3994);
   assign  _net_4619 = (in_do&_net_3994);
   assign  _net_4620 = (in_do&_net_3994);
   assign  _net_4621 = (in_do&_net_3994);
   assign  _net_4622 = (in_do&_net_3994);
   assign  _net_4623 = (in_do&_net_3994);
   assign  _net_4624 = (in_do&_net_3994);
   assign  _net_4625 = (in_do&_net_3994);
   assign  _net_4626 = (in_do&_net_3994);
   assign  _net_4627 = (in_do&_net_3994);
   assign  _net_4628 = (in_do&_net_3994);
   assign  _net_4629 = (in_do&_net_3994);
   assign  _net_4630 = (in_do&_net_3994);
   assign  _net_4631 = (in_do&_net_3994);
   assign  _net_4632 = (in_do&_net_3994);
   assign  _net_4633 = (in_do&_net_3994);
   assign  _net_4634 = (in_do&_net_3994);
   assign  _net_4635 = (in_do&_net_3994);
   assign  _net_4636 = (in_do&_net_3994);
   assign  _net_4637 = (in_do&_net_3994);
   assign  _net_4638 = (in_do&_net_3994);
   assign  _net_4639 = (in_do&_net_3994);
   assign  _net_4640 = (in_do&_net_3994);
   assign  _net_4641 = (in_do&_net_3994);
   assign  _net_4642 = (in_do&_net_3994);
   assign  _net_4643 = (in_do&_net_3994);
   assign  _net_4644 = (in_do&_net_3994);
   assign  _net_4645 = (in_do&_net_3994);
   assign  _net_4646 = (in_do&_net_3994);
   assign  _net_4647 = (in_do&_net_3994);
   assign  _net_4648 = (in_do&_net_3994);
   assign  _net_4649 = (in_do&_net_3994);
   assign  _net_4650 = (in_do&_net_3994);
   assign  _net_4651 = (in_do&_net_3994);
   assign  _net_4652 = (in_do&_net_3994);
   assign  _net_4653 = (in_do&_net_3994);
   assign  _net_4654 = (in_do&_net_3994);
   assign  _net_4655 = (in_do&_net_3994);
   assign  _net_4656 = (in_do&_net_3994);
   assign  _net_4657 = (in_do&_net_3994);
   assign  _net_4658 = (in_do&_net_3994);
   assign  _net_4659 = (in_do&_net_3994);
   assign  _net_4660 = (in_do&_net_3994);
   assign  _net_4661 = (in_do&_net_3994);
   assign  _net_4662 = (in_do&_net_3994);
   assign  _net_4663 = (in_do&_net_3994);
   assign  _net_4664 = (in_do&_net_3994);
   assign  _net_4665 = (in_do&_net_3994);
   assign  _net_4666 = (in_do&_net_3994);
   assign  _net_4667 = (in_do&_net_3994);
   assign  _net_4668 = (in_do&_net_3994);
   assign  _net_4669 = (in_do&_net_3994);
   assign  _net_4670 = (in_do&_net_3994);
   assign  _net_4671 = (in_do&_net_3994);
   assign  _net_4672 = (in_do&_net_3994);
   assign  _net_4673 = (in_do&_net_3994);
   assign  _net_4674 = (in_do&_net_3994);
   assign  _net_4675 = (in_do&_net_3994);
   assign  _net_4676 = (in_do&_net_3994);
   assign  _net_4677 = (in_do&_net_3994);
   assign  _net_4678 = (in_do&_net_3994);
   assign  _net_4679 = (in_do&_net_3994);
   assign  _net_4680 = (in_do&_net_3994);
   assign  _net_4681 = (in_do&_net_3994);
   assign  _net_4682 = (in_do&_net_3994);
   assign  _net_4683 = (in_do&_net_3994);
   assign  _net_4684 = (in_do&_net_3994);
   assign  _net_4685 = (in_do&_net_3994);
   assign  _net_4686 = (in_do&_net_3994);
   assign  _net_4687 = (in_do&_net_3994);
   assign  _net_4688 = (in_do&_net_3994);
   assign  _net_4689 = (in_do&_net_3994);
   assign  _net_4690 = (in_do&_net_3994);
   assign  _net_4691 = (in_do&_net_3994);
   assign  _net_4692 = (in_do&_net_3994);
   assign  _net_4693 = (in_do&_net_3994);
   assign  _net_4694 = (in_do&_net_3994);
   assign  _net_4695 = (in_do&_net_3994);
   assign  _net_4696 = (in_do&_net_3994);
   assign  _net_4697 = (in_do&_net_3994);
   assign  _net_4698 = (in_do&_net_3994);
   assign  _net_4699 = (in_do&_net_3994);
   assign  _net_4700 = (in_do&_net_3994);
   assign  _net_4701 = (in_do&_net_3994);
   assign  _net_4702 = (in_do&_net_3994);
   assign  _net_4703 = (in_do&_net_3994);
   assign  _net_4704 = (in_do&_net_3994);
   assign  _net_4705 = (in_do&_net_3994);
   assign  _net_4706 = (in_do&_net_3994);
   assign  _net_4707 = (in_do&_net_3994);
   assign  _net_4708 = (in_do&_net_3994);
   assign  _net_4709 = (in_do&_net_3994);
   assign  _net_4710 = (in_do&_net_3994);
   assign  _net_4711 = (in_do&_net_3994);
   assign  _net_4712 = (in_do&_net_3994);
   assign  _net_4713 = (in_do&_net_3994);
   assign  _net_4714 = (in_do&_net_3994);
   assign  _net_4715 = (in_do&_net_3994);
   assign  _net_4716 = (in_do&_net_3994);
   assign  _net_4717 = (in_do&_net_3994);
   assign  _net_4718 = (in_do&_net_3994);
   assign  _net_4719 = (in_do&_net_3994);
   assign  _net_4720 = (in_do&_net_3994);
   assign  _net_4721 = (in_do&_net_3994);
   assign  _net_4722 = (in_do&_net_3994);
   assign  _net_4723 = (in_do&_net_3994);
   assign  _net_4724 = (in_do&_net_3994);
   assign  _net_4725 = (in_do&_net_3994);
   assign  _net_4726 = (in_do&_net_3994);
   assign  _net_4727 = (in_do&_net_3994);
   assign  _net_4728 = (in_do&_net_3994);
   assign  _net_4729 = (in_do&_net_3994);
   assign  _net_4730 = (in_do&_net_3994);
   assign  _net_4731 = (in_do&_net_3994);
   assign  _net_4732 = (in_do&_net_3994);
   assign  _net_4733 = (in_do&_net_3994);
   assign  _net_4734 = (in_do&_net_3994);
   assign  _net_4735 = (in_do&_net_3994);
   assign  _net_4736 = (in_do&_net_3994);
   assign  _net_4737 = (in_do&_net_3994);
   assign  _net_4738 = (in_do&_net_3994);
   assign  _net_4739 = (in_do&_net_3994);
   assign  _net_4740 = (in_do&_net_3994);
   assign  _net_4741 = (in_do&_net_3994);
   assign  _net_4742 = (in_do&_net_3994);
   assign  _net_4743 = (in_do&_net_3994);
   assign  _net_4744 = (in_do&_net_3994);
   assign  _net_4745 = (in_do&_net_3994);
   assign  _net_4746 = (in_do&_net_3994);
   assign  _net_4747 = (in_do&_net_3994);
   assign  _net_4748 = (in_do&_net_3994);
   assign  _net_4749 = (in_do&_net_3994);
   assign  _net_4750 = (in_do&_net_3994);
   assign  _net_4751 = (in_do&_net_3994);
   assign  _net_4752 = (in_do&_net_3994);
   assign  _net_4753 = (in_do&_net_3994);
   assign  _net_4754 = (in_do&_net_3994);
   assign  _net_4755 = (in_do&_net_3994);
   assign  _net_4756 = (in_do&_net_3994);
   assign  _net_4757 = (in_do&_net_3994);
   assign  _net_4758 = (in_do&_net_3994);
   assign  _net_4759 = (in_do&_net_3994);
   assign  _net_4760 = (in_do&_net_3994);
   assign  _net_4761 = (in_do&_net_3994);
   assign  _net_4762 = (in_do&_net_3994);
   assign  _net_4763 = (in_do&_net_3994);
   assign  _net_4764 = (in_do&_net_3994);
   assign  _net_4765 = (in_do&_net_3994);
   assign  _net_4766 = (in_do&_net_3994);
   assign  _net_4767 = (in_do&_net_3994);
   assign  _net_4768 = (in_do&_net_3994);
   assign  _net_4769 = (in_do&_net_3994);
   assign  _net_4770 = (in_do&_net_3994);
   assign  _net_4771 = (in_do&_net_3994);
   assign  _net_4772 = (in_do&_net_3994);
   assign  _net_4773 = (in_do&_net_3994);
   assign  _net_4774 = (in_do&_net_3994);
   assign  _net_4775 = (in_do&_net_3994);
   assign  _net_4776 = (in_do&_net_3994);
   assign  _net_4777 = (in_do&_net_3994);
   assign  _net_4778 = (in_do&_net_3994);
   assign  _net_4779 = (in_do&_net_3994);
   assign  _net_4780 = (in_do&_net_3994);
   assign  _net_4781 = (in_do&_net_3994);
   assign  _net_4782 = (in_do&_net_3994);
   assign  _net_4783 = (in_do&_net_3994);
   assign  _net_4784 = (in_do&_net_3994);
   assign  _net_4785 = (in_do&_net_3994);
   assign  _net_4786 = (in_do&_net_3994);
   assign  _net_4787 = (in_do&_net_3994);
   assign  _net_4788 = (in_do&_net_3994);
   assign  _net_4789 = (in_do&_net_3994);
   assign  _net_4790 = (in_do&_net_3994);
   assign  _net_4791 = (in_do&_net_3994);
   assign  _net_4792 = (in_do&_net_3994);
   assign  _net_4793 = (in_do&_net_3994);
   assign  _net_4794 = (in_do&_net_3994);
   assign  _net_4795 = (in_do&_net_3994);
   assign  _net_4796 = (in_do&_net_3994);
   assign  _net_4797 = (in_do&_net_3994);
   assign  _net_4798 = (in_do&_net_3994);
   assign  _net_4799 = (in_do&_net_3994);
   assign  _net_4800 = (in_do&_net_3994);
   assign  _net_4801 = (in_do&_net_3994);
   assign  _net_4802 = (in_do&_net_3994);
   assign  _net_4803 = (in_do&_net_3994);
   assign  _net_4804 = (in_do&_net_3994);
   assign  _net_4805 = (in_do&_net_3994);
   assign  _net_4806 = (in_do&_net_3994);
   assign  _net_4807 = (in_do&_net_3994);
   assign  _net_4808 = (in_do&_net_3994);
   assign  _net_4809 = (in_do&_net_3994);
   assign  _net_4810 = (in_do&_net_3994);
   assign  _net_4811 = (in_do&_net_3994);
   assign  _net_4812 = (in_do&_net_3994);
   assign  _net_4813 = (in_do&_net_3994);
   assign  _net_4814 = (in_do&_net_3994);
   assign  _net_4815 = (in_do&_net_3994);
   assign  _net_4816 = (in_do&_net_3994);
   assign  _net_4817 = (in_do&_net_3994);
   assign  _net_4818 = (in_do&_net_3994);
   assign  _net_4819 = (in_do&_net_3994);
   assign  _net_4820 = (in_do&_net_3994);
   assign  _net_4821 = (in_do&_net_3994);
   assign  _net_4822 = (in_do&_net_3994);
   assign  _net_4823 = (in_do&_net_3994);
   assign  _net_4824 = (in_do&_net_3994);
   assign  _net_4825 = (in_do&_net_3994);
   assign  _net_4826 = (in_do&_net_3994);
   assign  _net_4827 = (in_do&_net_3994);
   assign  _net_4828 = (in_do&_net_3994);
   assign  _net_4829 = (in_do&_net_3994);
   assign  _net_4830 = (in_do&_net_3994);
   assign  _net_4831 = (in_do&_net_3994);
   assign  _net_4832 = (in_do&_net_3994);
   assign  _net_4833 = (in_do&_net_3994);
   assign  _net_4834 = (in_do&_net_3994);
   assign  _net_4835 = (in_do&_net_3994);
   assign  _net_4836 = (in_do&_net_3994);
   assign  _net_4837 = (in_do&_net_3994);
   assign  _net_4838 = (in_do&_net_3994);
   assign  _net_4839 = (in_do&_net_3994);
   assign  _net_4840 = (in_do&_net_3994);
   assign  _net_4841 = (in_do&_net_3994);
   assign  _net_4842 = (in_do&_net_3994);
   assign  _net_4843 = (in_do&_net_3994);
   assign  _net_4844 = (in_do&_net_3994);
   assign  _net_4845 = (in_do&_net_3994);
   assign  _net_4846 = (in_do&_net_3994);
   assign  _net_4847 = (in_do&_net_3994);
   assign  _net_4848 = (in_do&_net_3994);
   assign  _net_4849 = (in_do&_net_3994);
   assign  _net_4850 = (in_do&_net_3994);
   assign  _net_4851 = (in_do&_net_3994);
   assign  _net_4852 = (in_do&_net_3994);
   assign  _net_4853 = (in_do&_net_3994);
   assign  _net_4854 = (in_do&_net_3994);
   assign  _net_4855 = (in_do&_net_3994);
   assign  _net_4856 = (in_do&_net_3994);
   assign  _net_4857 = (in_do&_net_3994);
   assign  _net_4858 = (in_do&_net_3994);
   assign  _net_4859 = (in_do&_net_3994);
   assign  _net_4860 = (in_do&_net_3994);
   assign  _net_4861 = (in_do&_net_3994);
   assign  _net_4862 = (in_do&_net_3994);
   assign  _net_4863 = (in_do&_net_3994);
   assign  _net_4864 = (in_do&_net_3994);
   assign  _net_4865 = (in_do&_net_3994);
   assign  _net_4866 = (in_do&_net_3994);
   assign  _net_4867 = (in_do&_net_3994);
   assign  _net_4868 = (in_do&_net_3994);
   assign  _net_4869 = (in_do&_net_3994);
   assign  _net_4870 = (in_do&_net_3994);
   assign  _net_4871 = (in_do&_net_3994);
   assign  _net_4872 = (in_do&_net_3994);
   assign  _net_4873 = (in_do&_net_3994);
   assign  _net_4874 = (in_do&_net_3994);
   assign  _net_4875 = (in_do&_net_3994);
   assign  _net_4876 = (in_do&_net_3994);
   assign  _net_4877 = (in_do&_net_3994);
   assign  _net_4878 = (in_do&_net_3994);
   assign  _net_4879 = (in_do&_net_3994);
   assign  _net_4880 = (in_do&_net_3994);
   assign  _net_4881 = (in_do&_net_3994);
   assign  _net_4882 = (in_do&_net_3994);
   assign  _net_4883 = (in_do&_net_3994);
   assign  _net_4884 = (in_do&_net_3994);
   assign  _net_4885 = (in_do&_net_3994);
   assign  _net_4886 = (in_do&_net_3994);
   assign  _net_4887 = (in_do&_net_3994);
   assign  _net_4888 = (in_do&_net_3994);
   assign  _net_4889 = (in_do&_net_3994);
   assign  _net_4890 = (in_do&_net_3994);
   assign  _net_4891 = (in_do&_net_3994);
   assign  _net_4892 = (in_do&_net_3994);
   assign  _net_4893 = (in_do&_net_3994);
   assign  _net_4894 = (in_do&_net_3994);
   assign  _net_4895 = (in_do&_net_3994);
   assign  _net_4896 = (in_do&_net_3994);
   assign  _net_4897 = (in_do&_net_3994);
   assign  _net_4898 = (in_do&_net_3994);
   assign  _net_4899 = (in_do&_net_3994);
   assign  _net_4900 = (in_do&_net_3994);
   assign  _net_4901 = (in_do&_net_3994);
   assign  _net_4902 = (in_do&_net_3994);
   assign  _net_4903 = (in_do&_net_3994);
   assign  _net_4904 = (in_do&_net_3994);
   assign  _net_4905 = (in_do&_net_3994);
   assign  _net_4906 = (in_do&_net_3994);
   assign  _net_4907 = (in_do&_net_3994);
   assign  _net_4908 = (in_do&_net_3994);
   assign  _net_4909 = (in_do&_net_3994);
   assign  _net_4910 = (in_do&_net_3994);
   assign  _net_4911 = (in_do&_net_3994);
   assign  _net_4912 = (in_do&_net_3994);
   assign  _net_4913 = (in_do&_net_3994);
   assign  _net_4914 = (in_do&_net_3994);
   assign  _net_4915 = (in_do&_net_3994);
   assign  _net_4916 = (in_do&_net_3994);
   assign  _net_4917 = (in_do&_net_3994);
   assign  _net_4918 = (in_do&_net_3994);
   assign  _net_4919 = (in_do&_net_3994);
   assign  _net_4920 = (in_do&_net_3994);
   assign  _net_4921 = (in_do&_net_3994);
   assign  _net_4922 = (in_do&_net_3994);
   assign  _net_4923 = (in_do&_net_3994);
   assign  _net_4924 = (in_do&_net_3994);
   assign  _net_4925 = (in_do&_net_3994);
   assign  _net_4926 = (in_do&_net_3994);
   assign  _net_4927 = (in_do&_net_3994);
   assign  _net_4928 = (in_do&_net_3994);
   assign  _net_4929 = (in_do&_net_3994);
   assign  _net_4930 = (in_do&_net_3994);
   assign  _net_4931 = (in_do&_net_3994);
   assign  _net_4932 = (in_do&_net_3994);
   assign  _net_4933 = (in_do&_net_3994);
   assign  _net_4934 = (in_do&_net_3994);
   assign  _net_4935 = (in_do&_net_3994);
   assign  _net_4936 = (in_do&_net_3994);
   assign  _net_4937 = (in_do&_net_3994);
   assign  _net_4938 = (in_do&_net_3994);
   assign  _net_4939 = (in_do&_net_3994);
   assign  _net_4940 = (in_do&_net_3994);
   assign  _net_4941 = (in_do&_net_3994);
   assign  _net_4942 = (in_do&_net_3994);
   assign  _net_4943 = (in_do&_net_3994);
   assign  _net_4944 = (in_do&_net_3994);
   assign  _net_4945 = (in_do&_net_3994);
   assign  _net_4946 = (in_do&_net_3994);
   assign  _net_4947 = (in_do&_net_3994);
   assign  _net_4948 = (in_do&_net_3994);
   assign  _net_4949 = (in_do&_net_3994);
   assign  _net_4950 = (in_do&_net_3994);
   assign  _net_4951 = (in_do&_net_3994);
   assign  _net_4952 = (in_do&_net_3994);
   assign  _net_4953 = (in_do&_net_3994);
   assign  _net_4954 = (in_do&_net_3994);
   assign  _net_4955 = (in_do&_net_3994);
   assign  _net_4956 = (in_do&_net_3994);
   assign  _net_4957 = (in_do&_net_3994);
   assign  _net_4958 = (in_do&_net_3994);
   assign  _net_4959 = (in_do&_net_3994);
   assign  _net_4960 = (in_do&_net_3994);
   assign  _net_4961 = (in_do&_net_3994);
   assign  _net_4962 = (in_do&_net_3994);
   assign  _net_4963 = (in_do&_net_3994);
   assign  _net_4964 = (in_do&_net_3994);
   assign  _net_4965 = (in_do&_net_3994);
   assign  _net_4966 = (in_do&_net_3994);
   assign  _net_4967 = (in_do&_net_3994);
   assign  _net_4968 = (in_do&_net_3994);
   assign  _net_4969 = (in_do&_net_3994);
   assign  _net_4970 = (in_do&_net_3994);
   assign  _net_4971 = (in_do&_net_3994);
   assign  _net_4972 = (in_do&_net_3994);
   assign  _net_4973 = (in_do&_net_3994);
   assign  _net_4974 = (in_do&_net_3994);
   assign  _net_4975 = (in_do&_net_3994);
   assign  _net_4976 = (in_do&_net_3994);
   assign  _net_4977 = (in_do&_net_3994);
   assign  _net_4978 = (in_do&_net_3994);
   assign  _net_4979 = (in_do&_net_3994);
   assign  _net_4980 = (in_do&_net_3994);
   assign  _net_4981 = (in_do&_net_3994);
   assign  _net_4982 = (in_do&_net_3994);
   assign  _net_4983 = (in_do&_net_3994);
   assign  _net_4984 = (in_do&_net_3994);
   assign  _net_4985 = (in_do&_net_3994);
   assign  _net_4986 = (in_do&_net_3994);
   assign  _net_4987 = (in_do&_net_3994);
   assign  _net_4988 = (in_do&_net_3994);
   assign  _net_4989 = (in_do&_net_3994);
   assign  _net_4990 = (in_do&_net_3994);
   assign  _net_4991 = (in_do&_net_3994);
   assign  _net_4992 = (in_do&_net_3994);
   assign  _net_4993 = (in_do&_net_3994);
   assign  _net_4994 = (in_do&_net_3994);
   assign  _net_4995 = (in_do&_net_3994);
   assign  _net_4996 = (in_do&_net_3994);
   assign  _net_4997 = (in_do&_net_3994);
   assign  _net_4998 = (in_do&_net_3994);
   assign  _net_4999 = (in_do&_net_3994);
   assign  _net_5000 = (in_do&_net_3994);
   assign  _net_5001 = (in_do&_net_3994);
   assign  _net_5002 = (in_do&_net_3994);
   assign  _net_5003 = (in_do&_net_3994);
   assign  _net_5004 = (in_do&_net_3994);
   assign  _net_5005 = (in_do&_net_3994);
   assign  _net_5006 = (in_do&_net_3994);
   assign  _net_5007 = (in_do&_net_3994);
   assign  _net_5008 = (in_do&_net_3994);
   assign  _net_5009 = (in_do&_net_3994);
   assign  _net_5010 = (in_do&_net_3994);
   assign  _net_5011 = (in_do&_net_3994);
   assign  _net_5012 = (in_do&_net_3994);
   assign  _net_5013 = (in_do&_net_3994);
   assign  _net_5014 = (in_do&_net_3994);
   assign  _net_5015 = (in_do&_net_3994);
   assign  _net_5016 = (in_do&_net_3994);
   assign  _net_5017 = (in_do&_net_3994);
   assign  _net_5018 = (in_do&_net_3994);
   assign  _net_5019 = (in_do&_net_3994);
   assign  _net_5020 = (in_do&_net_3994);
   assign  _net_5021 = (in_do&_net_3994);
   assign  _net_5022 = (in_do&_net_3994);
   assign  _net_5023 = (in_do&_net_3994);
   assign  _net_5024 = (in_do&_net_3994);
   assign  _net_5025 = (in_do&_net_3994);
   assign  _net_5026 = (in_do&_net_3994);
   assign  _net_5027 = (in_do&_net_3994);
   assign  _net_5028 = (in_do&_net_3994);
   assign  _net_5029 = (in_do&_net_3994);
   assign  _net_5030 = (in_do&_net_3994);
   assign  _net_5031 = (in_do&_net_3994);
   assign  _net_5032 = (in_do&_net_3994);
   assign  _net_5033 = (in_do&_net_3994);
   assign  _net_5034 = (in_do&_net_3994);
   assign  _net_5035 = (in_do&_net_3994);
   assign  _net_5036 = (in_do&_net_3994);
   assign  _net_5037 = (in_do&_net_3994);
   assign  _net_5038 = (in_do&_net_3994);
   assign  _net_5039 = (in_do&_net_3994);
   assign  _net_5040 = (in_do&_net_3994);
   assign  _net_5041 = (in_do&_net_3994);
   assign  _net_5042 = (in_do&_net_3994);
   assign  _net_5043 = (in_do&_net_3994);
   assign  _net_5044 = (in_do&_net_3994);
   assign  _net_5045 = (in_do&_net_3994);
   assign  _net_5046 = (in_do&_net_3994);
   assign  _net_5047 = (in_do&_net_3994);
   assign  _net_5048 = (in_do&_net_3994);
   assign  _net_5049 = (in_do&_net_3994);
   assign  _net_5050 = (in_do&_net_3994);
   assign  _net_5051 = (in_do&_net_3994);
   assign  _net_5052 = (in_do&_net_3994);
   assign  _net_5053 = (in_do&_net_3994);
   assign  _net_5054 = (in_do&_net_3994);
   assign  _net_5055 = (in_do&_net_3994);
   assign  _net_5056 = (in_do&_net_3994);
   assign  _net_5057 = (in_do&_net_3994);
   assign  _net_5058 = (in_do&_net_3994);
   assign  _net_5059 = (in_do&_net_3994);
   assign  _net_5060 = (in_do&_net_3994);
   assign  _net_5061 = (in_do&_net_3994);
   assign  _net_5062 = (in_do&_net_3994);
   assign  _net_5063 = (in_do&_net_3994);
   assign  _net_5064 = (in_do&_net_3994);
   assign  _net_5065 = (in_do&_net_3994);
   assign  _net_5066 = (in_do&_net_3994);
   assign  _net_5067 = (in_do&_net_3994);
   assign  _net_5068 = (in_do&_net_3994);
   assign  _net_5069 = (in_do&_net_3994);
   assign  _net_5070 = (in_do&_net_3994);
   assign  _net_5071 = (in_do&_net_3994);
   assign  _net_5072 = (in_do&_net_3994);
   assign  _net_5073 = (in_do&_net_3994);
   assign  _net_5074 = (in_do&_net_3994);
   assign  _net_5075 = (in_do&_net_3994);
   assign  _net_5076 = (in_do&_net_3994);
   assign  _net_5077 = (in_do&_net_3994);
   assign  _net_5078 = (in_do&_net_3994);
   assign  _net_5079 = (in_do&_net_3994);
   assign  _net_5080 = (in_do&_net_3994);
   assign  _net_5081 = (in_do&_net_3994);
   assign  _net_5082 = (in_do&_net_3994);
   assign  _net_5083 = (in_do&_net_3994);
   assign  _net_5084 = (in_do&_net_3994);
   assign  _net_5085 = (in_do&_net_3994);
   assign  _net_5086 = (in_do&_net_3994);
   assign  _net_5087 = (in_do&_net_3994);
   assign  _net_5088 = (in_do&_net_3994);
   assign  _net_5089 = (in_do&_net_3994);
   assign  _net_5090 = (in_do&_net_3994);
   assign  _net_5091 = (in_do&_net_3994);
   assign  _net_5092 = (in_do&_net_3994);
   assign  _net_5093 = (in_do&_net_3994);
   assign  _net_5094 = (in_do&_net_3994);
   assign  _net_5095 = (in_do&_net_3994);
   assign  _net_5096 = (in_do&_net_3994);
   assign  _net_5097 = (in_do&_net_3994);
   assign  _net_5098 = (in_do&_net_3994);
   assign  _net_5099 = (in_do&_net_3994);
   assign  _net_5100 = (in_do&_net_3994);
   assign  _net_5101 = (in_do&_net_3994);
   assign  _net_5102 = (in_do&_net_3994);
   assign  _net_5103 = (in_do&_net_3994);
   assign  _net_5104 = (in_do&_net_3994);
   assign  _net_5105 = (in_do&_net_3994);
   assign  _net_5106 = (in_do&_net_3994);
   assign  _net_5107 = (in_do&_net_3994);
   assign  _net_5108 = (in_do&_net_3994);
   assign  _net_5109 = (in_do&_net_3994);
   assign  _net_5110 = (in_do&_net_3994);
   assign  _net_5111 = (in_do&_net_3994);
   assign  _net_5112 = (in_do&_net_3994);
   assign  _net_5113 = (in_do&_net_3994);
   assign  _net_5114 = (in_do&_net_3994);
   assign  _net_5115 = (in_do&_net_3994);
   assign  _net_5116 = (in_do&_net_3994);
   assign  _net_5117 = (in_do&_net_3994);
   assign  _net_5118 = (in_do&_net_3994);
   assign  _net_5119 = (in_do&_net_3994);
   assign  _net_5120 = (in_do&_net_3994);
   assign  _net_5121 = (in_do&_net_3994);
   assign  _net_5122 = (in_do&_net_3994);
   assign  _net_5123 = (in_do&_net_3994);
   assign  _net_5124 = (in_do&_net_3994);
   assign  _net_5125 = (in_do&_net_3994);
   assign  _net_5126 = (in_do&_net_3994);
   assign  _net_5127 = (in_do&_net_3994);
   assign  _net_5128 = (in_do&_net_3994);
   assign  _net_5129 = (in_do&_net_3994);
   assign  _net_5130 = (in_do&_net_3994);
   assign  _net_5131 = (in_do&_net_3994);
   assign  _net_5132 = (in_do&_net_3994);
   assign  _net_5133 = (in_do&_net_3994);
   assign  _net_5134 = (in_do&_net_3994);
   assign  _net_5135 = (in_do&_net_3994);
   assign  _net_5136 = (in_do&_net_3994);
   assign  _net_5137 = (in_do&_net_3994);
   assign  _net_5138 = (in_do&_net_3994);
   assign  _net_5139 = (in_do&_net_3994);
   assign  _net_5140 = (in_do&_net_3994);
   assign  _net_5141 = (in_do&_net_3994);
   assign  _net_5142 = (in_do&_net_3994);
   assign  _net_5143 = (in_do&_net_3994);
   assign  _net_5144 = (in_do&_net_3994);
   assign  _net_5145 = (in_do&_net_3994);
   assign  _net_5146 = (in_do&_net_3994);
   assign  _net_5147 = (in_do&_net_3994);
   assign  _net_5148 = (in_do&_net_3994);
   assign  _net_5149 = (in_do&_net_3994);
   assign  _net_5150 = (in_do&_net_3994);
   assign  _net_5151 = (in_do&_net_3994);
   assign  _net_5152 = (in_do&_net_3994);
   assign  _net_5153 = (in_do&_net_3994);
   assign  _net_5154 = (in_do&_net_3994);
   assign  _net_5155 = (in_do&_net_3994);
   assign  _net_5156 = (in_do&_net_3994);
   assign  _net_5157 = (in_do&_net_3994);
   assign  _net_5158 = (in_do&_net_3994);
   assign  _net_5159 = (in_do&_net_3994);
   assign  _net_5160 = (in_do&_net_3994);
   assign  _net_5161 = (in_do&_net_3994);
   assign  _net_5162 = (in_do&_net_3994);
   assign  _net_5163 = (in_do&_net_3994);
   assign  _net_5164 = (in_do&_net_3994);
   assign  _net_5165 = (in_do&_net_3994);
   assign  _net_5166 = (in_do&_net_3994);
   assign  _net_5167 = (in_do&_net_3994);
   assign  _net_5168 = (in_do&_net_3994);
   assign  _net_5169 = (in_do&_net_3994);
   assign  _net_5170 = (in_do&_net_3994);
   assign  _net_5171 = (in_do&_net_3994);
   assign  _net_5172 = (in_do&_net_3994);
   assign  _net_5173 = (in_do&_net_3994);
   assign  _net_5174 = (in_do&_net_3994);
   assign  _net_5175 = (in_do&_net_3994);
   assign  _net_5176 = (in_do&_net_3994);
   assign  _net_5177 = (in_do&_net_3994);
   assign  _net_5178 = (in_do&_net_3994);
   assign  _net_5179 = (in_do&_net_3994);
   assign  _net_5180 = (in_do&_net_3994);
   assign  _net_5181 = (in_do&_net_3994);
   assign  _net_5182 = (in_do&_net_3994);
   assign  _net_5183 = (in_do&_net_3994);
   assign  _net_5184 = (in_do&_net_3994);
   assign  _net_5185 = (in_do&_net_3994);
   assign  _net_5186 = (in_do&_net_3994);
   assign  _net_5187 = (in_do&_net_3994);
   assign  _net_5188 = (in_do&_net_3994);
   assign  _net_5189 = (in_do&_net_3994);
   assign  _net_5190 = (in_do&_net_3994);
   assign  _net_5191 = (in_do&_net_3994);
   assign  _net_5192 = (in_do&_net_3994);
   assign  _net_5193 = (in_do&_net_3994);
   assign  _net_5194 = (in_do&_net_3994);
   assign  _net_5195 = (in_do&_net_3994);
   assign  _net_5196 = (in_do&_net_3994);
   assign  _net_5197 = (in_do&_net_3994);
   assign  _net_5198 = (in_do&_net_3994);
   assign  _net_5199 = (in_do&_net_3994);
   assign  _net_5200 = (in_do&_net_3994);
   assign  _net_5201 = (in_do&_net_3994);
   assign  _net_5202 = (in_do&_net_3994);
   assign  _net_5203 = (in_do&_net_3994);
   assign  _net_5204 = (in_do&_net_3994);
   assign  _net_5205 = (in_do&_net_3994);
   assign  _net_5206 = (in_do&_net_3994);
   assign  _net_5207 = (in_do&_net_3994);
   assign  _net_5208 = (in_do&_net_3994);
   assign  _net_5209 = (in_do&_net_3994);
   assign  _net_5210 = (in_do&_net_3994);
   assign  _net_5211 = (in_do&_net_3994);
   assign  _net_5212 = (in_do&_net_3994);
   assign  _net_5213 = (in_do&_net_3994);
   assign  _net_5214 = (in_do&_net_3994);
   assign  _net_5215 = (in_do&_net_3994);
   assign  _net_5216 = (in_do&_net_3994);
   assign  _net_5217 = (in_do&_net_3994);
   assign  _net_5218 = (in_do&_net_3994);
   assign  _net_5219 = (in_do&_net_3994);
   assign  _net_5220 = (in_do&_net_3994);
   assign  _net_5221 = (in_do&_net_3994);
   assign  _net_5222 = (in_do&_net_3994);
   assign  _net_5223 = (in_do&_net_3994);
   assign  _net_5224 = (in_do&_net_3994);
   assign  _net_5225 = (in_do&_net_3994);
   assign  _net_5226 = (in_do&_net_3994);
   assign  _net_5227 = (in_do&_net_3994);
   assign  _net_5228 = (in_do&_net_3994);
   assign  _net_5229 = (in_do&_net_3994);
   assign  _net_5230 = (in_do&_net_3994);
   assign  _net_5231 = (in_do&_net_3994);
   assign  _net_5232 = (in_do&_net_3994);
   assign  _net_5233 = (in_do&_net_3994);
   assign  _net_5234 = (in_do&_net_3994);
   assign  _net_5235 = (in_do&_net_3994);
   assign  _net_5236 = (in_do&_net_3994);
   assign  _net_5237 = (in_do&_net_3994);
   assign  _net_5238 = (in_do&_net_3994);
   assign  _net_5239 = (in_do&_net_3994);
   assign  _net_5240 = (in_do&_net_3994);
   assign  _net_5241 = (in_do&_net_3994);
   assign  _net_5242 = (in_do&_net_3994);
   assign  _net_5243 = (in_do&_net_3994);
   assign  _net_5244 = (in_do&_net_3994);
   assign  _net_5245 = (in_do&_net_3994);
   assign  _net_5246 = (in_do&_net_3994);
   assign  _net_5247 = (in_do&_net_3994);
   assign  _net_5248 = (in_do&_net_3994);
   assign  _net_5249 = (in_do&_net_3994);
   assign  _net_5250 = (in_do&_net_3994);
   assign  _net_5251 = (in_do&_net_3994);
   assign  _net_5252 = (in_do&_net_3994);
   assign  _net_5253 = (in_do&_net_3994);
   assign  _net_5254 = (in_do&_net_3994);
   assign  _net_5255 = (in_do&_net_3994);
   assign  _net_5256 = (in_do&_net_3994);
   assign  _net_5257 = (in_do&_net_3994);
   assign  _net_5258 = (in_do&_net_3994);
   assign  _net_5259 = (in_do&_net_3994);
   assign  _net_5260 = (in_do&_net_3994);
   assign  _net_5261 = (in_do&_net_3994);
   assign  _net_5262 = (in_do&_net_3994);
   assign  _net_5263 = (in_do&_net_3994);
   assign  _net_5264 = (in_do&_net_3994);
   assign  _net_5265 = (in_do&_net_3994);
   assign  _net_5266 = (in_do&_net_3994);
   assign  _net_5267 = (in_do&_net_3994);
   assign  _net_5268 = (in_do&_net_3994);
   assign  _net_5269 = (in_do&_net_3994);
   assign  _net_5270 = (in_do&_net_3994);
   assign  _net_5271 = (in_do&_net_3994);
   assign  _net_5272 = (in_do&_net_3994);
   assign  _net_5273 = (in_do&_net_3994);
   assign  _net_5274 = (in_do&_net_3994);
   assign  _net_5275 = (in_do&_net_3994);
   assign  _net_5276 = (in_do&_net_3994);
   assign  _net_5277 = (in_do&_net_3994);
   assign  _net_5278 = (in_do&_net_3994);
   assign  _net_5279 = (in_do&_net_3994);
   assign  _net_5280 = (in_do&_net_3994);
   assign  _net_5281 = (in_do&_net_3994);
   assign  _net_5282 = (in_do&_net_3994);
   assign  _net_5283 = (in_do&_net_3994);
   assign  _net_5284 = (in_do&_net_3994);
   assign  _net_5285 = (in_do&_net_3994);
   assign  _net_5286 = (in_do&_net_3994);
   assign  _net_5287 = (in_do&_net_3994);
   assign  _net_5288 = (in_do&_net_3994);
   assign  _net_5289 = (in_do&_net_3994);
   assign  _net_5290 = (in_do&_net_3994);
   assign  _net_5291 = (in_do&_net_3994);
   assign  _net_5292 = (in_do&_net_3994);
   assign  _net_5293 = (in_do&_net_3994);
   assign  _net_5294 = (in_do&_net_3994);
   assign  _net_5295 = (in_do&_net_3994);
   assign  _net_5296 = (in_do&_net_3994);
   assign  _net_5297 = (in_do&_net_3994);
   assign  _net_5298 = (in_do&_net_3994);
   assign  _net_5299 = (in_do&_net_3994);
   assign  _net_5300 = (in_do&_net_3994);
   assign  _net_5301 = (in_do&_net_3994);
   assign  _net_5302 = (in_do&_net_3994);
   assign  _net_5303 = (in_do&_net_3994);
   assign  _net_5304 = (in_do&_net_3994);
   assign  _net_5305 = (in_do&_net_3994);
   assign  _net_5306 = (in_do&_net_3994);
   assign  _net_5307 = (in_do&_net_3994);
   assign  _net_5308 = (in_do&_net_3994);
   assign  _net_5309 = (in_do&_net_3994);
   assign  _net_5310 = (in_do&_net_3994);
   assign  _net_5311 = (in_do&_net_3994);
   assign  _net_5312 = (in_do&_net_3994);
   assign  _net_5313 = (in_do&_net_3994);
   assign  _net_5314 = (in_do&_net_3994);
   assign  _net_5315 = (in_do&_net_3994);
   assign  _net_5316 = (in_do&_net_3994);
   assign  _net_5317 = (in_do&_net_3994);
   assign  _net_5318 = (in_do&_net_3994);
   assign  _net_5319 = (in_do&_net_3994);
   assign  _net_5320 = (in_do&_net_3994);
   assign  _net_5321 = (in_do&_net_3994);
   assign  _net_5322 = (in_do&_net_3994);
   assign  _net_5323 = (in_do&_net_3994);
   assign  _net_5324 = (in_do&_net_3994);
   assign  _net_5325 = (in_do&_net_3994);
   assign  _net_5326 = (in_do&_net_3994);
   assign  _net_5327 = (in_do&_net_3994);
   assign  _net_5328 = (in_do&_net_3994);
   assign  _net_5329 = (in_do&_net_3994);
   assign  _net_5330 = (in_do&_net_3994);
   assign  _net_5331 = (in_do&_net_3994);
   assign  _net_5332 = (in_do&_net_3994);
   assign  _net_5333 = (in_do&_net_3994);
   assign  _net_5334 = (in_do&_net_3994);
   assign  _net_5335 = (in_do&_net_3994);
   assign  _net_5336 = (in_do&_net_3994);
   assign  _net_5337 = (in_do&_net_3994);
   assign  _net_5338 = (in_do&_net_3994);
   assign  _net_5339 = (in_do&_net_3994);
   assign  _net_5340 = (in_do&_net_3994);
   assign  _net_5341 = (in_do&_net_3994);
   assign  _net_5342 = (in_do&_net_3994);
   assign  _net_5343 = (in_do&_net_3994);
   assign  _net_5344 = (in_do&_net_3994);
   assign  _net_5345 = (in_do&_net_3994);
   assign  _net_5346 = (in_do&_net_3994);
   assign  _net_5347 = (in_do&_net_3994);
   assign  _net_5348 = (in_do&_net_3994);
   assign  _net_5349 = (in_do&_net_3994);
   assign  _net_5350 = (in_do&_net_3994);
   assign  _net_5351 = (in_do&_net_3994);
   assign  _net_5352 = (in_do&_net_3994);
   assign  _net_5353 = (in_do&_net_3994);
   assign  _net_5354 = (in_do&_net_3994);
   assign  _net_5355 = (in_do&_net_3994);
   assign  _net_5356 = (in_do&_net_3994);
   assign  _net_5357 = (in_do&_net_3994);
   assign  _net_5358 = (in_do&_net_3994);
   assign  _net_5359 = (in_do&_net_3994);
   assign  _net_5360 = (in_do&_net_3994);
   assign  _net_5361 = (in_do&_net_3994);
   assign  _net_5362 = (in_do&_net_3994);
   assign  _net_5363 = (in_do&_net_3994);
   assign  _net_5364 = (in_do&_net_3994);
   assign  _net_5365 = (in_do&_net_3994);
   assign  _net_5366 = (in_do&_net_3994);
   assign  _net_5367 = (in_do&_net_3994);
   assign  _net_5368 = (in_do&_net_3994);
   assign  _net_5369 = (in_do&_net_3994);
   assign  _net_5370 = (in_do&_net_3994);
   assign  _net_5371 = (in_do&_net_3994);
   assign  _net_5372 = (in_do&_net_3994);
   assign  _net_5373 = (in_do&_net_3994);
   assign  _net_5374 = (in_do&_net_3994);
   assign  _net_5375 = (in_do&_net_3994);
   assign  _net_5376 = (in_do&_net_3994);
   assign  _net_5377 = (in_do&_net_3994);
   assign  _net_5378 = (in_do&_net_3994);
   assign  _net_5379 = (in_do&_net_3994);
   assign  _net_5380 = (in_do&_net_3994);
   assign  _net_5381 = (in_do&_net_3994);
   assign  _net_5382 = (in_do&_net_3994);
   assign  _net_5383 = (in_do&_net_3994);
   assign  _net_5384 = (in_do&_net_3994);
   assign  _net_5385 = (in_do&_net_3994);
   assign  _net_5386 = (in_do&_net_3994);
   assign  _net_5387 = (in_do&_net_3994);
   assign  _net_5388 = (in_do&_net_3994);
   assign  _net_5389 = (in_do&_net_3994);
   assign  _net_5390 = (in_do&_net_3994);
   assign  _net_5391 = (in_do&_net_3994);
   assign  _net_5392 = (in_do&_net_3994);
   assign  _net_5393 = (in_do&_net_3994);
   assign  _net_5394 = (in_do&_net_3994);
   assign  _net_5395 = (in_do&_net_3994);
   assign  _net_5396 = (in_do&_net_3994);
   assign  _net_5397 = (in_do&_net_3994);
   assign  _net_5398 = (in_do&_net_3994);
   assign  _net_5399 = (in_do&_net_3994);
   assign  _net_5400 = (in_do&_net_3994);
   assign  _net_5401 = (in_do&_net_3994);
   assign  _net_5402 = (in_do&_net_3994);
   assign  _net_5403 = (in_do&_net_3994);
   assign  _net_5404 = (in_do&_net_3994);
   assign  _net_5405 = (in_do&_net_3994);
   assign  _net_5406 = (in_do&_net_3994);
   assign  _net_5407 = (in_do&_net_3994);
   assign  _net_5408 = (in_do&_net_3994);
   assign  _net_5409 = (in_do&_net_3994);
   assign  _net_5410 = (in_do&_net_3994);
   assign  _net_5411 = (in_do&_net_3994);
   assign  _net_5412 = (in_do&_net_3994);
   assign  _net_5413 = (in_do&_net_3994);
   assign  _net_5414 = (in_do&_net_3994);
   assign  _net_5415 = (in_do&_net_3994);
   assign  _net_5416 = (in_do&_net_3994);
   assign  _net_5417 = (in_do&_net_3994);
   assign  _net_5418 = (in_do&_net_3994);
   assign  _net_5419 = (in_do&_net_3994);
   assign  _net_5420 = (in_do&_net_3994);
   assign  _net_5421 = (in_do&_net_3994);
   assign  _net_5422 = (in_do&_net_3994);
   assign  _net_5423 = (in_do&_net_3994);
   assign  _net_5424 = (in_do&_net_3994);
   assign  _net_5425 = (in_do&_net_3994);
   assign  _net_5426 = (in_do&_net_3994);
   assign  _net_5427 = (in_do&_net_3994);
   assign  _net_5428 = (in_do&_net_3994);
   assign  _net_5429 = (in_do&_net_3994);
   assign  _net_5430 = (in_do&_net_3994);
   assign  _net_5431 = (in_do&_net_3994);
   assign  _net_5432 = (in_do&_net_3994);
   assign  _net_5433 = (in_do&_net_3994);
   assign  _net_5434 = (in_do&_net_3994);
   assign  _net_5435 = (in_do&_net_3994);
   assign  _net_5436 = (in_do&_net_3994);
   assign  _net_5437 = (in_do&_net_3994);
   assign  _net_5438 = (in_do&_net_3994);
   assign  _net_5439 = (in_do&_net_3994);
   assign  _net_5440 = (in_do&_net_3994);
   assign  _net_5441 = (in_do&_net_3994);
   assign  _net_5442 = (in_do&_net_3994);
   assign  _net_5443 = (in_do&_net_3994);
   assign  _net_5444 = (in_do&_net_3994);
   assign  _net_5445 = (in_do&_net_3994);
   assign  _net_5446 = (in_do&_net_3994);
   assign  _net_5447 = (in_do&_net_3994);
   assign  _net_5448 = (in_do&_net_3994);
   assign  _net_5449 = (in_do&_net_3994);
   assign  _net_5450 = (in_do&_net_3994);
   assign  _net_5451 = (in_do&_net_3994);
   assign  _net_5452 = (in_do&_net_3994);
   assign  _net_5453 = (in_do&_net_3994);
   assign  _net_5454 = (in_do&_net_3994);
   assign  _net_5455 = (in_do&_net_3994);
   assign  _net_5456 = (in_do&_net_3994);
   assign  _net_5457 = (in_do&_net_3994);
   assign  _net_5458 = (in_do&_net_3994);
   assign  _net_5459 = (in_do&_net_3994);
   assign  _net_5460 = (in_do&_net_3994);
   assign  _net_5461 = (in_do&_net_3994);
   assign  _net_5462 = (in_do&_net_3994);
   assign  _net_5463 = (in_do&_net_3994);
   assign  _net_5464 = (in_do&_net_3994);
   assign  _net_5465 = (in_do&_net_3994);
   assign  _net_5466 = (in_do&_net_3994);
   assign  _net_5467 = (in_do&_net_3994);
   assign  _net_5468 = (in_do&_net_3994);
   assign  _net_5469 = (in_do&_net_3994);
   assign  _net_5470 = (in_do&_net_3994);
   assign  _net_5471 = (in_do&_net_3994);
   assign  _net_5472 = (in_do&_net_3994);
   assign  _net_5473 = (in_do&_net_3994);
   assign  _net_5474 = (in_do&_net_3994);
   assign  _net_5475 = (in_do&_net_3994);
   assign  _net_5476 = (in_do&_net_3994);
   assign  _net_5477 = (in_do&_net_3994);
   assign  _net_5478 = (in_do&_net_3994);
   assign  _net_5479 = (in_do&_net_3994);
   assign  _net_5480 = (in_do&_net_3994);
   assign  _net_5481 = (in_do&_net_3994);
   assign  _net_5482 = (in_do&_net_3994);
   assign  _net_5483 = (in_do&_net_3994);
   assign  _net_5484 = (in_do&_net_3994);
   assign  _net_5485 = (in_do&_net_3994);
   assign  _net_5486 = (in_do&_net_3994);
   assign  _net_5487 = (in_do&_net_3994);
   assign  _net_5488 = (in_do&_net_3994);
   assign  _net_5489 = (in_do&_net_3994);
   assign  _net_5490 = (in_do&_net_3994);
   assign  _net_5491 = (in_do&_net_3994);
   assign  _net_5492 = (in_do&_net_3994);
   assign  _net_5493 = (in_do&_net_3994);
   assign  _net_5494 = (in_do&_net_3994);
   assign  _net_5495 = (in_do&_net_3994);
   assign  _net_5496 = (in_do&_net_3994);
   assign  _net_5497 = (in_do&_net_3994);
   assign  _net_5498 = (in_do&_net_3994);
   assign  _net_5499 = (in_do&_net_3994);
   assign  _net_5500 = (in_do&_net_3994);
   assign  _net_5501 = (in_do&_net_3994);
   assign  _net_5502 = (in_do&_net_3994);
   assign  _net_5503 = (in_do&_net_3994);
   assign  _net_5504 = (in_do&_net_3994);
   assign  _net_5505 = (in_do&_net_3994);
   assign  _net_5506 = (in_do&_net_3994);
   assign  _net_5507 = (in_do&_net_3994);
   assign  _net_5508 = (in_do&_net_3994);
   assign  _net_5509 = (in_do&_net_3994);
   assign  _net_5510 = (in_do&_net_3994);
   assign  _net_5511 = (in_do&_net_3994);
   assign  _net_5512 = (in_do&_net_3994);
   assign  _net_5513 = (in_do&_net_3994);
   assign  _net_5514 = (in_do&_net_3994);
   assign  _net_5515 = (in_do&_net_3994);
   assign  _net_5516 = (in_do&_net_3994);
   assign  _net_5517 = (in_do&_net_3994);
   assign  _net_5518 = (in_do&_net_3994);
   assign  _net_5519 = (in_do&_net_3994);
   assign  _net_5520 = (in_do&_net_3994);
   assign  _net_5521 = (in_do&_net_3994);
   assign  _net_5522 = (in_do&_net_3994);
   assign  _net_5523 = (in_do&_net_3994);
   assign  _net_5524 = (in_do&_net_3994);
   assign  _net_5525 = (in_do&_net_3994);
   assign  _net_5526 = (in_do&_net_3994);
   assign  _net_5527 = (in_do&_net_3994);
   assign  _net_5528 = (in_do&_net_3994);
   assign  _net_5529 = (in_do&_net_3994);
   assign  _net_5530 = (in_do&_net_3994);
   assign  _net_5531 = (in_do&_net_3994);
   assign  _net_5532 = (in_do&_net_3994);
   assign  _net_5533 = (in_do&_net_3994);
   assign  _net_5534 = (in_do&_net_3994);
   assign  _net_5535 = (in_do&_net_3994);
   assign  _net_5536 = (in_do&_net_3994);
   assign  _net_5537 = (in_do&_net_3994);
   assign  _net_5538 = (in_do&_net_3994);
   assign  _net_5539 = (in_do&_net_3994);
   assign  _net_5540 = (in_do&_net_3994);
   assign  _net_5541 = (in_do&_net_3994);
   assign  _net_5542 = (in_do&_net_3994);
   assign  _net_5543 = (in_do&_net_3994);
   assign  _net_5544 = (in_do&_net_3994);
   assign  _net_5545 = (in_do&_net_3994);
   assign  _net_5546 = (in_do&_net_3994);
   assign  _net_5547 = (in_do&_net_3994);
   assign  _net_5548 = (in_do&_net_3994);
   assign  _net_5549 = (in_do&_net_3994);
   assign  _net_5550 = (in_do&_net_3994);
   assign  _net_5551 = (in_do&_net_3994);
   assign  _net_5552 = (in_do&_net_3994);
   assign  _net_5553 = (in_do&_net_3994);
   assign  _net_5554 = (in_do&_net_3994);
   assign  _net_5555 = (in_do&_net_3994);
   assign  _net_5556 = (in_do&_net_3994);
   assign  _net_5557 = (in_do&_net_3994);
   assign  _net_5558 = (in_do&_net_3994);
   assign  _net_5559 = (in_do&_net_3994);
   assign  _net_5560 = (in_do&_net_3994);
   assign  _net_5561 = (in_do&_net_3994);
   assign  _net_5562 = (in_do&_net_3994);
   assign  _net_5563 = (in_do&_net_3994);
   assign  _net_5564 = (in_do&_net_3994);
   assign  _net_5565 = (in_do&_net_3994);
   assign  _net_5566 = (in_do&_net_3994);
   assign  _net_5567 = (in_do&_net_3994);
   assign  _net_5568 = (in_do&_net_3994);
   assign  _net_5569 = (in_do&_net_3994);
   assign  _net_5570 = (in_do&_net_3994);
   assign  _net_5571 = (in_do&_net_3994);
   assign  _net_5572 = (in_do&_net_3994);
   assign  _net_5573 = (in_do&_net_3994);
   assign  _net_5574 = (in_do&_net_3994);
   assign  _net_5575 = (in_do&_net_3994);
   assign  _net_5576 = (in_do&_net_3994);
   assign  _net_5577 = (in_do&_net_3994);
   assign  _net_5578 = (in_do&_net_3994);
   assign  _net_5579 = (in_do&_net_3994);
   assign  _net_5580 = (in_do&_net_3994);
   assign  _net_5581 = (in_do&_net_3994);
   assign  _net_5582 = (in_do&_net_3994);
   assign  _net_5583 = (in_do&_net_3994);
   assign  _net_5584 = (in_do&_net_3994);
   assign  _net_5585 = (in_do&_net_3994);
   assign  _net_5586 = (in_do&_net_3994);
   assign  _net_5587 = (in_do&_net_3994);
   assign  _net_5588 = (in_do&_net_3994);
   assign  _net_5589 = (in_do&_net_3994);
   assign  _net_5590 = (in_do&_net_3994);
   assign  _net_5591 = (in_do&_net_3994);
   assign  _net_5592 = (in_do&_net_3994);
   assign  _net_5593 = (in_do&_net_3994);
   assign  _net_5594 = (in_do&_net_3994);
   assign  _net_5595 = (in_do&_net_3994);
   assign  _net_5596 = (in_do&_net_3994);
   assign  _net_5597 = (in_do&_net_3994);
   assign  _net_5598 = (in_do&_net_3994);
   assign  _net_5599 = (in_do&_net_3994);
   assign  _net_5600 = (in_do&_net_3994);
   assign  _net_5601 = (in_do&_net_3994);
   assign  _net_5602 = (in_do&_net_3994);
   assign  _net_5603 = (in_do&_net_3994);
   assign  _net_5604 = (in_do&_net_3994);
   assign  _net_5605 = (in_do&_net_3994);
   assign  _net_5606 = (in_do&_net_3994);
   assign  _net_5607 = (in_do&_net_3994);
   assign  _net_5608 = (in_do&_net_3994);
   assign  _net_5609 = (in_do&_net_3994);
   assign  _net_5610 = (in_do&_net_3994);
   assign  _net_5611 = (in_do&_net_3994);
   assign  _net_5612 = (in_do&_net_3994);
   assign  _net_5613 = (in_do&_net_3994);
   assign  _net_5614 = (in_do&_net_3994);
   assign  _net_5615 = (in_do&_net_3994);
   assign  _net_5616 = (in_do&_net_3994);
   assign  _net_5617 = (in_do&_net_3994);
   assign  _net_5618 = (in_do&_net_3994);
   assign  _net_5619 = (in_do&_net_3994);
   assign  _net_5620 = (in_do&_net_3994);
   assign  _net_5621 = (in_do&_net_3994);
   assign  _net_5622 = (in_do&_net_3994);
   assign  _net_5623 = (in_do&_net_3994);
   assign  _net_5624 = (in_do&_net_3994);
   assign  _net_5625 = (in_do&_net_3994);
   assign  _net_5626 = (in_do&_net_3994);
   assign  _net_5627 = (in_do&_net_3994);
   assign  _net_5628 = (in_do&_net_3994);
   assign  _net_5629 = (in_do&_net_3994);
   assign  _net_5630 = (in_do&_net_3994);
   assign  _net_5631 = (in_do&_net_3994);
   assign  _net_5632 = (in_do&_net_3994);
   assign  _net_5633 = (in_do&_net_3994);
   assign  _net_5634 = (in_do&_net_3994);
   assign  _net_5635 = (in_do&_net_3994);
   assign  _net_5636 = (in_do&_net_3994);
   assign  _net_5637 = (in_do&_net_3994);
   assign  _net_5638 = (in_do&_net_3994);
   assign  _net_5639 = (in_do&_net_3994);
   assign  _net_5640 = (in_do&_net_3994);
   assign  _net_5641 = (in_do&_net_3994);
   assign  _net_5642 = (in_do&_net_3994);
   assign  _net_5643 = (in_do&_net_3994);
   assign  _net_5644 = (in_do&_net_3994);
   assign  _net_5645 = (in_do&_net_3994);
   assign  _net_5646 = (in_do&_net_3994);
   assign  _net_5647 = (in_do&_net_3994);
   assign  _net_5648 = (in_do&_net_3994);
   assign  _net_5649 = (in_do&_net_3994);
   assign  _net_5650 = (in_do&_net_3994);
   assign  _net_5651 = (in_do&_net_3994);
   assign  _net_5652 = (in_do&_net_3994);
   assign  _net_5653 = (in_do&_net_3994);
   assign  _net_5654 = (in_do&_net_3994);
   assign  _net_5655 = (in_do&_net_3994);
   assign  _net_5656 = (in_do&_net_3994);
   assign  _net_5657 = (in_do&_net_3994);
   assign  _net_5658 = (in_do&_net_3994);
   assign  _net_5659 = (in_do&_net_3994);
   assign  _net_5660 = (in_do&_net_3994);
   assign  _net_5661 = (in_do&_net_3994);
   assign  _net_5662 = (in_do&_net_3994);
   assign  _net_5663 = (in_do&_net_3994);
   assign  _net_5664 = (in_do&_net_3994);
   assign  _net_5665 = (in_do&_net_3994);
   assign  _net_5666 = (in_do&_net_3994);
   assign  _net_5667 = (in_do&_net_3994);
   assign  _net_5668 = (in_do&_net_3994);
   assign  _net_5669 = (in_do&_net_3994);
   assign  _net_5670 = (in_do&_net_3994);
   assign  _net_5671 = (in_do&_net_3994);
   assign  _net_5672 = (in_do&_net_3994);
   assign  _net_5673 = (in_do&_net_3994);
   assign  _net_5674 = (in_do&_net_3994);
   assign  _net_5675 = (in_do&_net_3994);
   assign  _net_5676 = (in_do&_net_3994);
   assign  _net_5677 = (in_do&_net_3994);
   assign  _net_5678 = (in_do&_net_3994);
   assign  _net_5679 = (in_do&_net_3994);
   assign  _net_5680 = (in_do&_net_3994);
   assign  _net_5681 = (in_do&_net_3994);
   assign  _net_5682 = (in_do&_net_3994);
   assign  _net_5683 = (in_do&_net_3994);
   assign  _net_5684 = (in_do&_net_3994);
   assign  _net_5685 = (in_do&_net_3994);
   assign  _net_5686 = (in_do&_net_3994);
   assign  _net_5687 = (in_do&_net_3994);
   assign  _net_5688 = (in_do&_net_3994);
   assign  _net_5689 = (in_do&_net_3994);
   assign  _net_5690 = (in_do&_net_3994);
   assign  _net_5691 = (in_do&_net_3994);
   assign  _net_5692 = (in_do&_net_3994);
   assign  _net_5693 = (in_do&_net_3994);
   assign  _net_5694 = (in_do&_net_3994);
   assign  _net_5695 = (in_do&_net_3994);
   assign  _net_5696 = (in_do&_net_3994);
   assign  _net_5697 = (in_do&_net_3994);
   assign  _net_5698 = (in_do&_net_3994);
   assign  _net_5699 = (in_do&_net_3994);
   assign  _net_5700 = (in_do&_net_3994);
   assign  _net_5701 = (in_do&_net_3994);
   assign  _net_5702 = (in_do&_net_3994);
   assign  _net_5703 = (in_do&_net_3994);
   assign  _net_5704 = (in_do&_net_3994);
   assign  _net_5705 = (in_do&_net_3994);
   assign  _net_5706 = (in_do&_net_3994);
   assign  _net_5707 = (in_do&_net_3994);
   assign  _net_5708 = (in_do&_net_3994);
   assign  _net_5709 = (in_do&_net_3994);
   assign  _net_5710 = (in_do&_net_3994);
   assign  _net_5711 = (in_do&_net_3994);
   assign  _net_5712 = (in_do&_net_3994);
   assign  _net_5713 = (in_do&_net_3994);
   assign  _net_5714 = (in_do&_net_3994);
   assign  _net_5715 = (in_do&_net_3994);
   assign  _net_5716 = (in_do&_net_3994);
   assign  _net_5717 = (in_do&_net_3994);
   assign  _net_5718 = (in_do&_net_3994);
   assign  _net_5719 = (in_do&_net_3994);
   assign  _net_5720 = (in_do&_net_3994);
   assign  _net_5721 = (in_do&_net_3994);
   assign  _net_5722 = (in_do&_net_3994);
   assign  _net_5723 = (in_do&_net_3994);
   assign  _net_5724 = (in_do&_net_3994);
   assign  _net_5725 = (in_do&_net_3994);
   assign  _net_5726 = (in_do&_net_3994);
   assign  _net_5727 = (in_do&_net_3994);
   assign  _net_5728 = (in_do&_net_3994);
   assign  _net_5729 = (in_do&_net_3994);
   assign  _net_5730 = (in_do&_net_3994);
   assign  _net_5731 = (in_do&_net_3994);
   assign  _net_5732 = (in_do&_net_3994);
   assign  _net_5733 = (in_do&_net_3994);
   assign  _net_5734 = (in_do&_net_3994);
   assign  _net_5735 = (in_do&_net_3994);
   assign  _net_5736 = (in_do&_net_3994);
   assign  _net_5737 = (in_do&_net_3994);
   assign  _net_5738 = (in_do&_net_3994);
   assign  _net_5739 = (in_do&_net_3994);
   assign  _net_5740 = (in_do&_net_3994);
   assign  _net_5741 = (in_do&_net_3994);
   assign  _net_5742 = (in_do&_net_3994);
   assign  _net_5743 = (in_do&_net_3994);
   assign  _net_5744 = (in_do&_net_3994);
   assign  _net_5745 = (in_do&_net_3994);
   assign  _net_5746 = (in_do&_net_3994);
   assign  _net_5747 = (in_do&_net_3994);
   assign  _net_5748 = (in_do&_net_3994);
   assign  _net_5749 = (in_do&_net_3994);
   assign  _net_5750 = (in_do&_net_3994);
   assign  _net_5751 = (in_do&_net_3994);
   assign  _net_5752 = (in_do&_net_3994);
   assign  _net_5753 = (in_do&_net_3994);
   assign  _net_5754 = (in_do&_net_3994);
   assign  _net_5755 = (in_do&_net_3994);
   assign  _net_5756 = (in_do&_net_3994);
   assign  _net_5757 = (in_do&_net_3994);
   assign  _net_5758 = (in_do&_net_3994);
   assign  _net_5759 = (in_do&_net_3994);
   assign  _net_5760 = (in_do&_net_3994);
   assign  _net_5761 = (in_do&_net_3994);
   assign  _net_5762 = (in_do&_net_3994);
   assign  _net_5763 = (in_do&_net_3994);
   assign  _net_5764 = (in_do&_net_3994);
   assign  _net_5765 = (in_do&_net_3994);
   assign  _net_5766 = (in_do&_net_3994);
   assign  _net_5767 = (in_do&_net_3994);
   assign  _net_5768 = (in_do&_net_3994);
   assign  _net_5769 = (in_do&_net_3994);
   assign  _net_5770 = (in_do&_net_3994);
   assign  _net_5771 = (in_do&_net_3994);
   assign  _net_5772 = (in_do&_net_3994);
   assign  _net_5773 = (in_do&_net_3994);
   assign  _net_5774 = (in_do&_net_3994);
   assign  _net_5775 = (in_do&_net_3994);
   assign  _net_5776 = (in_do&_net_3994);
   assign  _net_5777 = (in_do&_net_3994);
   assign  _net_5778 = (in_do&_net_3994);
   assign  _net_5779 = (in_do&_net_3994);
   assign  _net_5780 = (in_do&_net_3994);
   assign  _net_5781 = (in_do&_net_3994);
   assign  _net_5782 = (in_do&_net_3994);
   assign  _net_5783 = (in_do&_net_3994);
   assign  _net_5784 = (in_do&_net_3994);
   assign  _net_5785 = (in_do&_net_3994);
   assign  _net_5786 = (in_do&_net_3994);
   assign  _net_5787 = (in_do&_net_3994);
   assign  _net_5788 = (in_do&_net_3994);
   assign  _net_5789 = (in_do&_net_3994);
   assign  _net_5790 = (in_do&_net_3994);
   assign  _net_5791 = (in_do&_net_3994);
   assign  _net_5792 = (in_do&_net_3994);
   assign  _net_5793 = (in_do&_net_3994);
   assign  _net_5794 = (in_do&_net_3994);
   assign  _net_5795 = (in_do&_net_3994);
   assign  _net_5796 = (in_do&_net_3994);
   assign  _net_5797 = (in_do&_net_3994);
   assign  _net_5798 = (in_do&_net_3994);
   assign  _net_5799 = (in_do&_net_3994);
   assign  _net_5800 = (in_do&_net_3994);
   assign  _net_5801 = (in_do&_net_3994);
   assign  _net_5802 = (in_do&_net_3994);
   assign  _net_5803 = (in_do&_net_3994);
   assign  _net_5804 = (in_do&_net_3994);
   assign  _net_5805 = (in_do&_net_3994);
   assign  _net_5806 = (in_do&_net_3994);
   assign  _net_5807 = (in_do&_net_3994);
   assign  _net_5808 = (in_do&_net_3994);
   assign  _net_5809 = (in_do&_net_3994);
   assign  _net_5810 = (in_do&_net_3994);
   assign  _net_5811 = (in_do&_net_3994);
   assign  _net_5812 = (in_do&_net_3994);
   assign  _net_5813 = (in_do&_net_3994);
   assign  _net_5814 = (in_do&_net_3994);
   assign  _net_5815 = (in_do&_net_3994);
   assign  _net_5816 = (in_do&_net_3994);
   assign  _net_5817 = (in_do&_net_3994);
   assign  _net_5818 = (in_do&_net_3994);
   assign  _net_5819 = (in_do&_net_3994);
   assign  _net_5820 = (in_do&_net_3994);
   assign  _net_5821 = (in_do&_net_3994);
   assign  _net_5822 = (in_do&_net_3994);
   assign  _net_5823 = (in_do&_net_3994);
   assign  _net_5824 = (in_do&_net_3994);
   assign  _net_5825 = (in_do&_net_3994);
   assign  _net_5826 = (in_do&_net_3994);
   assign  _net_5827 = (in_do&_net_3994);
   assign  _net_5828 = (in_do&_net_3994);
   assign  _net_5829 = (in_do&_net_3994);
   assign  _net_5830 = (in_do&_net_3994);
   assign  _net_5831 = (in_do&_net_3994);
   assign  _net_5832 = (in_do&_net_3994);
   assign  _net_5833 = (in_do&_net_3994);
   assign  _net_5834 = (in_do&_net_3994);
   assign  _net_5835 = (in_do&_net_3994);
   assign  _net_5836 = (in_do&_net_3994);
   assign  _net_5837 = (in_do&_net_3994);
   assign  _net_5838 = (in_do&_net_3994);
   assign  _net_5839 = (in_do&_net_3994);
   assign  _net_5840 = (in_do&_net_3994);
   assign  _net_5841 = (in_do&_net_3994);
   assign  _net_5842 = (in_do&_net_3994);
   assign  _net_5843 = (in_do&_net_3994);
   assign  _net_5844 = (in_do&_net_3994);
   assign  _net_5845 = (in_do&_net_3994);
   assign  _net_5846 = (in_do&_net_3994);
   assign  _net_5847 = (in_do&_net_3994);
   assign  _net_5848 = (in_do&_net_3994);
   assign  _net_5849 = (in_do&_net_3994);
   assign  _net_5850 = (in_do&_net_3994);
   assign  _net_5851 = (in_do&_net_3994);
   assign  _net_5852 = (in_do&_net_3994);
   assign  _net_5853 = (in_do&_net_3994);
   assign  _net_5854 = (in_do&_net_3994);
   assign  _net_5855 = (in_do&_net_3994);
   assign  _net_5856 = (in_do&_net_3994);
   assign  _net_5857 = (in_do&_net_3994);
   assign  _net_5858 = (in_do&_net_3994);
   assign  _net_5859 = (in_do&_net_3994);
   assign  _net_5860 = (in_do&_net_3994);
   assign  _net_5861 = (in_do&_net_3994);
   assign  _net_5862 = (in_do&_net_3994);
   assign  _net_5863 = (in_do&_net_3994);
   assign  _net_5864 = (in_do&_net_3994);
   assign  _net_5865 = (in_do&_net_3994);
   assign  _net_5866 = (in_do&_net_3994);
   assign  _net_5867 = (in_do&_net_3994);
   assign  _net_5868 = (in_do&_net_3994);
   assign  _net_5869 = (in_do&_net_3994);
   assign  _net_5870 = (in_do&_net_3994);
   assign  _net_5871 = (in_do&_net_3994);
   assign  _net_5872 = (in_do&_net_3994);
   assign  _net_5873 = (in_do&_net_3994);
   assign  _net_5874 = (in_do&_net_3994);
   assign  _net_5875 = (in_do&_net_3994);
   assign  _net_5876 = (in_do&_net_3994);
   assign  _net_5877 = (in_do&_net_3994);
   assign  _net_5878 = (in_do&_net_3994);
   assign  _net_5879 = (in_do&_net_3994);
   assign  _net_5880 = (in_do&_net_3994);
   assign  _net_5881 = (in_do&_net_3994);
   assign  _net_5882 = (in_do&_net_3994);
   assign  _net_5883 = (in_do&_net_3994);
   assign  _net_5884 = (in_do&_net_3994);
   assign  _net_5885 = (in_do&_net_3994);
   assign  _net_5886 = (in_do&_net_3994);
   assign  _net_5887 = (in_do&_net_3994);
   assign  _net_5888 = (in_do&_net_3994);
   assign  _net_5889 = (in_do&_net_3994);
   assign  _net_5890 = (in_do&_net_3994);
   assign  _net_5891 = (in_do&_net_3994);
   assign  _net_5892 = (in_do&_net_3994);
   assign  _net_5893 = (in_do&_net_3994);
   assign  _net_5894 = (in_do&_net_3994);
   assign  _net_5895 = (in_do&_net_3994);
   assign  _net_5896 = (in_do&_net_3994);
   assign  _net_5897 = (in_do&_net_3994);
   assign  _net_5898 = (in_do&_net_3994);
   assign  _net_5899 = (in_do&_net_3994);
   assign  _net_5900 = (in_do&_net_3994);
   assign  _net_5901 = (in_do&_net_3994);
   assign  _net_5902 = (in_do&_net_3994);
   assign  _net_5903 = (in_do&_net_3994);
   assign  _net_5904 = (in_do&_net_3994);
   assign  _net_5905 = (in_do&_net_3994);
   assign  _net_5906 = (in_do&_net_3994);
   assign  _net_5907 = (in_do&_net_3994);
   assign  _net_5908 = (in_do&_net_3994);
   assign  _net_5909 = (in_do&_net_3994);
   assign  _net_5910 = (in_do&_net_3994);
   assign  _net_5911 = (in_do&_net_3994);
   assign  _net_5912 = (in_do&_net_3994);
   assign  _net_5913 = (in_do&_net_3994);
   assign  _net_5914 = (in_do&_net_3994);
   assign  _net_5915 = (in_do&_net_3994);
   assign  _net_5916 = (in_do&_net_3994);
   assign  _net_5917 = (in_do&_net_3994);
   assign  _net_5918 = (in_do&_net_3994);
   assign  _net_5919 = (in_do&_net_3994);
   assign  _net_5920 = (in_do&_net_3994);
   assign  _net_5921 = (in_do&_net_3994);
   assign  _net_5922 = (in_do&_net_3994);
   assign  _net_5923 = (in_do&_net_3994);
   assign  _net_5924 = (in_do&_net_3994);
   assign  _net_5925 = (in_do&_net_3994);
   assign  _net_5926 = (in_do&_net_3994);
   assign  _net_5927 = (in_do&_net_3994);
   assign  _net_5928 = (in_do&_net_3994);
   assign  _net_5929 = (in_do&_net_3994);
   assign  _net_5930 = (in_do&_net_3994);
   assign  _net_5931 = (in_do&_net_3994);
   assign  _net_5932 = (in_do&_net_3994);
   assign  _net_5933 = (in_do&_net_3994);
   assign  _net_5934 = (in_do&_net_3994);
   assign  _net_5935 = (in_do&_net_3994);
   assign  _net_5936 = (in_do&_net_3994);
   assign  _net_5937 = (in_do&_net_3994);
   assign  _net_5938 = (in_do&_net_3994);
   assign  _net_5939 = (in_do&_net_3994);
   assign  _net_5940 = (in_do&_net_3994);
   assign  _net_5941 = (in_do&_net_3994);
   assign  _net_5942 = (in_do&_net_3994);
   assign  _net_5943 = (in_do&_net_3994);
   assign  _net_5944 = (in_do&_net_3994);
   assign  _net_5945 = (in_do&_net_3994);
   assign  _net_5946 = (in_do&_net_3994);
   assign  _net_5947 = (in_do&_net_3994);
   assign  _net_5948 = (in_do&_net_3994);
   assign  _net_5949 = (in_do&_net_3994);
   assign  _net_5950 = (in_do&_net_3994);
   assign  _net_5951 = (in_do&_net_3994);
   assign  _net_5952 = (in_do&_net_3994);
   assign  _net_5953 = (in_do&_net_3994);
   assign  _net_5954 = (in_do&_net_3994);
   assign  _net_5955 = (in_do&_net_3994);
   assign  _net_5956 = (in_do&_net_3994);
   assign  _net_5957 = (in_do&_net_3994);
   assign  _net_5958 = (in_do&_net_3994);
   assign  _net_5959 = (in_do&_net_3994);
   assign  _net_5960 = (in_do&_net_3994);
   assign  _net_5961 = (in_do&_net_3994);
   assign  _net_5962 = (in_do&_net_3994);
   assign  _net_5963 = (in_do&_net_3994);
   assign  _net_5964 = (in_do&_net_3994);
   assign  _net_5965 = (in_do&_net_3994);
   assign  _net_5966 = (in_do&_net_3994);
   assign  _net_5967 = (in_do&_net_3994);
   assign  _net_5968 = (in_do&_net_3994);
   assign  _net_5969 = (in_do&_net_3994);
   assign  _net_5970 = (in_do&_net_3994);
   assign  _net_5971 = (in_do&_net_3994);
   assign  _net_5972 = (in_do&_net_3994);
   assign  _net_5973 = (in_do&_net_3994);
   assign  _net_5974 = (in_do&_net_3994);
   assign  _net_5975 = (in_do&_net_3994);
   assign  _net_5976 = (in_do&_net_3994);
   assign  _net_5977 = (in_do&_net_3994);
   assign  _net_5978 = (in_do&_net_3994);
   assign  _net_5979 = (in_do&_net_3994);
   assign  _net_5980 = (in_do&_net_3994);
   assign  _net_5981 = (in_do&_net_3994);
   assign  _net_5982 = (in_do&_net_3994);
   assign  _net_5983 = (in_do&_net_3994);
   assign  _net_5984 = (in_do&_net_3994);
   assign  _net_5985 = (in_do&_net_3994);
   assign  _net_5986 = (in_do&_net_3994);
   assign  _net_5987 = (in_do&_net_3994);
   assign  _net_5988 = (in_do&_net_3994);
   assign  _net_5989 = (in_do&_net_3994);
   assign  _net_5990 = (in_do&_net_3994);
   assign  _net_5991 = (in_do&_net_3994);
   assign  _net_5992 = (in_do&_net_3994);
   assign  _net_5993 = (in_do&_net_3994);
   assign  _net_5994 = (in_do&_net_3994);
   assign  _net_5995 = (in_do&_net_3994);
   assign  _net_5996 = (in_do&_net_3994);
   assign  _net_5997 = (in_do&_net_3994);
   assign  _net_5998 = (in_do&_net_3994);
   assign  _net_5999 = (in_do&_net_3994);
   assign  _net_6000 = (in_do&_net_3994);
   assign  _net_6001 = (in_do&_net_3994);
   assign  _net_6002 = (in_do&_net_3994);
   assign  _net_6003 = (in_do&_net_3994);
   assign  _net_6004 = (in_do&_net_3994);
   assign  _net_6005 = (in_do&_net_3994);
   assign  _net_6006 = (in_do&_net_3994);
   assign  _net_6007 = (in_do&_net_3994);
   assign  _net_6008 = (in_do&_net_3994);
   assign  _net_6009 = (in_do&_net_3994);
   assign  _net_6010 = (in_do&_net_3994);
   assign  _net_6011 = (in_do&_net_3994);
   assign  _net_6012 = (in_do&_net_3994);
   assign  _net_6013 = (in_do&_net_3994);
   assign  _net_6014 = (in_do&_net_3994);
   assign  _net_6015 = (in_do&_net_3994);
   assign  _net_6016 = (in_do&_net_3994);
   assign  _net_6017 = (in_do&_net_3994);
   assign  _net_6018 = (in_do&_net_3994);
   assign  _net_6019 = (in_do&_net_3994);
   assign  _net_6020 = (in_do&_net_3994);
   assign  _net_6021 = (in_do&_net_3994);
   assign  _net_6022 = (in_do&_net_3994);
   assign  _net_6023 = (in_do&_net_3994);
   assign  _net_6024 = (in_do&_net_3994);
   assign  _net_6025 = (in_do&_net_3994);
   assign  _net_6026 = (in_do&_net_3994);
   assign  _net_6027 = (in_do&_net_3994);
   assign  _net_6028 = (in_do&_net_3994);
   assign  _net_6029 = (in_do&_net_3994);
   assign  _net_6030 = (in_do&_net_3994);
   assign  _net_6031 = (in_do&_net_3994);
   assign  _net_6032 = (in_do&_net_3994);
   assign  _net_6033 = (in_do&_net_3994);
   assign  _net_6034 = (in_do&_net_3994);
   assign  _net_6035 = (in_do&_net_3994);
   assign  _net_6036 = (in_do&_net_3994);
   assign  _net_6037 = (in_do&_net_3994);
   assign  _net_6038 = (in_do&_net_3994);
   assign  _net_6039 = (in_do&_net_3994);
   assign  _net_6040 = (in_do&_net_3994);
   assign  _net_6041 = (in_do&_net_3994);
   assign  _net_6042 = (in_do&_net_3994);
   assign  _net_6043 = (in_do&_net_3994);
   assign  _net_6044 = (in_do&_net_3994);
   assign  _net_6045 = (in_do&_net_3994);
   assign  _net_6046 = (in_do&_net_3994);
   assign  _net_6047 = (in_do&_net_3994);
   assign  _net_6048 = (in_do&_net_3994);
   assign  _net_6049 = (in_do&_net_3994);
   assign  _net_6050 = (in_do&_net_3994);
   assign  _net_6051 = (in_do&_net_3994);
   assign  _net_6052 = (in_do&_net_3994);
   assign  _net_6053 = (in_do&_net_3994);
   assign  _net_6054 = (in_do&_net_3994);
   assign  _net_6055 = (in_do&_net_3994);
   assign  _net_6056 = (in_do&_net_3994);
   assign  _net_6057 = (in_do&_net_3994);
   assign  _net_6058 = (in_do&_net_3994);
   assign  _net_6059 = (in_do&_net_3994);
   assign  _net_6060 = (in_do&_net_3994);
   assign  _net_6061 = (in_do&_net_3994);
   assign  _net_6062 = (in_do&_net_3994);
   assign  _net_6063 = (in_do&_net_3994);
   assign  _net_6064 = (in_do&_net_3994);
   assign  _net_6065 = (in_do&_net_3994);
   assign  _net_6066 = (in_do&_net_3994);
   assign  _net_6067 = (in_do&_net_3994);
   assign  _net_6068 = (in_do&_net_3994);
   assign  _net_6069 = (in_do&_net_3994);
   assign  _net_6070 = (in_do&_net_3994);
   assign  _net_6071 = (in_do&_net_3994);
   assign  _net_6072 = (in_do&_net_3994);
   assign  _net_6073 = (in_do&_net_3994);
   assign  _net_6074 = (in_do&_net_3994);
   assign  _net_6075 = (in_do&_net_3994);
   assign  _net_6076 = (in_do&_net_3994);
   assign  _net_6077 = (in_do&_net_3994);
   assign  _net_6078 = (in_do&_net_3994);
   assign  _net_6079 = (in_do&_net_3994);
   assign  _net_6080 = (in_do&_net_3994);
   assign  _net_6081 = (in_do&_net_3994);
   assign  _net_6082 = (in_do&_net_3994);
   assign  _net_6083 = (in_do&_net_3994);
   assign  _net_6084 = (in_do&_net_3994);
   assign  _net_6085 = (in_do&_net_3994);
   assign  _net_6086 = (in_do&_net_3994);
   assign  _net_6087 = (in_do&_net_3994);
   assign  _net_6088 = (in_do&_net_3994);
   assign  _net_6089 = (in_do&_net_3994);
   assign  _net_6090 = (in_do&_net_3994);
   assign  _net_6091 = (in_do&_net_3994);
   assign  _net_6092 = (in_do&_net_3994);
   assign  _net_6093 = (in_do&_net_3994);
   assign  _net_6094 = (in_do&_net_3994);
   assign  _net_6095 = (in_do&_net_3994);
   assign  _net_6096 = (in_do&_net_3994);
   assign  _net_6097 = (in_do&_net_3994);
   assign  _net_6098 = (in_do&_net_3994);
   assign  _net_6099 = (in_do&_net_3994);
   assign  _net_6100 = (in_do&_net_3994);
   assign  _net_6101 = (in_do&_net_3994);
   assign  _net_6102 = (in_do&_net_3994);
   assign  _net_6103 = (in_do&_net_3994);
   assign  _net_6104 = (in_do&_net_3994);
   assign  _net_6105 = (in_do&_net_3994);
   assign  _net_6106 = (in_do&_net_3994);
   assign  _net_6107 = (in_do&_net_3994);
   assign  _net_6108 = (in_do&_net_3994);
   assign  _net_6109 = (in_do&_net_3994);
   assign  _net_6110 = (in_do&_net_3994);
   assign  _net_6111 = (in_do&_net_3994);
   assign  _net_6112 = (in_do&_net_3994);
   assign  _net_6113 = (in_do&_net_3994);
   assign  _net_6114 = (in_do&_net_3994);
   assign  _net_6115 = (in_do&_net_3994);
   assign  _net_6116 = (in_do&_net_3994);
   assign  _net_6117 = (in_do&_net_3994);
   assign  _net_6118 = (in_do&_net_3994);
   assign  _net_6119 = (in_do&_net_3994);
   assign  _net_6120 = (in_do&_net_3994);
   assign  _net_6121 = (in_do&_net_3994);
   assign  _net_6122 = (in_do&_net_3994);
   assign  _net_6123 = (in_do&_net_3994);
   assign  _net_6124 = (in_do&_net_3994);
   assign  _net_6125 = (in_do&_net_3994);
   assign  _net_6126 = (in_do&_net_3994);
   assign  _net_6127 = (in_do&_net_3994);
   assign  _net_6128 = (in_do&_net_3994);
   assign  _net_6129 = (in_do&_net_3994);
   assign  _net_6130 = (in_do&_net_3994);
   assign  _net_6131 = (in_do&_net_3994);
   assign  _net_6132 = (in_do&_net_3994);
   assign  _net_6133 = (in_do&_net_3994);
   assign  _net_6134 = (in_do&_net_3994);
   assign  _net_6135 = (in_do&_net_3994);
   assign  _net_6136 = (in_do&_net_3994);
   assign  _net_6137 = (in_do&_net_3994);
   assign  _net_6138 = (in_do&_net_3994);
   assign  _net_6139 = (in_do&_net_3994);
   assign  _net_6140 = (in_do&_net_3994);
   assign  _net_6141 = (in_do&_net_3994);
   assign  _net_6142 = (in_do&_net_3994);
   assign  _net_6143 = (in_do&_net_3994);
   assign  _net_6144 = (in_do&_net_3994);
   assign  _net_6145 = (in_do&_net_3994);
   assign  _net_6146 = (in_do&_net_3994);
   assign  _net_6147 = (in_do&_net_3994);
   assign  _net_6148 = (in_do&_net_3994);
   assign  _net_6149 = (in_do&_net_3994);
   assign  _net_6150 = (in_do&_net_3994);
   assign  _net_6151 = (in_do&_net_3994);
   assign  _net_6152 = (in_do&_net_3994);
   assign  _net_6153 = (in_do&_net_3994);
   assign  _net_6154 = (in_do&_net_3994);
   assign  _net_6155 = (in_do&_net_3994);
   assign  _net_6156 = (in_do&_net_3994);
   assign  _net_6157 = (in_do&_net_3994);
   assign  _net_6158 = (in_do&_net_3994);
   assign  _net_6159 = (in_do&_net_3994);
   assign  _net_6160 = (in_do&_net_3994);
   assign  _net_6161 = (in_do&_net_3994);
   assign  _net_6162 = (in_do&_net_3994);
   assign  _net_6163 = (in_do&_net_3994);
   assign  _net_6164 = (in_do&_net_3994);
   assign  _net_6165 = (in_do&_net_3994);
   assign  _net_6166 = (in_do&_net_3994);
   assign  _net_6167 = (in_do&_net_3994);
   assign  _net_6168 = (in_do&_net_3994);
   assign  _net_6169 = (in_do&_net_3994);
   assign  _net_6170 = (in_do&_net_3994);
   assign  _net_6171 = (in_do&_net_3994);
   assign  _net_6172 = (in_do&_net_3994);
   assign  _net_6173 = (in_do&_net_3994);
   assign  _net_6174 = (in_do&_net_3994);
   assign  _net_6175 = (in_do&_net_3994);
   assign  _net_6176 = (in_do&_net_3994);
   assign  _net_6177 = (in_do&_net_3994);
   assign  _net_6178 = (in_do&_net_3994);
   assign  _net_6179 = (in_do&_net_3994);
   assign  _net_6180 = (in_do&_net_3994);
   assign  _net_6181 = (in_do&_net_3994);
   assign  _net_6182 = (in_do&_net_3994);
   assign  _net_6183 = (in_do&_net_3994);
   assign  _net_6184 = (in_do&_net_3994);
   assign  _net_6185 = (in_do&_net_3994);
   assign  _net_6186 = (in_do&_net_3994);
   assign  _net_6187 = (in_do&_net_3994);
   assign  _net_6188 = (in_do&_net_3994);
   assign  _net_6189 = (in_do&_net_3994);
   assign  _net_6190 = (in_do&_net_3994);
   assign  _net_6191 = (in_do&_net_3994);
   assign  _net_6192 = (in_do&_net_3994);
   assign  _net_6193 = (in_do&_net_3994);
   assign  _net_6194 = (in_do&_net_3994);
   assign  _net_6195 = (in_do&_net_3994);
   assign  _net_6196 = (in_do&_net_3994);
   assign  _net_6197 = (in_do&_net_3994);
   assign  _net_6198 = (in_do&_net_3994);
   assign  _net_6199 = (in_do&_net_3994);
   assign  _net_6200 = (in_do&_net_3994);
   assign  _net_6201 = (in_do&_net_3994);
   assign  _net_6202 = (in_do&_net_3994);
   assign  _net_6203 = (in_do&_net_3994);
   assign  _net_6204 = (in_do&_net_3994);
   assign  _net_6205 = (in_do&_net_3994);
   assign  _net_6206 = (in_do&_net_3994);
   assign  _net_6207 = (in_do&_net_3994);
   assign  _net_6208 = (in_do&_net_3994);
   assign  _net_6209 = (in_do&_net_3994);
   assign  _net_6210 = (in_do&_net_3994);
   assign  _net_6211 = (in_do&_net_3994);
   assign  _net_6212 = (in_do&_net_3994);
   assign  _net_6213 = (in_do&_net_3994);
   assign  _net_6214 = (in_do&_net_3994);
   assign  _net_6215 = (in_do&_net_3994);
   assign  _net_6216 = (in_do&_net_3994);
   assign  _net_6217 = (in_do&_net_3994);
   assign  _net_6218 = (in_do&_net_3994);
   assign  _net_6219 = (in_do&_net_3994);
   assign  _net_6220 = (in_do&_net_3994);
   assign  _net_6221 = (in_do&_net_3994);
   assign  _net_6222 = (in_do&_net_3994);
   assign  _net_6223 = (in_do&_net_3994);
   assign  _net_6224 = (in_do&_net_3994);
   assign  _net_6225 = (in_do&_net_3994);
   assign  _net_6226 = (in_do&_net_3994);
   assign  _net_6227 = (in_do&_net_3994);
   assign  _net_6228 = (in_do&_net_3994);
   assign  _net_6229 = (in_do&_net_3994);
   assign  _net_6230 = (in_do&_net_3994);
   assign  _net_6231 = (in_do&_net_3994);
   assign  _net_6232 = (in_do&_net_3994);
   assign  _net_6233 = (in_do&_net_3994);
   assign  _net_6234 = (in_do&_net_3994);
   assign  _net_6235 = (in_do&_net_3994);
   assign  _net_6236 = (in_do&_net_3994);
   assign  _net_6237 = (in_do&_net_3994);
   assign  _net_6238 = (in_do&_net_3994);
   assign  _net_6239 = (in_do&_net_3994);
   assign  _net_6240 = (in_do&_net_3994);
   assign  _net_6241 = (in_do&_net_3994);
   assign  _net_6242 = (in_do&_net_3994);
   assign  _net_6243 = (in_do&_net_3994);
   assign  _net_6244 = (in_do&_net_3994);
   assign  _net_6245 = (in_do&_net_3994);
   assign  _net_6246 = (in_do&_net_3994);
   assign  _net_6247 = (in_do&_net_3994);
   assign  _net_6248 = (in_do&_net_3994);
   assign  _net_6249 = (in_do&_net_3994);
   assign  _net_6250 = (in_do&_net_3994);
   assign  _net_6251 = (in_do&_net_3994);
   assign  _net_6252 = (in_do&_net_3994);
   assign  _net_6253 = (in_do&_net_3994);
   assign  _net_6254 = (in_do&_net_3994);
   assign  _net_6255 = (in_do&_net_3994);
   assign  _net_6256 = (in_do&_net_3994);
   assign  _net_6257 = (in_do&_net_3994);
   assign  _net_6258 = (in_do&_net_3994);
   assign  _net_6259 = (in_do&_net_3994);
   assign  _net_6260 = (in_do&_net_3994);
   assign  _net_6261 = (in_do&_net_3994);
   assign  _net_6262 = (in_do&_net_3994);
   assign  _net_6263 = (in_do&_net_3994);
   assign  _net_6264 = (in_do&_net_3994);
   assign  _net_6265 = (in_do&_net_3994);
   assign  _net_6266 = (in_do&_net_3994);
   assign  _net_6267 = (in_do&_net_3994);
   assign  _net_6268 = (in_do&_net_3994);
   assign  _net_6269 = (in_do&_net_3994);
   assign  _net_6270 = (in_do&_net_3994);
   assign  _net_6271 = (in_do&_net_3994);
   assign  _net_6272 = (in_do&_net_3994);
   assign  _net_6273 = (in_do&_net_3994);
   assign  _net_6274 = (in_do&_net_3994);
   assign  _net_6275 = (in_do&_net_3994);
   assign  _net_6276 = (in_do&_net_3994);
   assign  _net_6277 = (in_do&_net_3994);
   assign  _net_6278 = (in_do&_net_3994);
   assign  _net_6279 = (in_do&_net_3994);
   assign  _net_6280 = (in_do&_net_3994);
   assign  _net_6281 = (in_do&_net_3994);
   assign  _net_6282 = (in_do&_net_3994);
   assign  _net_6283 = (in_do&_net_3994);
   assign  _net_6284 = (in_do&_net_3994);
   assign  _net_6285 = (in_do&_net_3994);
   assign  _net_6286 = (in_do&_net_3994);
   assign  _net_6287 = (in_do&_net_3994);
   assign  _net_6288 = (in_do&_net_3994);
   assign  _net_6289 = (in_do&_net_3994);
   assign  _net_6290 = (in_do&_net_3994);
   assign  _net_6291 = (in_do&_net_3994);
   assign  _net_6292 = (in_do&_net_3994);
   assign  _net_6293 = (in_do&_net_3994);
   assign  _net_6294 = (in_do&_net_3994);
   assign  _net_6295 = (in_do&_net_3994);
   assign  _net_6296 = (in_do&_net_3994);
   assign  _net_6297 = (in_do&_net_3994);
   assign  _net_6298 = (in_do&_net_3994);
   assign  _net_6299 = (in_do&_net_3994);
   assign  _net_6300 = (in_do&_net_3994);
   assign  _net_6301 = (in_do&_net_3994);
   assign  _net_6302 = (in_do&_net_3994);
   assign  _net_6303 = (in_do&_net_3994);
   assign  _net_6304 = (in_do&_net_3994);
   assign  _net_6305 = (in_do&_net_3994);
   assign  _net_6306 = (in_do&_net_3994);
   assign  _net_6307 = (in_do&_net_3994);
   assign  _net_6308 = (in_do&_net_3994);
   assign  _net_6309 = (in_do&_net_3994);
   assign  _net_6310 = (in_do&_net_3994);
   assign  _net_6311 = (in_do&_net_3994);
   assign  _net_6312 = (in_do&_net_3994);
   assign  _net_6313 = (in_do&_net_3994);
   assign  _net_6314 = (in_do&_net_3994);
   assign  _net_6315 = (in_do&_net_3994);
   assign  _net_6316 = (in_do&_net_3994);
   assign  _net_6317 = (in_do&_net_3994);
   assign  _net_6318 = (in_do&_net_3994);
   assign  _net_6319 = (in_do&_net_3994);
   assign  _net_6320 = (in_do&_net_3994);
   assign  _net_6321 = (in_do&_net_3994);
   assign  _net_6322 = (in_do&_net_3994);
   assign  _net_6323 = (in_do&_net_3994);
   assign  _net_6324 = (in_do&_net_3994);
   assign  _net_6325 = (in_do&_net_3994);
   assign  _net_6326 = (in_do&_net_3994);
   assign  _net_6327 = (in_do&_net_3994);
   assign  _net_6328 = (in_do&_net_3994);
   assign  _net_6329 = (in_do&_net_3994);
   assign  _net_6330 = (in_do&_net_3994);
   assign  _net_6331 = (in_do&_net_3994);
   assign  _net_6332 = (in_do&_net_3994);
   assign  _net_6333 = (in_do&_net_3994);
   assign  _net_6334 = (in_do&_net_3994);
   assign  _net_6335 = (in_do&_net_3994);
   assign  _net_6336 = (in_do&_net_3994);
   assign  _net_6337 = (in_do&_net_3994);
   assign  _net_6338 = (in_do&_net_3994);
   assign  _net_6339 = (in_do&_net_3994);
   assign  _net_6340 = (in_do&_net_3994);
   assign  _net_6341 = (in_do&_net_3994);
   assign  _net_6342 = (in_do&_net_3994);
   assign  _net_6343 = (in_do&_net_3994);
   assign  _net_6344 = (in_do&_net_3994);
   assign  _net_6345 = (in_do&_net_3994);
   assign  _net_6346 = (in_do&_net_3994);
   assign  _net_6347 = (in_do&_net_3994);
   assign  _net_6348 = (in_do&_net_3994);
   assign  _net_6349 = (in_do&_net_3994);
   assign  _net_6350 = (in_do&_net_3994);
   assign  _net_6351 = (in_do&_net_3994);
   assign  _net_6352 = (in_do&_net_3994);
   assign  _net_6353 = (in_do&_net_3994);
   assign  _net_6354 = (in_do&_net_3994);
   assign  _net_6355 = (in_do&_net_3994);
   assign  _net_6356 = (in_do&_net_3994);
   assign  _net_6357 = (in_do&_net_3994);
   assign  _net_6358 = (in_do&_net_3994);
   assign  _net_6359 = (in_do&_net_3994);
   assign  _net_6360 = (in_do&_net_3994);
   assign  _net_6361 = (in_do&_net_3994);
   assign  _net_6362 = (in_do&_net_3994);
   assign  _net_6363 = (in_do&_net_3994);
   assign  _net_6364 = (in_do&_net_3994);
   assign  _net_6365 = (in_do&_net_3994);
   assign  _net_6366 = (in_do&_net_3994);
   assign  _net_6367 = (in_do&_net_3994);
   assign  _net_6368 = (in_do&_net_3994);
   assign  _net_6369 = (in_do&_net_3994);
   assign  _net_6370 = (in_do&_net_3994);
   assign  _net_6371 = (in_do&_net_3994);
   assign  _net_6372 = (in_do&_net_3994);
   assign  _net_6373 = (in_do&_net_3994);
   assign  _net_6374 = (in_do&_net_3994);
   assign  _net_6375 = (in_do&_net_3994);
   assign  _net_6376 = (in_do&_net_3994);
   assign  _net_6377 = (in_do&_net_3994);
   assign  _net_6378 = (in_do&_net_3994);
   assign  _net_6379 = (in_do&_net_3994);
   assign  _net_6380 = (in_do&_net_3994);
   assign  _net_6381 = (in_do&_net_3994);
   assign  _net_6382 = (in_do&_net_3994);
   assign  _net_6383 = (in_do&_net_3994);
   assign  _net_6384 = (in_do&_net_3994);
   assign  _net_6385 = (in_do&_net_3994);
   assign  _net_6386 = (in_do&_net_3994);
   assign  _net_6387 = (in_do&_net_3994);
   assign  _net_6388 = (in_do&_net_3994);
   assign  _net_6389 = (in_do&_net_3994);
   assign  _net_6390 = (in_do&_net_3994);
   assign  _net_6391 = (in_do&_net_3994);
   assign  _net_6392 = (in_do&_net_3994);
   assign  _net_6393 = (in_do&_net_3994);
   assign  _net_6394 = (in_do&_net_3994);
   assign  _net_6395 = (in_do&_net_3994);
   assign  _net_6396 = (in_do&_net_3994);
   assign  _net_6397 = (in_do&_net_3994);
   assign  _net_6398 = (in_do&_net_3994);
   assign  _net_6399 = (in_do&_net_3994);
   assign  _net_6400 = (in_do&_net_3994);
   assign  _net_6401 = (in_do&_net_3994);
   assign  _net_6402 = (in_do&_net_3994);
   assign  _net_6403 = (in_do&_net_3994);
   assign  _net_6404 = (in_do&_net_3994);
   assign  _net_6405 = (in_do&_net_3994);
   assign  _net_6406 = (in_do&_net_3994);
   assign  _net_6407 = (in_do&_net_3994);
   assign  _net_6408 = (in_do&_net_3994);
   assign  _net_6409 = (in_do&_net_3994);
   assign  _net_6410 = (in_do&_net_3994);
   assign  _net_6411 = (in_do&_net_3994);
   assign  _net_6412 = (in_do&_net_3994);
   assign  _net_6413 = (in_do&_net_3994);
   assign  _net_6414 = (in_do&_net_3994);
   assign  _net_6415 = (in_do&_net_3994);
   assign  _net_6416 = (in_do&_net_3994);
   assign  _net_6417 = (in_do&_net_3994);
   assign  _net_6418 = (in_do&_net_3994);
   assign  _net_6419 = (in_do&_net_3994);
   assign  _net_6420 = (in_do&_net_3994);
   assign  _net_6421 = (in_do&_net_3994);
   assign  _net_6422 = (in_do&_net_3994);
   assign  _net_6423 = (in_do&_net_3994);
   assign  _net_6424 = (in_do&_net_3994);
   assign  _net_6425 = (in_do&_net_3994);
   assign  _net_6426 = (in_do&_net_3994);
   assign  _net_6427 = (in_do&_net_3994);
   assign  _net_6428 = (in_do&_net_3994);
   assign  _net_6429 = (in_do&_net_3994);
   assign  _net_6430 = (in_do&_net_3994);
   assign  _net_6431 = (in_do&_net_3994);
   assign  _net_6432 = (in_do&_net_3994);
   assign  _net_6433 = (in_do&_net_3994);
   assign  _net_6434 = (in_do&_net_3994);
   assign  _net_6435 = (in_do&_net_3994);
   assign  _net_6436 = (in_do&_net_3994);
   assign  _net_6437 = (in_do&_net_3994);
   assign  _net_6438 = (in_do&_net_3994);
   assign  _net_6439 = (in_do&_net_3994);
   assign  _net_6440 = (in_do&_net_3994);
   assign  _net_6441 = (in_do&_net_3994);
   assign  _net_6442 = (in_do&_net_3994);
   assign  _net_6443 = (in_do&_net_3994);
   assign  _net_6444 = (in_do&_net_3994);
   assign  _net_6445 = (in_do&_net_3994);
   assign  _net_6446 = (in_do&_net_3994);
   assign  _net_6447 = (in_do&_net_3994);
   assign  _net_6448 = (in_do&_net_3994);
   assign  _net_6449 = (in_do&_net_3994);
   assign  _net_6450 = (in_do&_net_3994);
   assign  _net_6451 = (in_do&_net_3994);
   assign  _net_6452 = (in_do&_net_3994);
   assign  _net_6453 = (in_do&_net_3994);
   assign  _net_6454 = (in_do&_net_3994);
   assign  _net_6455 = (in_do&_net_3994);
   assign  _net_6456 = (in_do&_net_3994);
   assign  _net_6457 = (in_do&_net_3994);
   assign  _net_6458 = (in_do&_net_3994);
   assign  _net_6459 = (in_do&_net_3994);
   assign  _net_6460 = (in_do&_net_3994);
   assign  _net_6461 = (in_do&_net_3994);
   assign  _net_6462 = (in_do&_net_3994);
   assign  _net_6463 = (in_do&_net_3994);
   assign  _net_6464 = (in_do&_net_3994);
   assign  _net_6465 = (in_do&_net_3994);
   assign  _net_6466 = (in_do&_net_3994);
   assign  _net_6467 = (in_do&_net_3994);
   assign  _net_6468 = (in_do&_net_3994);
   assign  _net_6469 = (in_do&_net_3994);
   assign  _net_6470 = (in_do&_net_3994);
   assign  _net_6471 = (in_do&_net_3994);
   assign  _net_6472 = (in_do&_net_3994);
   assign  _net_6473 = (in_do&_net_3994);
   assign  _net_6474 = (in_do&_net_3994);
   assign  _net_6475 = (in_do&_net_3994);
   assign  _net_6476 = (in_do&_net_3994);
   assign  _net_6477 = (in_do&_net_3994);
   assign  _net_6478 = (in_do&_net_3994);
   assign  _net_6479 = (in_do&_net_3994);
   assign  _net_6480 = (in_do&_net_3994);
   assign  _net_6481 = (in_do&_net_3994);
   assign  _net_6482 = (in_do&_net_3994);
   assign  _net_6483 = (in_do&_net_3994);
   assign  _net_6484 = (in_do&_net_3994);
   assign  _net_6485 = (in_do&_net_3994);
   assign  _net_6486 = (in_do&_net_3994);
   assign  _net_6487 = (in_do&_net_3994);
   assign  _net_6488 = (in_do&_net_3994);
   assign  _net_6489 = (in_do&_net_3994);
   assign  _net_6490 = (in_do&_net_3994);
   assign  _net_6491 = (in_do&_net_3994);
   assign  _net_6492 = (in_do&_net_3994);
   assign  _net_6493 = (in_do&_net_3994);
   assign  _net_6494 = (in_do&_net_3994);
   assign  _net_6495 = (in_do&_net_3994);
   assign  _net_6496 = (in_do&_net_3994);
   assign  _net_6497 = (in_do&_net_3994);
   assign  _net_6498 = (in_do&_net_3994);
   assign  _net_6499 = (in_do&_net_3994);
   assign  _net_6500 = (in_do&_net_3994);
   assign  _net_6501 = (in_do&_net_3994);
   assign  _net_6502 = (in_do&_net_3994);
   assign  _net_6503 = (in_do&_net_3994);
   assign  _net_6504 = (in_do&_net_3994);
   assign  _net_6505 = (in_do&_net_3994);
   assign  _net_6506 = (in_do&_net_3994);
   assign  _net_6507 = (in_do&_net_3994);
   assign  _net_6508 = (in_do&_net_3994);
   assign  _net_6509 = (in_do&_net_3994);
   assign  _net_6510 = (in_do&_net_3994);
   assign  _net_6511 = (in_do&_net_3994);
   assign  _net_6512 = (in_do&_net_3994);
   assign  _net_6513 = (in_do&_net_3994);
   assign  _net_6514 = (in_do&_net_3994);
   assign  _net_6515 = (in_do&_net_3994);
   assign  _net_6516 = (in_do&_net_3994);
   assign  _net_6517 = (in_do&_net_3994);
   assign  _net_6518 = (in_do&_net_3994);
   assign  _net_6519 = (in_do&_net_3994);
   assign  _net_6520 = (in_do&_net_3994);
   assign  _net_6521 = (in_do&_net_3994);
   assign  _net_6522 = (in_do&_net_3994);
   assign  _net_6523 = (in_do&_net_3994);
   assign  _net_6524 = (in_do&_net_3994);
   assign  _net_6525 = (in_do&_net_3994);
   assign  _net_6526 = (in_do&_net_3994);
   assign  _net_6527 = (in_do&_net_3994);
   assign  _net_6528 = (in_do&_net_3994);
   assign  _net_6529 = (in_do&_net_3994);
   assign  _net_6530 = (in_do&_net_3994);
   assign  _net_6531 = (in_do&_net_3994);
   assign  _net_6532 = (in_do&_net_3994);
   assign  _net_6533 = (in_do&_net_3994);
   assign  _net_6534 = (in_do&_net_3994);
   assign  _net_6535 = (in_do&_net_3994);
   assign  _net_6536 = (in_do&_net_3994);
   assign  _net_6537 = (in_do&_net_3994);
   assign  _net_6538 = (in_do&_net_3994);
   assign  _net_6539 = (in_do&_net_3994);
   assign  _net_6540 = (in_do&_net_3994);
   assign  _net_6541 = (in_do&_net_3994);
   assign  _net_6542 = (in_do&_net_3994);
   assign  _net_6543 = (in_do&_net_3994);
   assign  _net_6544 = (in_do&_net_3994);
   assign  _net_6545 = (in_do&_net_3994);
   assign  _net_6546 = (in_do&_net_3994);
   assign  _net_6547 = (in_do&_net_3994);
   assign  _net_6548 = (in_do&_net_3994);
   assign  _net_6549 = (in_do&_net_3994);
   assign  _net_6550 = (in_do&_net_3994);
   assign  _net_6551 = (in_do&_net_3994);
   assign  _net_6552 = (in_do&_net_3994);
   assign  _net_6553 = (in_do&_net_3994);
   assign  _net_6554 = (in_do&_net_3994);
   assign  _net_6555 = (in_do&_net_3994);
   assign  _net_6556 = (in_do&_net_3994);
   assign  _net_6557 = (in_do&_net_3994);
   assign  _net_6558 = (in_do&_net_3994);
   assign  _net_6559 = (in_do&_net_3994);
   assign  _net_6560 = (in_do&_net_3994);
   assign  _net_6561 = (in_do&_net_3994);
   assign  _net_6562 = (in_do&_net_3994);
   assign  _net_6563 = (in_do&_net_3994);
   assign  _net_6564 = (in_do&_net_3994);
   assign  _net_6565 = (in_do&_net_3994);
   assign  _net_6566 = (in_do&_net_3994);
   assign  _net_6567 = (in_do&_net_3994);
   assign  _net_6568 = (in_do&_net_3994);
   assign  _net_6569 = (in_do&_net_3994);
   assign  _net_6570 = (in_do&_net_3994);
   assign  _net_6571 = (in_do&_net_3994);
   assign  _net_6572 = (in_do&_net_3994);
   assign  _net_6573 = (in_do&_net_3994);
   assign  _net_6574 = (in_do&_net_3994);
   assign  _net_6575 = (in_do&_net_3994);
   assign  _net_6576 = (in_do&_net_3994);
   assign  _net_6577 = (in_do&_net_3994);
   assign  _net_6578 = (in_do&_net_3994);
   assign  _net_6579 = (in_do&_net_3994);
   assign  _net_6580 = (in_do&_net_3994);
   assign  _net_6581 = (in_do&_net_3994);
   assign  _net_6582 = (in_do&_net_3994);
   assign  _net_6583 = (in_do&_net_3994);
   assign  _net_6584 = (in_do&_net_3994);
   assign  _net_6585 = (in_do&_net_3994);
   assign  _net_6586 = (in_do&_net_3994);
   assign  _net_6587 = (in_do&_net_3994);
   assign  _net_6588 = (in_do&_net_3994);
   assign  _net_6589 = (in_do&_net_3994);
   assign  _net_6590 = (in_do&_net_3994);
   assign  _net_6591 = (in_do&_net_3994);
   assign  _net_6592 = (in_do&_net_3994);
   assign  _net_6593 = (in_do&_net_3994);
   assign  _net_6594 = (in_do&_net_3994);
   assign  _net_6595 = (in_do&_net_3994);
   assign  _net_6596 = (in_do&_net_3994);
   assign  _net_6597 = (in_do&_net_3994);
   assign  _net_6598 = (in_do&_net_3994);
   assign  _net_6599 = (in_do&_net_3994);
   assign  _net_6600 = (in_do&_net_3994);
   assign  _net_6601 = (in_do&_net_3994);
   assign  _net_6602 = (in_do&_net_3994);
   assign  _net_6603 = (in_do&_net_3994);
   assign  _net_6604 = (in_do&_net_3994);
   assign  _net_6605 = (in_do&_net_3994);
   assign  _net_6606 = (in_do&_net_3994);
   assign  _net_6607 = (in_do&_net_3994);
   assign  _net_6608 = (in_do&_net_3994);
   assign  _net_6609 = (in_do&_net_3994);
   assign  _net_6610 = (in_do&_net_3994);
   assign  _net_6611 = (in_do&_net_3994);
   assign  _net_6612 = (in_do&_net_3994);
   assign  _net_6613 = (in_do&_net_3994);
   assign  _net_6614 = (in_do&_net_3994);
   assign  _net_6615 = (in_do&_net_3994);
   assign  _net_6616 = (in_do&_net_3994);
   assign  _net_6617 = (in_do&_net_3994);
   assign  _net_6618 = (in_do&_net_3994);
   assign  _net_6619 = (in_do&_net_3994);
   assign  _net_6620 = (in_do&_net_3994);
   assign  _net_6621 = (in_do&_net_3994);
   assign  _net_6622 = (in_do&_net_3994);
   assign  _net_6623 = (in_do&_net_3994);
   assign  _net_6624 = (in_do&_net_3994);
   assign  _net_6625 = (in_do&_net_3994);
   assign  _net_6626 = (in_do&_net_3994);
   assign  _net_6627 = (in_do&_net_3994);
   assign  _net_6628 = (in_do&_net_3994);
   assign  _net_6629 = (in_do&_net_3994);
   assign  _net_6630 = (in_do&_net_3994);
   assign  _net_6631 = (in_do&_net_3994);
   assign  _net_6632 = (in_do&_net_3994);
   assign  _net_6633 = (in_do&_net_3994);
   assign  _net_6634 = (in_do&_net_3994);
   assign  _net_6635 = (in_do&_net_3994);
   assign  _net_6636 = (in_do&_net_3994);
   assign  _net_6637 = (in_do&_net_3994);
   assign  _net_6638 = (in_do&_net_3994);
   assign  _net_6639 = (in_do&_net_3994);
   assign  _net_6640 = (in_do&_net_3994);
   assign  _net_6641 = (in_do&_net_3994);
   assign  _net_6642 = (in_do&_net_3994);
   assign  _net_6643 = (in_do&_net_3994);
   assign  _net_6644 = (in_do&_net_3994);
   assign  _net_6645 = (in_do&_net_3994);
   assign  _net_6646 = (in_do&_net_3994);
   assign  _net_6647 = (in_do&_net_3994);
   assign  _net_6648 = (in_do&_net_3994);
   assign  _net_6649 = (in_do&_net_3994);
   assign  _net_6650 = (in_do&_net_3994);
   assign  _net_6651 = (in_do&_net_3994);
   assign  _net_6652 = (in_do&_net_3994);
   assign  _net_6653 = (in_do&_net_3994);
   assign  _net_6654 = (in_do&_net_3994);
   assign  _net_6655 = (in_do&_net_3994);
   assign  _net_6656 = (in_do&_net_3994);
   assign  _net_6657 = (in_do&_net_3994);
   assign  _net_6658 = (in_do&_net_3994);
   assign  _net_6659 = (in_do&_net_3994);
   assign  _net_6660 = (in_do&_net_3994);
   assign  _net_6661 = (in_do&_net_3994);
   assign  _net_6662 = (in_do&_net_3994);
   assign  _net_6663 = (in_do&_net_3994);
   assign  _net_6664 = (in_do&_net_3994);
   assign  _net_6665 = (in_do&_net_3994);
   assign  _net_6666 = (in_do&_net_3994);
   assign  _net_6667 = (in_do&_net_3994);
   assign  _net_6668 = (in_do&_net_3994);
   assign  _net_6669 = (in_do&_net_3994);
   assign  _net_6670 = (in_do&_net_3994);
   assign  _net_6671 = (in_do&_net_3994);
   assign  _net_6672 = (in_do&_net_3994);
   assign  _net_6673 = (in_do&_net_3994);
   assign  _net_6674 = (in_do&_net_3994);
   assign  _net_6675 = (in_do&_net_3994);
   assign  _net_6676 = (in_do&_net_3994);
   assign  _net_6677 = (in_do&_net_3994);
   assign  _net_6678 = (in_do&_net_3994);
   assign  _net_6679 = (in_do&_net_3994);
   assign  _net_6680 = (in_do&_net_3994);
   assign  _net_6681 = (in_do&_net_3994);
   assign  _net_6682 = (in_do&_net_3994);
   assign  _net_6683 = (in_do&_net_3994);
   assign  _net_6684 = (in_do&_net_3994);
   assign  _net_6685 = (in_do&_net_3994);
   assign  _net_6686 = (in_do&_net_3994);
   assign  _net_6687 = (in_do&_net_3994);
   assign  _net_6688 = (in_do&_net_3994);
   assign  _net_6689 = (in_do&_net_3994);
   assign  _net_6690 = (in_do&_net_3994);
   assign  _net_6691 = (in_do&_net_3994);
   assign  _net_6692 = (in_do&_net_3994);
   assign  _net_6693 = (in_do&_net_3994);
   assign  _net_6694 = (in_do&_net_3994);
   assign  _net_6695 = (in_do&_net_3994);
   assign  _net_6696 = (in_do&_net_3994);
   assign  _net_6697 = (in_do&_net_3994);
   assign  _net_6698 = (in_do&_net_3994);
   assign  _net_6699 = (in_do&_net_3994);
   assign  _net_6700 = (in_do&_net_3994);
   assign  _net_6701 = (in_do&_net_3994);
   assign  _net_6702 = (in_do&_net_3994);
   assign  _net_6703 = (in_do&_net_3994);
   assign  _net_6704 = (in_do&_net_3994);
   assign  _net_6705 = (in_do&_net_3994);
   assign  _net_6706 = (in_do&_net_3994);
   assign  _net_6707 = (in_do&_net_3994);
   assign  _net_6708 = (in_do&_net_3994);
   assign  _net_6709 = (in_do&_net_3994);
   assign  _net_6710 = (in_do&_net_3994);
   assign  _net_6711 = (in_do&_net_3994);
   assign  _net_6712 = (in_do&_net_3994);
   assign  _net_6713 = (in_do&_net_3994);
   assign  _net_6714 = (in_do&_net_3994);
   assign  _net_6715 = (in_do&_net_3994);
   assign  _net_6716 = (in_do&_net_3994);
   assign  _net_6717 = (in_do&_net_3994);
   assign  _net_6718 = (in_do&_net_3994);
   assign  _net_6719 = (in_do&_net_3994);
   assign  _net_6720 = (in_do&_net_3994);
   assign  _net_6721 = (in_do&_net_3994);
   assign  _net_6722 = (in_do&_net_3994);
   assign  _net_6723 = (in_do&_net_3994);
   assign  _net_6724 = (in_do&_net_3994);
   assign  _net_6725 = (in_do&_net_3994);
   assign  _net_6726 = (in_do&_net_3994);
   assign  _net_6727 = (in_do&_net_3994);
   assign  _net_6728 = (in_do&_net_3994);
   assign  _net_6729 = (in_do&_net_3994);
   assign  _net_6730 = (in_do&_net_3994);
   assign  _net_6731 = (in_do&_net_3994);
   assign  _net_6732 = (in_do&_net_3994);
   assign  _net_6733 = (in_do&_net_3994);
   assign  _net_6734 = (in_do&_net_3994);
   assign  _net_6735 = (in_do&_net_3994);
   assign  _net_6736 = (in_do&_net_3994);
   assign  _net_6737 = (in_do&_net_3994);
   assign  _net_6738 = (in_do&_net_3994);
   assign  _net_6739 = (in_do&_net_3994);
   assign  _net_6740 = (in_do&_net_3994);
   assign  _net_6741 = (in_do&_net_3994);
   assign  _net_6742 = (in_do&_net_3994);
   assign  _net_6743 = (in_do&_net_3994);
   assign  _net_6744 = (in_do&_net_3994);
   assign  _net_6745 = (in_do&_net_3994);
   assign  _net_6746 = (in_do&_net_3994);
   assign  _net_6747 = (in_do&_net_3994);
   assign  _net_6748 = (in_do&_net_3994);
   assign  _net_6749 = (in_do&_net_3994);
   assign  _net_6750 = (in_do&_net_3994);
   assign  _net_6751 = (in_do&_net_3994);
   assign  _net_6752 = (in_do&_net_3994);
   assign  _net_6753 = (in_do&_net_3994);
   assign  _net_6754 = (in_do&_net_3994);
   assign  _net_6755 = (in_do&_net_3994);
   assign  _net_6756 = (in_do&_net_3994);
   assign  _net_6757 = (in_do&_net_3994);
   assign  _net_6758 = (in_do&_net_3994);
   assign  _net_6759 = (in_do&_net_3994);
   assign  _net_6760 = (in_do&_net_3994);
   assign  _net_6761 = (in_do&_net_3994);
   assign  _net_6762 = (in_do&_net_3994);
   assign  _net_6763 = (in_do&_net_3994);
   assign  _net_6764 = (in_do&_net_3994);
   assign  _net_6765 = (in_do&_net_3994);
   assign  _net_6766 = (in_do&_net_3994);
   assign  _net_6767 = (in_do&_net_3994);
   assign  _net_6768 = (in_do&_net_3994);
   assign  _net_6769 = (in_do&_net_3994);
   assign  _net_6770 = (in_do&_net_3994);
   assign  _net_6771 = (in_do&_net_3994);
   assign  _net_6772 = (in_do&_net_3994);
   assign  _net_6773 = (in_do&_net_3994);
   assign  _net_6774 = (in_do&_net_3994);
   assign  _net_6775 = (in_do&_net_3994);
   assign  _net_6776 = (in_do&_net_3994);
   assign  _net_6777 = (in_do&_net_3994);
   assign  _net_6778 = (in_do&_net_3994);
   assign  _net_6779 = (in_do&_net_3994);
   assign  _net_6780 = (in_do&_net_3994);
   assign  _net_6781 = (in_do&_net_3994);
   assign  _net_6782 = (in_do&_net_3994);
   assign  _net_6783 = (in_do&_net_3994);
   assign  _net_6784 = (in_do&_net_3994);
   assign  _net_6785 = (in_do&_net_3994);
   assign  _net_6786 = (in_do&_net_3994);
   assign  _net_6787 = (in_do&_net_3994);
   assign  _net_6788 = (in_do&_net_3994);
   assign  _net_6789 = (in_do&_net_3994);
   assign  _net_6790 = (in_do&_net_3994);
   assign  _net_6791 = (in_do&_net_3994);
   assign  _net_6792 = (in_do&_net_3994);
   assign  _net_6793 = (in_do&_net_3994);
   assign  _net_6794 = (in_do&_net_3994);
   assign  _net_6795 = (in_do&_net_3994);
   assign  _net_6796 = (in_do&_net_3994);
   assign  _net_6797 = (in_do&_net_3994);
   assign  _net_6798 = (in_do&_net_3994);
   assign  _net_6799 = (in_do&_net_3994);
   assign  _net_6800 = (in_do&_net_3994);
   assign  _net_6801 = (in_do&_net_3994);
   assign  _net_6802 = (in_do&_net_3994);
   assign  _net_6803 = (in_do&_net_3994);
   assign  _net_6804 = (in_do&_net_3994);
   assign  _net_6805 = (in_do&_net_3994);
   assign  _net_6806 = (in_do&_net_3994);
   assign  _net_6807 = (in_do&_net_3994);
   assign  _net_6808 = (in_do&_net_3994);
   assign  _net_6809 = (in_do&_net_3994);
   assign  _net_6810 = (in_do&_net_3994);
   assign  _net_6811 = (in_do&_net_3994);
   assign  _net_6812 = (in_do&_net_3994);
   assign  _net_6813 = (in_do&_net_3994);
   assign  _net_6814 = (in_do&_net_3994);
   assign  _net_6815 = (in_do&_net_3994);
   assign  _net_6816 = (in_do&_net_3994);
   assign  _net_6817 = (in_do&_net_3994);
   assign  _net_6818 = (in_do&_net_3994);
   assign  _net_6819 = (in_do&_net_3994);
   assign  _net_6820 = (in_do&_net_3994);
   assign  _net_6821 = (in_do&_net_3994);
   assign  _net_6822 = (in_do&_net_3994);
   assign  _net_6823 = (in_do&_net_3994);
   assign  _net_6824 = (in_do&_net_3994);
   assign  _net_6825 = (in_do&_net_3994);
   assign  _net_6826 = (in_do&_net_3994);
   assign  _net_6827 = (in_do&_net_3994);
   assign  _net_6828 = (in_do&_net_3994);
   assign  _net_6829 = (in_do&_net_3994);
   assign  _net_6830 = (in_do&_net_3994);
   assign  _net_6831 = (in_do&_net_3994);
   assign  _net_6832 = (in_do&_net_3994);
   assign  _net_6833 = (in_do&_net_3994);
   assign  _net_6834 = (in_do&_net_3994);
   assign  _net_6835 = (in_do&_net_3994);
   assign  _net_6836 = (in_do&_net_3994);
   assign  _net_6837 = (in_do&_net_3994);
   assign  _net_6838 = (in_do&_net_3994);
   assign  _net_6839 = (in_do&_net_3994);
   assign  _net_6840 = (in_do&_net_3994);
   assign  _net_6841 = (in_do&_net_3994);
   assign  _net_6842 = (in_do&_net_3994);
   assign  _net_6843 = (in_do&_net_3994);
   assign  _net_6844 = (in_do&_net_3994);
   assign  _net_6845 = (in_do&_net_3994);
   assign  _net_6846 = (in_do&_net_3994);
   assign  _net_6847 = (in_do&_net_3994);
   assign  _net_6848 = (in_do&_net_3994);
   assign  _net_6849 = (in_do&_net_3994);
   assign  _net_6850 = (in_do&_net_3994);
   assign  _net_6851 = (in_do&_net_3994);
   assign  _net_6852 = (in_do&_net_3994);
   assign  _net_6853 = (in_do&_net_3994);
   assign  _net_6854 = (in_do&_net_3994);
   assign  _net_6855 = (in_do&_net_3994);
   assign  _net_6856 = (in_do&_net_3994);
   assign  _net_6857 = (in_do&_net_3994);
   assign  _net_6858 = (in_do&_net_3994);
   assign  _net_6859 = (in_do&_net_3994);
   assign  _net_6860 = (in_do&_net_3994);
   assign  _net_6861 = (in_do&_net_3994);
   assign  _net_6862 = (in_do&_net_3994);
   assign  _net_6863 = (in_do&_net_3994);
   assign  _net_6864 = (in_do&_net_3994);
   assign  _net_6865 = (in_do&_net_3994);
   assign  _net_6866 = (in_do&_net_3994);
   assign  _net_6867 = (in_do&_net_3994);
   assign  _net_6868 = (in_do&_net_3994);
   assign  _net_6869 = (in_do&_net_3994);
   assign  _net_6870 = (in_do&_net_3994);
   assign  _net_6871 = (in_do&_net_3994);
   assign  _net_6872 = (in_do&_net_3994);
   assign  _net_6873 = (in_do&_net_3994);
   assign  _net_6874 = (in_do&_net_3994);
   assign  _net_6875 = (in_do&_net_3994);
   assign  _net_6876 = (in_do&_net_3994);
   assign  _net_6877 = (in_do&_net_3994);
   assign  _net_6878 = (in_do&_net_3994);
   assign  _net_6879 = (in_do&_net_3994);
   assign  _net_6880 = (in_do&_net_3994);
   assign  _net_6881 = (in_do&_net_3994);
   assign  _net_6882 = (in_do&_net_3994);
   assign  _net_6883 = (in_do&_net_3994);
   assign  _net_6884 = (in_do&_net_3994);
   assign  _net_6885 = (in_do&_net_3994);
   assign  _net_6886 = (in_do&_net_3994);
   assign  _net_6887 = (in_do&_net_3994);
   assign  _net_6888 = (in_do&_net_3994);
   assign  _net_6889 = (in_do&_net_3994);
   assign  _net_6890 = (in_do&_net_3994);
   assign  _net_6891 = (in_do&_net_3994);
   assign  _net_6892 = (in_do&_net_3994);
   assign  _net_6893 = (in_do&_net_3994);
   assign  _net_6894 = (in_do&_net_3994);
   assign  _net_6895 = (in_do&_net_3994);
   assign  _net_6896 = (in_do&_net_3994);
   assign  _net_6897 = (in_do&_net_3994);
   assign  _net_6898 = (in_do&_net_3994);
   assign  _net_6899 = (in_do&_net_3994);
   assign  _net_6900 = (in_do&_net_3994);
   assign  _net_6901 = (in_do&_net_3994);
   assign  _net_6902 = (in_do&_net_3994);
   assign  _net_6903 = (in_do&_net_3994);
   assign  _net_6904 = (in_do&_net_3994);
   assign  _net_6905 = (in_do&_net_3994);
   assign  _net_6906 = (in_do&_net_3994);
   assign  _net_6907 = (in_do&_net_3994);
   assign  _net_6908 = (in_do&_net_3994);
   assign  _net_6909 = (in_do&_net_3994);
   assign  _net_6910 = (in_do&_net_3994);
   assign  _net_6911 = (in_do&_net_3994);
   assign  _net_6912 = (in_do&_net_3994);
   assign  _net_6913 = (in_do&_net_3994);
   assign  _net_6914 = (in_do&_net_3994);
   assign  _net_6915 = (in_do&_net_3994);
   assign  _net_6916 = (in_do&_net_3994);
   assign  _net_6917 = (in_do&_net_3994);
   assign  _net_6918 = (in_do&_net_3994);
   assign  _net_6919 = (in_do&_net_3994);
   assign  _net_6920 = (in_do&_net_3994);
   assign  _net_6921 = (in_do&_net_3994);
   assign  _net_6922 = (in_do&_net_3994);
   assign  _net_6923 = (in_do&_net_3994);
   assign  _net_6924 = (in_do&_net_3994);
   assign  _net_6925 = (in_do&_net_3994);
   assign  _net_6926 = (in_do&_net_3994);
   assign  _net_6927 = (in_do&_net_3994);
   assign  _net_6928 = (in_do&_net_3994);
   assign  _net_6929 = (in_do&_net_3994);
   assign  _net_6930 = (in_do&_net_3994);
   assign  _net_6931 = (in_do&_net_3994);
   assign  _net_6932 = (in_do&_net_3994);
   assign  _net_6933 = (in_do&_net_3994);
   assign  _net_6934 = (in_do&_net_3994);
   assign  _net_6935 = (in_do&_net_3994);
   assign  _net_6936 = (in_do&_net_3994);
   assign  _net_6937 = (in_do&_net_3994);
   assign  _net_6938 = (in_do&_net_3994);
   assign  _net_6939 = (in_do&_net_3994);
   assign  _net_6940 = (in_do&_net_3994);
   assign  _net_6941 = (in_do&_net_3994);
   assign  _net_6942 = (in_do&_net_3994);
   assign  _net_6943 = (in_do&_net_3994);
   assign  _net_6944 = (in_do&_net_3994);
   assign  _net_6945 = (in_do&_net_3994);
   assign  _net_6946 = (in_do&_net_3994);
   assign  _net_6947 = (in_do&_net_3994);
   assign  _net_6948 = (in_do&_net_3994);
   assign  _net_6949 = (in_do&_net_3994);
   assign  _net_6950 = (in_do&_net_3994);
   assign  _net_6951 = (in_do&_net_3994);
   assign  _net_6952 = (in_do&_net_3994);
   assign  _net_6953 = (in_do&_net_3994);
   assign  _net_6954 = (in_do&_net_3994);
   assign  _net_6955 = (in_do&_net_3994);
   assign  _net_6956 = (in_do&_net_3994);
   assign  _net_6957 = (in_do&_net_3994);
   assign  _net_6958 = (in_do&_net_3994);
   assign  _net_6959 = (in_do&_net_3994);
   assign  _net_6960 = (in_do&_net_3994);
   assign  _net_6961 = (in_do&_net_3994);
   assign  _net_6962 = (in_do&_net_3994);
   assign  _net_6963 = (in_do&_net_3994);
   assign  _net_6964 = (in_do&_net_3994);
   assign  _net_6965 = (in_do&_net_3994);
   assign  _net_6966 = (in_do&_net_3994);
   assign  _net_6967 = (in_do&_net_3994);
   assign  _net_6968 = (in_do&_net_3994);
   assign  _net_6969 = (in_do&_net_3994);
   assign  _net_6970 = (in_do&_net_3994);
   assign  _net_6971 = (in_do&_net_3994);
   assign  _net_6972 = (in_do&_net_3994);
   assign  _net_6973 = (in_do&_net_3994);
   assign  _net_6974 = (in_do&_net_3994);
   assign  _net_6975 = (in_do&_net_3994);
   assign  _net_6976 = (in_do&_net_3994);
   assign  _net_6977 = (in_do&_net_3994);
   assign  _net_6978 = (in_do&_net_3994);
   assign  _net_6979 = (in_do&_net_3994);
   assign  _net_6980 = (in_do&_net_3994);
   assign  _net_6981 = (in_do&_net_3994);
   assign  _net_6982 = (in_do&_net_3994);
   assign  _net_6983 = (in_do&_net_3994);
   assign  _net_6984 = (in_do&_net_3994);
   assign  _net_6985 = (in_do&_net_3994);
   assign  _net_6986 = (in_do&_net_3994);
   assign  _net_6987 = (in_do&_net_3994);
   assign  _net_6988 = (in_do&_net_3994);
   assign  _net_6989 = (in_do&_net_3994);
   assign  _net_6990 = (in_do&_net_3994);
   assign  _net_6991 = (in_do&_net_3994);
   assign  _net_6992 = (in_do&_net_3994);
   assign  _net_6993 = (in_do&_net_3994);
   assign  _net_6994 = (in_do&_net_3994);
   assign  _net_6995 = (in_do&_net_3994);
   assign  _net_6996 = (in_do&_net_3994);
   assign  _net_6997 = (in_do&_net_3994);
   assign  _net_6998 = (in_do&_net_3994);
   assign  _net_6999 = (in_do&_net_3994);
   assign  _net_7000 = (in_do&_net_3994);
   assign  _net_7001 = (in_do&_net_3994);
   assign  _net_7002 = (in_do&_net_3994);
   assign  _net_7003 = (in_do&_net_3994);
   assign  _net_7004 = (in_do&_net_3994);
   assign  _net_7005 = (in_do&_net_3994);
   assign  _net_7006 = (in_do&_net_3994);
   assign  _net_7007 = (in_do&_net_3994);
   assign  _net_7008 = (in_do&_net_3994);
   assign  _net_7009 = (in_do&_net_3994);
   assign  _net_7010 = (in_do&_net_3994);
   assign  _net_7011 = (in_do&_net_3994);
   assign  _net_7012 = (in_do&_net_3994);
   assign  _net_7013 = (in_do&_net_3994);
   assign  _net_7014 = (in_do&_net_3994);
   assign  _net_7015 = (in_do&_net_3994);
   assign  _net_7016 = (in_do&_net_3994);
   assign  _net_7017 = (in_do&_net_3994);
   assign  _net_7018 = (in_do&_net_3994);
   assign  _net_7019 = (in_do&_net_3994);
   assign  _net_7020 = (in_do&_net_3994);
   assign  _net_7021 = (in_do&_net_3994);
   assign  _net_7022 = (in_do&_net_3994);
   assign  _net_7023 = (in_do&_net_3994);
   assign  _net_7024 = (in_do&_net_3994);
   assign  _net_7025 = (in_do&_net_3994);
   assign  _net_7026 = (in_do&_net_3994);
   assign  _net_7027 = (in_do&_net_3994);
   assign  _net_7028 = (in_do&_net_3994);
   assign  _net_7029 = (in_do&_net_3994);
   assign  _net_7030 = (in_do&_net_3994);
   assign  _net_7031 = (in_do&_net_3994);
   assign  _net_7032 = (in_do&_net_3994);
   assign  _net_7033 = (in_do&_net_3994);
   assign  _net_7034 = (in_do&_net_3994);
   assign  _net_7035 = (in_do&_net_3994);
   assign  _net_7036 = (in_do&_net_3994);
   assign  _net_7037 = (in_do&_net_3994);
   assign  _net_7038 = (in_do&_net_3994);
   assign  _net_7039 = (in_do&_net_3994);
   assign  _net_7040 = (in_do&_net_3994);
   assign  _net_7041 = (in_do&_net_3994);
   assign  _net_7042 = (in_do&_net_3994);
   assign  _net_7043 = (in_do&_net_3994);
   assign  _net_7044 = (in_do&_net_3994);
   assign  _net_7045 = (in_do&_net_3994);
   assign  _net_7046 = (in_do&_net_3994);
   assign  _net_7047 = (in_do&_net_3994);
   assign  _net_7048 = (in_do&_net_3994);
   assign  _net_7049 = (in_do&_net_3994);
   assign  _net_7050 = (in_do&_net_3994);
   assign  _net_7051 = (in_do&_net_3994);
   assign  _net_7052 = (in_do&_net_3994);
   assign  _net_7053 = (in_do&_net_3994);
   assign  _net_7054 = (in_do&_net_3994);
   assign  _net_7055 = (in_do&_net_3994);
   assign  _net_7056 = (in_do&_net_3994);
   assign  _net_7057 = (in_do&_net_3994);
   assign  _net_7058 = (in_do&_net_3994);
   assign  _net_7059 = (in_do&_net_3994);
   assign  _net_7060 = (in_do&_net_3994);
   assign  _net_7061 = (in_do&_net_3994);
   assign  _net_7062 = (in_do&_net_3994);
   assign  _net_7063 = (in_do&_net_3994);
   assign  _net_7064 = (in_do&_net_3994);
   assign  _net_7065 = (in_do&_net_3994);
   assign  _net_7066 = (in_do&_net_3994);
   assign  _net_7067 = (in_do&_net_3994);
   assign  _net_7068 = (in_do&_net_3994);
   assign  _net_7069 = (in_do&_net_3994);
   assign  _net_7070 = (in_do&_net_3994);
   assign  _net_7071 = (in_do&_net_3994);
   assign  _net_7072 = (in_do&_net_3994);
   assign  _net_7073 = (in_do&_net_3994);
   assign  _net_7074 = (in_do&_net_3994);
   assign  _net_7075 = (in_do&_net_3994);
   assign  _net_7076 = (in_do&_net_3994);
   assign  _net_7077 = (in_do&_net_3994);
   assign  _net_7078 = (in_do&_net_3994);
   assign  _net_7079 = (in_do&_net_3994);
   assign  _net_7080 = (in_do&_net_3994);
   assign  _net_7081 = (in_do&_net_3994);
   assign  _net_7082 = (in_do&_net_3994);
   assign  _net_7083 = (in_do&_net_3994);
   assign  _net_7084 = (in_do&_net_3994);
   assign  _net_7085 = (in_do&_net_3994);
   assign  _net_7086 = (in_do&_net_3994);
   assign  _net_7087 = (in_do&_net_3994);
   assign  _net_7088 = (in_do&_net_3994);
   assign  _net_7089 = (in_do&_net_3994);
   assign  _net_7090 = (in_do&_net_3994);
   assign  _net_7091 = (in_do&_net_3994);
   assign  _net_7092 = (in_do&_net_3994);
   assign  _net_7093 = (in_do&_net_3994);
   assign  _net_7094 = (in_do&_net_3994);
   assign  _net_7095 = (in_do&_net_3994);
   assign  _net_7096 = (in_do&_net_3994);
   assign  _net_7097 = (in_do&_net_3994);
   assign  _net_7098 = (in_do&_net_3994);
   assign  _net_7099 = (in_do&_net_3994);
   assign  _net_7100 = (in_do&_net_3994);
   assign  _net_7101 = (in_do&_net_3994);
   assign  _net_7102 = (in_do&_net_3994);
   assign  _net_7103 = (in_do&_net_3994);
   assign  _net_7104 = (in_do&_net_3994);
   assign  _net_7105 = (in_do&_net_3994);
   assign  _net_7106 = (in_do&_net_3994);
   assign  _net_7107 = (in_do&_net_3994);
   assign  _net_7108 = (in_do&_net_3994);
   assign  _net_7109 = (in_do&_net_3994);
   assign  _net_7110 = (in_do&_net_3994);
   assign  _net_7111 = (in_do&_net_3994);
   assign  _net_7112 = (in_do&_net_3994);
   assign  _net_7113 = (in_do&_net_3994);
   assign  _net_7114 = (in_do&_net_3994);
   assign  _net_7115 = (in_do&_net_3994);
   assign  _net_7116 = (in_do&_net_3994);
   assign  _net_7117 = (in_do&_net_3994);
   assign  _net_7118 = (in_do&_net_3994);
   assign  _net_7119 = (in_do&_net_3994);
   assign  _net_7120 = (in_do&_net_3994);
   assign  _net_7121 = (in_do&_net_3994);
   assign  _net_7122 = (in_do&_net_3994);
   assign  _net_7123 = (in_do&_net_3994);
   assign  _net_7124 = (in_do&_net_3994);
   assign  _net_7125 = (in_do&_net_3994);
   assign  _net_7126 = (in_do&_net_3994);
   assign  _net_7127 = (in_do&_net_3994);
   assign  _net_7128 = (in_do&_net_3994);
   assign  _net_7129 = (in_do&_net_3994);
   assign  _net_7130 = (in_do&_net_3994);
   assign  _net_7131 = (in_do&_net_3994);
   assign  _net_7132 = (in_do&_net_3994);
   assign  _net_7133 = (in_do&_net_3994);
   assign  _net_7134 = (in_do&_net_3994);
   assign  _net_7135 = (in_do&_net_3994);
   assign  _net_7136 = (in_do&_net_3994);
   assign  _net_7137 = (in_do&_net_3994);
   assign  _net_7138 = (in_do&_net_3994);
   assign  _net_7139 = (in_do&_net_3994);
   assign  _net_7140 = (in_do&_net_3994);
   assign  _net_7141 = (in_do&_net_3994);
   assign  _net_7142 = (in_do&_net_3994);
   assign  _net_7143 = (in_do&_net_3994);
   assign  _net_7144 = (in_do&_net_3994);
   assign  _net_7145 = (in_do&_net_3994);
   assign  _net_7146 = (in_do&_net_3994);
   assign  _net_7147 = (in_do&_net_3994);
   assign  _net_7148 = (in_do&_net_3994);
   assign  _net_7149 = (in_do&_net_3994);
   assign  _net_7150 = (in_do&_net_3994);
   assign  _net_7151 = (in_do&_net_3994);
   assign  _net_7152 = (in_do&_net_3994);
   assign  _net_7153 = (in_do&_net_3994);
   assign  _net_7154 = (in_do&_net_3994);
   assign  _net_7155 = (in_do&_net_3994);
   assign  _net_7156 = (in_do&_net_3994);
   assign  _net_7157 = (in_do&_net_3994);
   assign  _net_7158 = (in_do&_net_3994);
   assign  _net_7159 = (in_do&_net_3994);
   assign  _net_7160 = (in_do&_net_3994);
   assign  _net_7161 = (in_do&_net_3994);
   assign  _net_7162 = (in_do&_net_3994);
   assign  _net_7163 = (in_do&_net_3994);
   assign  _net_7164 = (in_do&_net_3994);
   assign  _net_7165 = (in_do&_net_3994);
   assign  _net_7166 = (in_do&_net_3994);
   assign  _net_7167 = (in_do&_net_3994);
   assign  _net_7168 = (in_do&_net_3994);
   assign  _net_7169 = (in_do&_net_3994);
   assign  _net_7170 = (in_do&_net_3994);
   assign  _net_7171 = (in_do&_net_3994);
   assign  _net_7172 = (in_do&_net_3994);
   assign  _net_7173 = (in_do&_net_3994);
   assign  _net_7174 = (in_do&_net_3994);
   assign  _net_7175 = (in_do&_net_3994);
   assign  _net_7176 = (in_do&_net_3994);
   assign  _net_7177 = (in_do&_net_3994);
   assign  _net_7178 = (in_do&_net_3994);
   assign  _net_7179 = (in_do&_net_3994);
   assign  _net_7180 = (in_do&_net_3994);
   assign  _net_7181 = (in_do&_net_3994);
   assign  _net_7182 = (in_do&_net_3994);
   assign  _net_7183 = (in_do&_net_3994);
   assign  _net_7184 = (in_do&_net_3994);
   assign  _net_7185 = (in_do&_net_3994);
   assign  _net_7186 = (in_do&_net_3994);
   assign  _net_7187 = (in_do&_net_3994);
   assign  _net_7188 = (in_do&_net_3994);
   assign  _net_7189 = (in_do&_net_3994);
   assign  _net_7190 = (in_do&_net_3994);
   assign  _net_7191 = (in_do&_net_3994);
   assign  _net_7192 = (in_do&_net_3994);
   assign  _net_7193 = (in_do&_net_3994);
   assign  _net_7194 = (in_do&_net_3994);
   assign  _net_7195 = (in_do&_net_3994);
   assign  _net_7196 = (in_do&_net_3994);
   assign  _net_7197 = (in_do&_net_3994);
   assign  _net_7198 = (in_do&_net_3994);
   assign  _net_7199 = (in_do&_net_3994);
   assign  _net_7200 = (in_do&_net_3994);
   assign  _net_7201 = (in_do&_net_3994);
   assign  _net_7202 = (in_do&_net_3994);
   assign  _net_7203 = (in_do&_net_3994);
   assign  _net_7204 = (in_do&_net_3994);
   assign  _net_7205 = (in_do&_net_3994);
   assign  _net_7206 = (in_do&_net_3994);
   assign  _net_7207 = (in_do&_net_3994);
   assign  _net_7208 = (in_do&_net_3994);
   assign  _net_7209 = (in_do&_net_3994);
   assign  _net_7210 = (in_do&_net_3994);
   assign  _net_7211 = (in_do&_net_3994);
   assign  _net_7212 = (in_do&_net_3994);
   assign  _net_7213 = (in_do&_net_3994);
   assign  _net_7214 = (in_do&_net_3994);
   assign  _net_7215 = (in_do&_net_3994);
   assign  _net_7216 = (in_do&_net_3994);
   assign  _net_7217 = (in_do&_net_3994);
   assign  _net_7218 = (in_do&_net_3994);
   assign  _net_7219 = (in_do&_net_3994);
   assign  _net_7220 = (in_do&_net_3994);
   assign  _net_7221 = (in_do&_net_3994);
   assign  _net_7222 = (in_do&_net_3994);
   assign  _net_7223 = (in_do&_net_3994);
   assign  _net_7224 = (in_do&_net_3994);
   assign  _net_7225 = (in_do&_net_3994);
   assign  _net_7226 = (in_do&_net_3994);
   assign  _net_7227 = (in_do&_net_3994);
   assign  _net_7228 = (in_do&_net_3994);
   assign  _net_7229 = (in_do&_net_3994);
   assign  _net_7230 = (in_do&_net_3994);
   assign  _net_7231 = (in_do&_net_3994);
   assign  _net_7232 = (in_do&_net_3994);
   assign  _net_7233 = (in_do&_net_3994);
   assign  _net_7234 = (in_do&_net_3994);
   assign  _net_7235 = (in_do&_net_3994);
   assign  _net_7236 = (in_do&_net_3994);
   assign  _net_7237 = (in_do&_net_3994);
   assign  _net_7238 = (in_do&_net_3994);
   assign  _net_7239 = (in_do&_net_3994);
   assign  _net_7240 = (in_do&_net_3994);
   assign  _net_7241 = (in_do&_net_3994);
   assign  _net_7242 = (in_do&_net_3994);
   assign  _net_7243 = (in_do&_net_3994);
   assign  _net_7244 = (in_do&_net_3994);
   assign  _net_7245 = (in_do&_net_3994);
   assign  _net_7246 = (in_do&_net_3994);
   assign  _net_7247 = (in_do&_net_3994);
   assign  _net_7248 = (in_do&_net_3994);
   assign  _net_7249 = (in_do&_net_3994);
   assign  _net_7250 = (in_do&_net_3994);
   assign  _net_7251 = (in_do&_net_3994);
   assign  _net_7252 = (in_do&_net_3994);
   assign  _net_7253 = (in_do&_net_3994);
   assign  _net_7254 = (in_do&_net_3994);
   assign  _net_7255 = (in_do&_net_3994);
   assign  _net_7256 = (in_do&_net_3994);
   assign  _net_7257 = (in_do&_net_3994);
   assign  _net_7258 = (in_do&_net_3994);
   assign  _net_7259 = (in_do&_net_3994);
   assign  _net_7260 = (in_do&_net_3994);
   assign  _net_7261 = (in_do&_net_3994);
   assign  _net_7262 = (in_do&_net_3994);
   assign  _net_7263 = (in_do&_net_3994);
   assign  _net_7264 = (in_do&_net_3994);
   assign  _net_7265 = (in_do&_net_3994);
   assign  _net_7266 = (in_do&_net_3994);
   assign  _net_7267 = (in_do&_net_3994);
   assign  _net_7268 = (in_do&_net_3994);
   assign  _net_7269 = (in_do&_net_3994);
   assign  _net_7270 = (in_do&_net_3994);
   assign  _net_7271 = (in_do&_net_3994);
   assign  _net_7272 = (in_do&_net_3994);
   assign  _net_7273 = (in_do&_net_3994);
   assign  _net_7274 = (in_do&_net_3994);
   assign  _net_7275 = (in_do&_net_3994);
   assign  _net_7276 = (in_do&_net_3994);
   assign  _net_7277 = (in_do&_net_3994);
   assign  _net_7278 = (in_do&_net_3994);
   assign  _net_7279 = (in_do&_net_3994);
   assign  _net_7280 = (in_do&_net_3994);
   assign  _net_7281 = (in_do&_net_3994);
   assign  _net_7282 = (in_do&_net_3994);
   assign  _net_7283 = (in_do&_net_3994);
   assign  _net_7284 = (in_do&_net_3994);
   assign  _net_7285 = (in_do&_net_3994);
   assign  _net_7286 = (in_do&_net_3994);
   assign  _net_7287 = (in_do&_net_3994);
   assign  _net_7288 = (in_do&_net_3994);
   assign  _net_7289 = (in_do&_net_3994);
   assign  _net_7290 = (in_do&_net_3994);
   assign  _net_7291 = (in_do&_net_3994);
   assign  _net_7292 = (in_do&_net_3994);
   assign  _net_7293 = (in_do&_net_3994);
   assign  _net_7294 = (in_do&_net_3994);
   assign  _net_7295 = (in_do&_net_3994);
   assign  _net_7296 = (in_do&_net_3994);
   assign  _net_7297 = (in_do&_net_3994);
   assign  _net_7298 = (in_do&_net_3994);
   assign  _net_7299 = (in_do&_net_3994);
   assign  _net_7300 = (in_do&_net_3994);
   assign  _net_7301 = (in_do&_net_3994);
   assign  _net_7302 = (in_do&_net_3994);
   assign  _net_7303 = (in_do&_net_3994);
   assign  _net_7304 = (in_do&_net_3994);
   assign  _net_7305 = (in_do&_net_3994);
   assign  _net_7306 = (in_do&_net_3994);
   assign  _net_7307 = (in_do&_net_3994);
   assign  _net_7308 = (in_do&_net_3994);
   assign  _net_7309 = (in_do&_net_3994);
   assign  _net_7310 = (in_do&_net_3994);
   assign  _net_7311 = (in_do&_net_3994);
   assign  _net_7312 = (in_do&_net_3994);
   assign  _net_7313 = (in_do&_net_3994);
   assign  _net_7314 = (in_do&_net_3994);
   assign  _net_7315 = (in_do&_net_3994);
   assign  _net_7316 = (in_do&_net_3994);
   assign  _net_7317 = (in_do&_net_3994);
   assign  _net_7318 = (in_do&_net_3994);
   assign  _net_7319 = (in_do&_net_3994);
   assign  _net_7320 = (in_do&_net_3994);
   assign  _net_7321 = (in_do&_net_3994);
   assign  _net_7322 = (in_do&_net_3994);
   assign  _net_7323 = (in_do&_net_3994);
   assign  _net_7324 = (in_do&_net_3994);
   assign  _net_7325 = (in_do&_net_3994);
   assign  _net_7326 = (in_do&_net_3994);
   assign  _net_7327 = (in_do&_net_3994);
   assign  _net_7328 = (in_do&_net_3994);
   assign  _net_7329 = (in_do&_net_3994);
   assign  _net_7330 = (in_do&_net_3994);
   assign  _net_7331 = (in_do&_net_3994);
   assign  _net_7332 = (in_do&_net_3994);
   assign  _net_7333 = (in_do&_net_3994);
   assign  _net_7334 = (in_do&_net_3994);
   assign  _net_7335 = (in_do&_net_3994);
   assign  _net_7336 = (in_do&_net_3994);
   assign  _net_7337 = (in_do&_net_3994);
   assign  _net_7338 = (in_do&_net_3994);
   assign  _net_7339 = (in_do&_net_3994);
   assign  _net_7340 = (in_do&_net_3994);
   assign  _net_7341 = (in_do&_net_3994);
   assign  _net_7342 = (in_do&_net_3994);
   assign  _net_7343 = (in_do&_net_3994);
   assign  _net_7344 = (in_do&_net_3994);
   assign  _net_7345 = (in_do&_net_3994);
   assign  _net_7346 = (in_do&_net_3994);
   assign  _net_7347 = (in_do&_net_3994);
   assign  _net_7348 = (in_do&_net_3994);
   assign  _net_7349 = (in_do&_net_3994);
   assign  _net_7350 = (in_do&_net_3994);
   assign  _net_7351 = (in_do&_net_3994);
   assign  _net_7352 = (in_do&_net_3994);
   assign  _net_7353 = (in_do&_net_3994);
   assign  _net_7354 = (in_do&_net_3994);
   assign  _net_7355 = (in_do&_net_3994);
   assign  _net_7356 = (in_do&_net_3994);
   assign  _net_7357 = (in_do&_net_3994);
   assign  _net_7358 = (in_do&_net_3994);
   assign  _net_7359 = (in_do&_net_3994);
   assign  _net_7360 = (in_do&_net_3994);
   assign  _net_7361 = (in_do&_net_3994);
   assign  _net_7362 = (in_do&_net_3994);
   assign  _net_7363 = (in_do&_net_3994);
   assign  _net_7364 = (in_do&_net_3994);
   assign  _net_7365 = (in_do&_net_3994);
   assign  _net_7366 = (in_do&_net_3994);
   assign  _net_7367 = (in_do&_net_3994);
   assign  _net_7368 = (in_do&_net_3994);
   assign  _net_7369 = (in_do&_net_3994);
   assign  _net_7370 = (in_do&_net_3994);
   assign  _net_7371 = (in_do&_net_3994);
   assign  _net_7372 = (in_do&_net_3994);
   assign  _net_7373 = (in_do&_net_3994);
   assign  _net_7374 = (in_do&_net_3994);
   assign  _net_7375 = (in_do&_net_3994);
   assign  _net_7376 = (in_do&_net_3994);
   assign  _net_7377 = (in_do&_net_3994);
   assign  _net_7378 = (in_do&_net_3994);
   assign  _net_7379 = (in_do&_net_3994);
   assign  _net_7380 = (in_do&_net_3994);
   assign  _net_7381 = (in_do&_net_3994);
   assign  _net_7382 = (in_do&_net_3994);
   assign  _net_7383 = (in_do&_net_3994);
   assign  _net_7384 = (in_do&_net_3994);
   assign  _net_7385 = (in_do&_net_3994);
   assign  _net_7386 = (in_do&_net_3994);
   assign  _net_7387 = (in_do&_net_3994);
   assign  _net_7388 = (in_do&_net_3994);
   assign  _net_7389 = (in_do&_net_3994);
   assign  _net_7390 = (in_do&_net_3994);
   assign  _net_7391 = (in_do&_net_3994);
   assign  _net_7392 = (in_do&_net_3994);
   assign  _net_7393 = (in_do&_net_3994);
   assign  _net_7394 = (in_do&_net_3994);
   assign  _net_7395 = (in_do&_net_3994);
   assign  _net_7396 = (in_do&_net_3994);
   assign  _net_7397 = (in_do&_net_3994);
   assign  _net_7398 = (in_do&_net_3994);
   assign  _net_7399 = (in_do&_net_3994);
   assign  _net_7400 = (in_do&_net_3994);
   assign  _net_7401 = (in_do&_net_3994);
   assign  _net_7402 = (in_do&_net_3994);
   assign  _net_7403 = (in_do&_net_3994);
   assign  _net_7404 = (in_do&_net_3994);
   assign  _net_7405 = (in_do&_net_3994);
   assign  _net_7406 = (in_do&_net_3994);
   assign  _net_7407 = (in_do&_net_3994);
   assign  _net_7408 = (in_do&_net_3994);
   assign  _net_7409 = (in_do&_net_3994);
   assign  _net_7410 = (in_do&_net_3994);
   assign  _net_7411 = (in_do&_net_3994);
   assign  _net_7412 = (in_do&_net_3994);
   assign  _net_7413 = (in_do&_net_3994);
   assign  _net_7414 = (in_do&_net_3994);
   assign  _net_7415 = (in_do&_net_3994);
   assign  _net_7416 = (in_do&_net_3994);
   assign  _net_7417 = (in_do&_net_3994);
   assign  _net_7418 = (in_do&_net_3994);
   assign  _net_7419 = (in_do&_net_3994);
   assign  _net_7420 = (in_do&_net_3994);
   assign  _net_7421 = (in_do&_net_3994);
   assign  _net_7422 = (in_do&_net_3994);
   assign  _net_7423 = (in_do&_net_3994);
   assign  _net_7424 = (in_do&_net_3994);
   assign  _net_7425 = (in_do&_net_3994);
   assign  _net_7426 = (in_do&_net_3994);
   assign  _net_7427 = (in_do&_net_3994);
   assign  _net_7428 = (in_do&_net_3994);
   assign  _net_7429 = (in_do&_net_3994);
   assign  _net_7430 = (in_do&_net_3994);
   assign  _net_7431 = (in_do&_net_3994);
   assign  _net_7432 = (in_do&_net_3994);
   assign  _net_7433 = (in_do&_net_3994);
   assign  _net_7434 = (in_do&_net_3994);
   assign  _net_7435 = (in_do&_net_3994);
   assign  _net_7436 = (in_do&_net_3994);
   assign  _net_7437 = (in_do&_net_3994);
   assign  _net_7438 = (in_do&_net_3994);
   assign  _net_7439 = (in_do&_net_3994);
   assign  _net_7440 = (in_do&_net_3994);
   assign  _net_7441 = (in_do&_net_3994);
   assign  _net_7442 = (in_do&_net_3994);
   assign  _net_7443 = (in_do&_net_3994);
   assign  _net_7444 = (in_do&_net_3994);
   assign  _net_7445 = (in_do&_net_3994);
   assign  _net_7446 = (in_do&_net_3994);
   assign  _net_7447 = (in_do&_net_3994);
   assign  _net_7448 = (in_do&_net_3994);
   assign  _net_7449 = (in_do&_net_3994);
   assign  _net_7450 = (in_do&_net_3994);
   assign  _net_7451 = (in_do&_net_3994);
   assign  _net_7452 = (in_do&_net_3994);
   assign  _net_7453 = (in_do&_net_3994);
   assign  _net_7454 = (in_do&_net_3994);
   assign  _net_7455 = (in_do&_net_3994);
   assign  _net_7456 = (in_do&_net_3994);
   assign  _net_7457 = (in_do&_net_3994);
   assign  _net_7458 = (in_do&_net_3994);
   assign  _net_7459 = (in_do&_net_3994);
   assign  _net_7460 = (in_do&_net_3994);
   assign  _net_7461 = (in_do&_net_3994);
   assign  _net_7462 = (in_do&_net_3994);
   assign  _net_7463 = (in_do&_net_3994);
   assign  _net_7464 = (in_do&_net_3994);
   assign  _net_7465 = (in_do&_net_3994);
   assign  _net_7466 = (in_do&_net_3994);
   assign  _net_7467 = (in_do&_net_3994);
   assign  _net_7468 = (in_do&_net_3994);
   assign  _net_7469 = (in_do&_net_3994);
   assign  _net_7470 = (in_do&_net_3994);
   assign  _net_7471 = (in_do&_net_3994);
   assign  _net_7472 = (in_do&_net_3994);
   assign  _net_7473 = (in_do&_net_3994);
   assign  _net_7474 = (in_do&_net_3994);
   assign  _net_7475 = (in_do&_net_3994);
   assign  _net_7476 = (in_do&_net_3994);
   assign  _net_7477 = (in_do&_net_3994);
   assign  _net_7478 = (in_do&_net_3994);
   assign  _net_7479 = (in_do&_net_3994);
   assign  _net_7480 = (in_do&_net_3994);
   assign  _net_7481 = (in_do&_net_3994);
   assign  _net_7482 = (in_do&_net_3994);
   assign  _net_7483 = (in_do&_net_3994);
   assign  _net_7484 = (in_do&_net_3994);
   assign  _net_7485 = (in_do&_net_3994);
   assign  _net_7486 = (in_do&_net_3994);
   assign  _net_7487 = (in_do&_net_3994);
   assign  _net_7488 = (in_do&_net_3994);
   assign  _net_7489 = (in_do&_net_3994);
   assign  _net_7490 = (in_do&_net_3994);
   assign  _net_7491 = (in_do&_net_3994);
   assign  _net_7492 = (in_do&_net_3994);
   assign  _net_7493 = (in_do&_net_3994);
   assign  _net_7494 = (in_do&_net_3994);
   assign  _net_7495 = (in_do&_net_3994);
   assign  _net_7496 = (in_do&_net_3994);
   assign  _net_7497 = (in_do&_net_3994);
   assign  _net_7498 = (in_do&_net_3994);
   assign  _net_7499 = (in_do&_net_3994);
   assign  _net_7500 = (in_do&_net_3994);
   assign  _net_7501 = (in_do&_net_3994);
   assign  _net_7502 = (in_do&_net_3994);
   assign  _net_7503 = (in_do&_net_3994);
   assign  _net_7504 = (in_do&_net_3994);
   assign  _net_7505 = (in_do&_net_3994);
   assign  _net_7506 = (in_do&_net_3994);
   assign  _net_7507 = (in_do&_net_3994);
   assign  _net_7508 = (in_do&_net_3994);
   assign  _net_7509 = (in_do&_net_3994);
   assign  _net_7510 = (in_do&_net_3994);
   assign  _net_7511 = (in_do&_net_3994);
   assign  _net_7512 = (in_do&_net_3994);
   assign  _net_7513 = (in_do&_net_3994);
   assign  _net_7514 = (in_do&_net_3994);
   assign  _net_7515 = (in_do&_net_3994);
   assign  _net_7516 = (in_do&_net_3994);
   assign  _net_7517 = (in_do&_net_3994);
   assign  _net_7518 = (in_do&_net_3994);
   assign  _net_7519 = (in_do&_net_3994);
   assign  _net_7520 = (in_do&_net_3994);
   assign  _net_7521 = (in_do&_net_3994);
   assign  _net_7522 = (in_do&_net_3994);
   assign  _net_7523 = (in_do&_net_3994);
   assign  _net_7524 = (in_do&_net_3994);
   assign  _net_7525 = (in_do&_net_3994);
   assign  _net_7526 = (in_do&_net_3994);
   assign  _net_7527 = (in_do&_net_3994);
   assign  _net_7528 = (in_do&_net_3994);
   assign  _net_7529 = (in_do&_net_3994);
   assign  _net_7530 = (in_do&_net_3994);
   assign  _net_7531 = (in_do&_net_3994);
   assign  _net_7532 = (in_do&_net_3994);
   assign  _net_7533 = (in_do&_net_3994);
   assign  _net_7534 = (in_do&_net_3994);
   assign  _net_7535 = (in_do&_net_3994);
   assign  _net_7536 = (in_do&_net_3994);
   assign  _net_7537 = (in_do&_net_3994);
   assign  _net_7538 = (in_do&_net_3994);
   assign  _net_7539 = (in_do&_net_3994);
   assign  _net_7540 = (in_do&_net_3994);
   assign  _net_7541 = (in_do&_net_3994);
   assign  _net_7542 = (in_do&_net_3994);
   assign  _net_7543 = (in_do&_net_3994);
   assign  _net_7544 = (in_do&_net_3994);
   assign  _net_7545 = (in_do&_net_3994);
   assign  _net_7546 = (in_do&_net_3994);
   assign  _net_7547 = (in_do&_net_3994);
   assign  _net_7548 = (in_do&_net_3994);
   assign  _net_7549 = (in_do&_net_3994);
   assign  _net_7550 = (in_do&_net_3994);
   assign  _net_7551 = (in_do&_net_3994);
   assign  _net_7552 = (in_do&_net_3994);
   assign  _net_7553 = (in_do&_net_3994);
   assign  _net_7554 = (in_do&_net_3994);
   assign  _net_7555 = (in_do&_net_3994);
   assign  _net_7556 = (in_do&_net_3994);
   assign  _net_7557 = (in_do&_net_3994);
   assign  _net_7558 = (in_do&_net_3994);
   assign  _net_7559 = (in_do&_net_3994);
   assign  _net_7560 = (in_do&_net_3994);
   assign  _net_7561 = (in_do&_net_3994);
   assign  _net_7562 = (in_do&_net_3994);
   assign  _net_7563 = (in_do&_net_3994);
   assign  _net_7564 = (in_do&_net_3994);
   assign  _net_7565 = (in_do&_net_3994);
   assign  _net_7566 = (in_do&_net_3994);
   assign  _net_7567 = (in_do&_net_3994);
   assign  _net_7568 = (in_do&_net_3994);
   assign  _net_7569 = (in_do&_net_3994);
   assign  _net_7570 = (in_do&_net_3994);
   assign  _net_7571 = (in_do&_net_3994);
   assign  _net_7572 = (in_do&_net_3994);
   assign  _net_7573 = (in_do&_net_3994);
   assign  _net_7574 = (in_do&_net_3994);
   assign  _net_7575 = (in_do&_net_3994);
   assign  _net_7576 = (in_do&_net_3994);
   assign  _net_7577 = (in_do&_net_3994);
   assign  _net_7578 = (in_do&_net_3994);
   assign  _net_7579 = (in_do&_net_3994);
   assign  _net_7580 = (in_do&_net_3994);
   assign  _net_7581 = (in_do&_net_3994);
   assign  _net_7582 = (in_do&_net_3994);
   assign  _net_7583 = (in_do&_net_3994);
   assign  _net_7584 = (in_do&_net_3994);
   assign  _net_7585 = (in_do&_net_3994);
   assign  _net_7586 = (in_do&_net_3994);
   assign  _net_7587 = (in_do&_net_3994);
   assign  _net_7588 = (in_do&_net_3994);
   assign  _net_7589 = (in_do&_net_3994);
   assign  _net_7590 = (in_do&_net_3994);
   assign  _net_7591 = (in_do&_net_3994);
   assign  _net_7592 = (in_do&_net_3994);
   assign  _net_7593 = (in_do&_net_3994);
   assign  _net_7594 = (in_do&_net_3994);
   assign  _net_7595 = (in_do&_net_3994);
   assign  _net_7596 = (in_do&_net_3994);
   assign  _net_7597 = (in_do&_net_3994);
   assign  _net_7598 = (in_do&_net_3994);
   assign  _net_7599 = (in_do&_net_3994);
   assign  _net_7600 = (in_do&_net_3994);
   assign  _net_7601 = (in_do&_net_3994);
   assign  _net_7602 = (in_do&_net_3994);
   assign  _net_7603 = (in_do&_net_3994);
   assign  _net_7604 = (in_do&_net_3994);
   assign  _net_7605 = (in_do&_net_3994);
   assign  _net_7606 = (in_do&_net_3994);
   assign  _net_7607 = (in_do&_net_3994);
   assign  _net_7608 = (in_do&_net_3994);
   assign  _net_7609 = (in_do&_net_3994);
   assign  _net_7610 = (in_do&_net_3994);
   assign  _net_7611 = (in_do&_net_3994);
   assign  _net_7612 = (in_do&_net_3994);
   assign  _net_7613 = (in_do&_net_3994);
   assign  _net_7614 = (in_do&_net_3994);
   assign  _net_7615 = (in_do&_net_3994);
   assign  _net_7616 = (in_do&_net_3994);
   assign  _net_7617 = (in_do&_net_3994);
   assign  _net_7618 = (in_do&_net_3994);
   assign  _net_7619 = (in_do&_net_3994);
   assign  _net_7620 = (in_do&_net_3994);
   assign  _net_7621 = (in_do&_net_3994);
   assign  _net_7622 = (in_do&_net_3994);
   assign  _net_7623 = (in_do&_net_3994);
   assign  _net_7624 = (in_do&_net_3994);
   assign  _net_7625 = (in_do&_net_3994);
   assign  _net_7626 = (in_do&_net_3994);
   assign  _net_7627 = (in_do&_net_3994);
   assign  _net_7628 = (in_do&_net_3994);
   assign  _net_7629 = (in_do&_net_3994);
   assign  _net_7630 = (in_do&_net_3994);
   assign  _net_7631 = (in_do&_net_3994);
   assign  _net_7632 = (in_do&_net_3994);
   assign  _net_7633 = (in_do&_net_3994);
   assign  _net_7634 = (in_do&_net_3994);
   assign  _net_7635 = (in_do&_net_3994);
   assign  _net_7636 = (in_do&_net_3994);
   assign  _net_7637 = (in_do&_net_3994);
   assign  _net_7638 = (in_do&_net_3994);
   assign  _net_7639 = (in_do&_net_3994);
   assign  _net_7640 = (in_do&_net_3994);
   assign  _net_7641 = (in_do&_net_3994);
   assign  _net_7642 = (in_do&_net_3994);
   assign  _net_7643 = (in_do&_net_3994);
   assign  _net_7644 = (in_do&_net_3994);
   assign  _net_7645 = (in_do&_net_3994);
   assign  _net_7646 = (in_do&_net_3994);
   assign  _net_7647 = (in_do&_net_3994);
   assign  _net_7648 = (in_do&_net_3994);
   assign  _net_7649 = (in_do&_net_3994);
   assign  _net_7650 = (in_do&_net_3994);
   assign  _net_7651 = (in_do&_net_3994);
   assign  _net_7652 = (in_do&_net_3994);
   assign  _net_7653 = (in_do&_net_3994);
   assign  _net_7654 = (in_do&_net_3994);
   assign  _net_7655 = (in_do&_net_3994);
   assign  _net_7656 = (in_do&_net_3994);
   assign  _net_7657 = (in_do&_net_3994);
   assign  _net_7658 = (in_do&_net_3994);
   assign  _net_7659 = (in_do&_net_3994);
   assign  _net_7660 = (in_do&_net_3994);
   assign  _net_7661 = (in_do&_net_3994);
   assign  _net_7662 = (in_do&_net_3994);
   assign  _net_7663 = (in_do&_net_3994);
   assign  _net_7664 = (in_do&_net_3994);
   assign  _net_7665 = (in_do&_net_3994);
   assign  _net_7666 = (in_do&_net_3994);
   assign  _net_7667 = (in_do&_net_3994);
   assign  _net_7668 = (in_do&_net_3994);
   assign  _net_7669 = (in_do&_net_3994);
   assign  _net_7670 = (in_do&_net_3994);
   assign  _net_7671 = (in_do&_net_3994);
   assign  _net_7672 = (in_do&_net_3994);
   assign  _net_7673 = (in_do&_net_3994);
   assign  _net_7674 = (in_do&_net_3994);
   assign  _net_7675 = (in_do&_net_3994);
   assign  _net_7676 = (in_do&_net_3994);
   assign  _net_7677 = (in_do&_net_3994);
   assign  _net_7678 = (in_do&_net_3994);
   assign  _net_7679 = (in_do&_net_3994);
   assign  _net_7680 = (in_do&_net_3994);
   assign  _net_7681 = (in_do&_net_3994);
   assign  _net_7682 = (in_do&_net_3994);
   assign  _net_7683 = (in_do&_net_3994);
   assign  _net_7684 = (in_do&_net_3994);
   assign  _net_7685 = (in_do&_net_3994);
   assign  _net_7686 = (in_do&_net_3994);
   assign  _net_7687 = (in_do&_net_3994);
   assign  _net_7688 = (in_do&_net_3994);
   assign  _net_7689 = (in_do&_net_3994);
   assign  _net_7690 = (in_do&_net_3994);
   assign  _net_7691 = (in_do&_net_3994);
   assign  _net_7692 = (in_do&_net_3994);
   assign  _net_7693 = (in_do&_net_3994);
   assign  _net_7694 = (in_do&_net_3994);
   assign  _net_7695 = (in_do&_net_3994);
   assign  _net_7696 = (in_do&_net_3994);
   assign  _net_7697 = (in_do&_net_3994);
   assign  _net_7698 = (in_do&_net_3994);
   assign  _net_7699 = (in_do&_net_3994);
   assign  _net_7700 = (in_do&_net_3994);
   assign  _net_7701 = (in_do&_net_3994);
   assign  _net_7702 = (in_do&_net_3994);
   assign  _net_7703 = (in_do&_net_3994);
   assign  _net_7704 = (in_do&_net_3994);
   assign  _net_7705 = (in_do&_net_3994);
   assign  _net_7706 = (in_do&_net_3994);
   assign  _net_7707 = (in_do&_net_3994);
   assign  _net_7708 = (in_do&_net_3994);
   assign  _net_7709 = (in_do&_net_3994);
   assign  _net_7710 = (in_do&_net_3994);
   assign  _net_7711 = (in_do&_net_3994);
   assign  _net_7712 = (in_do&_net_3994);
   assign  _net_7713 = (in_do&_net_3994);
   assign  _net_7714 = (in_do&_net_3994);
   assign  _net_7715 = (in_do&_net_3994);
   assign  _net_7716 = (in_do&_net_3994);
   assign  _net_7717 = (in_do&_net_3994);
   assign  _net_7718 = (in_do&_net_3994);
   assign  _net_7719 = (in_do&_net_3994);
   assign  _net_7720 = (in_do&_net_3994);
   assign  _net_7721 = (in_do&_net_3994);
   assign  _net_7722 = (in_do&_net_3994);
   assign  _net_7723 = (in_do&_net_3994);
   assign  _net_7724 = (in_do&_net_3994);
   assign  _net_7725 = (in_do&_net_3994);
   assign  _net_7726 = (in_do&_net_3994);
   assign  _net_7727 = (in_do&_net_3994);
   assign  _net_7728 = (in_do&_net_3994);
   assign  _net_7729 = (in_do&_net_3994);
   assign  _net_7730 = (in_do&_net_3994);
   assign  _net_7731 = (in_do&_net_3994);
   assign  _net_7732 = (in_do&_net_3994);
   assign  _net_7733 = (in_do&_net_3994);
   assign  _net_7734 = (in_do&_net_3994);
   assign  _net_7735 = (in_do&_net_3994);
   assign  _net_7736 = (in_do&_net_3994);
   assign  _net_7737 = (in_do&_net_3994);
   assign  _net_7738 = (in_do&_net_3994);
   assign  _net_7739 = (in_do&_net_3994);
   assign  _net_7740 = (in_do&_net_3994);
   assign  _net_7741 = (in_do&_net_3994);
   assign  _net_7742 = (in_do&_net_3994);
   assign  _net_7743 = (in_do&_net_3994);
   assign  _net_7744 = (in_do&_net_3994);
   assign  _net_7745 = (in_do&_net_3994);
   assign  _net_7746 = (in_do&_net_3994);
   assign  _net_7747 = (in_do&_net_3994);
   assign  _net_7748 = (in_do&_net_3994);
   assign  _net_7749 = (in_do&_net_3994);
   assign  _net_7750 = (in_do&_net_3994);
   assign  _net_7751 = (in_do&_net_3994);
   assign  _net_7752 = (in_do&_net_3994);
   assign  _net_7753 = (in_do&_net_3994);
   assign  _net_7754 = (in_do&_net_3994);
   assign  _net_7755 = (in_do&_net_3994);
   assign  _net_7756 = (in_do&_net_3994);
   assign  _net_7757 = (in_do&_net_3994);
   assign  _net_7758 = (in_do&_net_3994);
   assign  _net_7759 = (in_do&_net_3994);
   assign  _net_7760 = (in_do&_net_3994);
   assign  _net_7761 = (in_do&_net_3994);
   assign  _net_7762 = (in_do&_net_3994);
   assign  _net_7763 = (in_do&_net_3994);
   assign  _net_7764 = (in_do&_net_3994);
   assign  _net_7765 = (in_do&_net_3994);
   assign  _net_7766 = (in_do&_net_3994);
   assign  _net_7767 = (in_do&_net_3994);
   assign  _net_7768 = (in_do&_net_3994);
   assign  _net_7769 = (in_do&_net_3994);
   assign  _net_7770 = (in_do&_net_3994);
   assign  _net_7771 = (in_do&_net_3994);
   assign  _net_7772 = (in_do&_net_3994);
   assign  _net_7773 = (in_do&_net_3994);
   assign  _net_7774 = (in_do&_net_3994);
   assign  _net_7775 = (in_do&_net_3994);
   assign  _net_7776 = (in_do&_net_3994);
   assign  _net_7777 = (in_do&_net_3994);
   assign  _net_7778 = (in_do&_net_3994);
   assign  _net_7779 = (in_do&_net_3994);
   assign  _net_7780 = (in_do&_net_3994);
   assign  _net_7781 = (in_do&_net_3994);
   assign  _net_7782 = (in_do&_net_3994);
   assign  _net_7783 = (in_do&_net_3994);
   assign  _net_7784 = (in_do&_net_3994);
   assign  _net_7785 = (in_do&_net_3994);
   assign  _net_7786 = (in_do&_net_3994);
   assign  _net_7787 = (in_do&_net_3994);
   assign  _net_7788 = (in_do&_net_3994);
   assign  _net_7789 = (in_do&_net_3994);
   assign  _net_7790 = (in_do&_net_3994);
   assign  _net_7791 = (in_do&_net_3994);
   assign  _net_7792 = (in_do&_net_3994);
   assign  _net_7793 = (in_do&_net_3994);
   assign  _net_7794 = (in_do&_net_3994);
   assign  _net_7795 = (in_do&_net_3994);
   assign  _net_7796 = (in_do&_net_3994);
   assign  _net_7797 = (in_do&_net_3994);
   assign  _net_7798 = (in_do&_net_3994);
   assign  _net_7799 = (in_do&_net_3994);
   assign  _net_7800 = (in_do&_net_3994);
   assign  _net_7801 = (in_do&_net_3994);
   assign  _net_7802 = (in_do&_net_3994);
   assign  _net_7803 = (in_do&_net_3994);
   assign  _net_7804 = (in_do&_net_3994);
   assign  _net_7805 = (in_do&_net_3994);
   assign  _net_7806 = (in_do&_net_3994);
   assign  _net_7807 = (in_do&_net_3994);
   assign  _net_7808 = (in_do&_net_3994);
   assign  _net_7809 = (in_do&_net_3994);
   assign  _net_7810 = (in_do&_net_3994);
   assign  _net_7811 = (in_do&_net_3994);
   assign  _net_7812 = (in_do&_net_3994);
   assign  _net_7813 = (in_do&_net_3994);
   assign  _net_7814 = (in_do&_net_3994);
   assign  _net_7815 = (in_do&_net_3994);
   assign  _net_7816 = (in_do&_net_3994);
   assign  _net_7817 = (in_do&_net_3994);
   assign  _net_7818 = (in_do&_net_3994);
   assign  _net_7819 = (in_do&_net_3994);
   assign  _net_7820 = (in_do&_net_3994);
   assign  _net_7821 = (in_do&_net_3994);
   assign  _net_7822 = (in_do&_net_3994);
   assign  _net_7823 = (in_do&_net_3994);
   assign  _net_7824 = (in_do&_net_3994);
   assign  _net_7825 = (in_do&_net_3994);
   assign  _net_7826 = (in_do&_net_3994);
   assign  _net_7827 = (in_do&_net_3994);
   assign  _net_7828 = (in_do&_net_3994);
   assign  _net_7829 = (in_do&_net_3994);
   assign  _net_7830 = (in_do&_net_3994);
   assign  _net_7831 = (in_do&_net_3994);
   assign  _net_7832 = (in_do&_net_3994);
   assign  _net_7833 = (in_do&_net_3994);
   assign  _net_7834 = (in_do&_net_3994);
   assign  _net_7835 = (in_do&_net_3994);
   assign  _net_7836 = (in_do&_net_3994);
   assign  _net_7837 = (in_do&_net_3994);
   assign  _net_7838 = (in_do&_net_3994);
   assign  _net_7839 = (in_do&_net_3994);
   assign  _net_7840 = (in_do&_net_3994);
   assign  _net_7841 = (in_do&_net_3994);
   assign  _net_7842 = (in_do&_net_3994);
   assign  _net_7843 = (in_do&_net_3994);
   assign  _net_7844 = (in_do&_net_3994);
   assign  _net_7845 = (in_do&_net_3994);
   assign  _net_7846 = (in_do&_net_3994);
   assign  _net_7847 = (in_do&_net_3994);
   assign  _net_7848 = (in_do&_net_3994);
   assign  _net_7849 = (in_do&_net_3994);
   assign  _net_7850 = (in_do&_net_3994);
   assign  _net_7851 = (in_do&_net_3994);
   assign  _net_7852 = (in_do&_net_3994);
   assign  _net_7853 = (in_do&_net_3994);
   assign  _net_7854 = (in_do&_net_3994);
   assign  _net_7855 = (in_do&_net_3994);
   assign  _net_7856 = (in_do&_net_3994);
   assign  _net_7857 = (in_do&_net_3994);
   assign  _net_7858 = (in_do&_net_3994);
   assign  _net_7859 = (in_do&_net_3994);
   assign  _net_7860 = (in_do&_net_3994);
   assign  _net_7861 = (in_do&_net_3994);
   assign  _net_7862 = (in_do&_net_3994);
   assign  _net_7863 = (in_do&_net_3994);
   assign  _net_7864 = (in_do&_net_3994);
   assign  _net_7865 = (in_do&_net_3994);
   assign  _net_7866 = (in_do&_net_3994);
   assign  _net_7867 = (in_do&_net_3994);
   assign  _net_7868 = (in_do&_net_3994);
   assign  _net_7869 = (in_do&_net_3994);
   assign  _net_7870 = (in_do&_net_3994);
   assign  _net_7871 = (in_do&_net_3994);
   assign  _net_7872 = (in_do&_net_3994);
   assign  _net_7873 = (in_do&_net_3994);
   assign  _net_7874 = (in_do&_net_3994);
   assign  _net_7875 = (in_do&_net_3994);
   assign  _net_7876 = (in_do&_net_3994);
   assign  _net_7877 = (in_do&_net_3994);
   assign  _net_7878 = (in_do&_net_3994);
   assign  _net_7879 = (in_do&_net_3994);
   assign  _net_7880 = (in_do&_net_3994);
   assign  _net_7881 = (in_do&_net_3994);
   assign  _net_7882 = (in_do&_net_3994);
   assign  _net_7883 = (in_do&_net_3994);
   assign  _net_7884 = (in_do&_net_3994);
   assign  _net_7885 = (in_do&_net_3994);
   assign  _net_7886 = (in_do&_net_3994);
   assign  _net_7887 = (in_do&_net_3994);
   assign  _net_7888 = (in_do&_net_3994);
   assign  _net_7889 = (in_do&_net_3994);
   assign  _net_7890 = (in_do&_net_3994);
   assign  _net_7891 = (in_do&_net_3994);
   assign  _net_7892 = (in_do&_net_3994);
   assign  _net_7893 = (in_do&_net_3994);
   assign  _net_7894 = (in_do&_net_3994);
   assign  _net_7895 = (in_do&_net_3994);
   assign  _net_7896 = (in_do&_net_3994);
   assign  _net_7897 = (in_do&_net_3994);
   assign  _net_7898 = (in_do&_net_3994);
   assign  _net_7899 = (in_do&_net_3994);
   assign  _net_7900 = (in_do&_net_3994);
   assign  _net_7901 = (in_do&_net_3994);
   assign  _net_7902 = (in_do&_net_3994);
   assign  _net_7903 = (in_do&_net_3994);
   assign  _net_7904 = (in_do&_net_3994);
   assign  _net_7905 = (in_do&_net_3994);
   assign  _net_7906 = (in_do&_net_3994);
   assign  _net_7907 = (in_do&_net_3994);
   assign  _net_7908 = (in_do&_net_3994);
   assign  _net_7909 = (in_do&_net_3994);
   assign  _net_7910 = (in_do&_net_3994);
   assign  _net_7911 = (in_do&_net_3994);
   assign  _net_7912 = (in_do&_net_3994);
   assign  _net_7913 = (in_do&_net_3994);
   assign  _net_7914 = (in_do&_net_3994);
   assign  _net_7915 = (in_do&_net_3994);
   assign  _net_7916 = (in_do&_net_3994);
   assign  _net_7917 = (in_do&_net_3994);
   assign  _net_7918 = (in_do&_net_3994);
   assign  _net_7919 = (in_do&_net_3994);
   assign  _net_7920 = (in_do&_net_3994);
   assign  _net_7921 = (in_do&_net_3994);
   assign  _net_7922 = (in_do&_net_3994);
   assign  _net_7923 = (in_do&_net_3994);
   assign  _net_7924 = (in_do&_net_3994);
   assign  _net_7925 = (in_do&_net_3994);
   assign  _net_7926 = (in_do&_net_3994);
   assign  _net_7927 = (in_do&_net_3994);
   assign  _net_7928 = (in_do&_net_3994);
   assign  _net_7929 = (in_do&_net_3994);
   assign  _net_7930 = (in_do&_net_3994);
   assign  _net_7931 = (in_do&_net_3994);
   assign  _net_7932 = (in_do&_net_3994);
   assign  _net_7933 = (in_do&_net_3994);
   assign  _net_7934 = (in_do&_net_3994);
   assign  _net_7935 = (in_do&_net_3994);
   assign  _net_7936 = (in_do&_net_3994);
   assign  _net_7937 = (in_do&_net_3994);
   assign  _net_7938 = (in_do&_net_3994);
   assign  _net_7939 = (in_do&_net_3994);
   assign  _net_7940 = (in_do&_net_3994);
   assign  _net_7941 = (in_do&_net_3994);
   assign  _net_7942 = (in_do&_net_3994);
   assign  _net_7943 = (in_do&_net_3994);
   assign  _net_7944 = (in_do&_net_3994);
   assign  _net_7945 = (in_do&_net_3994);
   assign  _net_7946 = (in_do&_net_3994);
   assign  _net_7947 = (in_do&_net_3994);
   assign  _net_7948 = (in_do&_net_3994);
   assign  _net_7949 = (in_do&_net_3994);
   assign  _net_7950 = (in_do&_net_3994);
   assign  _net_7951 = (in_do&_net_3994);
   assign  _net_7952 = (in_do&_net_3994);
   assign  _net_7953 = (in_do&_net_3994);
   assign  _net_7954 = (in_do&_net_3994);
   assign  _net_7955 = (in_do&_net_3994);
   assign  _net_7956 = (in_do&_net_3994);
   assign  _net_7957 = (in_do&_net_3994);
   assign  _net_7958 = (in_do&_net_3994);
   assign  _net_7959 = (in_do&_net_3994);
   assign  _net_7960 = (in_do&_net_3994);
   assign  _net_7961 = (in_do&_net_3994);
   assign  _net_7962 = (in_do&_net_3994);
   assign  _net_7963 = (in_do&_net_3994);
   assign  _net_7964 = (in_do&_net_3994);
   assign  _net_7965 = (in_do&_net_3994);
   assign  _net_7966 = (in_do&_net_3994);
   assign  _net_7967 = (in_do&_net_3994);
   assign  _net_7968 = (in_do&_net_3994);
   assign  _net_7969 = (in_do&_net_3994);
   assign  _net_7970 = (in_do&_net_3994);
   assign  _net_7971 = (in_do&_net_3994);
   assign  _net_7972 = (in_do&_net_3994);
   assign  _net_7973 = (in_do&_net_3994);
   assign  _net_7974 = (in_do&_net_3994);
   assign  _net_7975 = (in_do&_net_3994);
   assign  _net_7976 = (in_do&_net_3994);
   assign  _net_7977 = (in_do&_net_3994);
   assign  _net_7978 = (in_do&_net_3994);
   assign  _net_7979 = (in_do&_net_3994);
   assign  _net_7980 = (in_do&_net_3994);
   assign  _net_7981 = (in_do&_net_3994);
   assign  _net_7982 = (in_do&_net_3994);
   assign  _net_7983 = (in_do&_net_3994);
   assign  _net_7984 = (in_do&_net_3994);
   assign  _net_7985 = (in_do&_net_3994);
   assign  data_out_org33 = ((_net_1)?_add_map_x_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_data_org:10'b0);
   assign  data_out_org34 = ((_net_1)?_add_map_x_data_org:10'b0)|
    ((_net_0)?_add_map_x_data_org_near:10'b0);
   assign  data_out_org35 = ((_net_1)?_add_map_x_1_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_1_data_org:10'b0);
   assign  data_out_org36 = ((_net_1)?_add_map_x_1_data_org:10'b0)|
    ((_net_0)?_add_map_x_1_data_org_near:10'b0);
   assign  data_out_org37 = ((_net_1)?_add_map_x_2_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_2_data_org:10'b0);
   assign  data_out_org38 = ((_net_1)?_add_map_x_2_data_org:10'b0)|
    ((_net_0)?_add_map_x_2_data_org_near:10'b0);
   assign  data_out_org39 = ((_net_1)?_add_map_x_3_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_3_data_org:10'b0);
   assign  data_out_org40 = ((_net_1)?_add_map_x_3_data_org:10'b0)|
    ((_net_0)?_add_map_x_3_data_org_near:10'b0);
   assign  data_out_org41 = ((_net_1)?_add_map_x_4_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_4_data_org:10'b0);
   assign  data_out_org42 = ((_net_1)?_add_map_x_4_data_org:10'b0)|
    ((_net_0)?_add_map_x_4_data_org_near:10'b0);
   assign  data_out_org43 = ((_net_1)?_add_map_x_5_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_5_data_org:10'b0);
   assign  data_out_org44 = ((_net_1)?_add_map_x_5_data_org:10'b0)|
    ((_net_0)?_add_map_x_5_data_org_near:10'b0);
   assign  data_out_org45 = ((_net_1)?_add_map_x_6_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_6_data_org:10'b0);
   assign  data_out_org46 = ((_net_1)?_add_map_x_6_data_org:10'b0)|
    ((_net_0)?_add_map_x_6_data_org_near:10'b0);
   assign  data_out_org47 = ((_net_1)?_add_map_x_7_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_7_data_org:10'b0);
   assign  data_out_org48 = ((_net_1)?_add_map_x_7_data_org:10'b0)|
    ((_net_0)?_add_map_x_7_data_org_near:10'b0);
   assign  data_out_org49 = ((_net_1)?_add_map_x_8_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_8_data_org:10'b0);
   assign  data_out_org50 = ((_net_1)?_add_map_x_8_data_org:10'b0)|
    ((_net_0)?_add_map_x_8_data_org_near:10'b0);
   assign  data_out_org51 = ((_net_1)?_add_map_x_9_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_9_data_org:10'b0);
   assign  data_out_org52 = ((_net_1)?_add_map_x_9_data_org:10'b0)|
    ((_net_0)?_add_map_x_9_data_org_near:10'b0);
   assign  data_out_org53 = ((_net_1)?_add_map_x_10_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_10_data_org:10'b0);
   assign  data_out_org54 = ((_net_1)?_add_map_x_10_data_org:10'b0)|
    ((_net_0)?_add_map_x_10_data_org_near:10'b0);
   assign  data_out_org55 = ((_net_1)?_add_map_x_11_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_11_data_org:10'b0);
   assign  data_out_org56 = ((_net_1)?_add_map_x_11_data_org:10'b0)|
    ((_net_0)?_add_map_x_11_data_org_near:10'b0);
   assign  data_out_org57 = ((_net_1)?_add_map_x_12_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_12_data_org:10'b0);
   assign  data_out_org58 = ((_net_1)?_add_map_x_12_data_org:10'b0)|
    ((_net_0)?_add_map_x_12_data_org_near:10'b0);
   assign  data_out_org59 = ((_net_1)?_add_map_x_13_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_13_data_org:10'b0);
   assign  data_out_org60 = ((_net_1)?_add_map_x_13_data_org:10'b0)|
    ((_net_0)?_add_map_x_13_data_org_near:10'b0);
   assign  data_out_org61 = ((_net_1)?_add_map_x_14_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_14_data_org:10'b0);
   assign  data_out_org62 = ((_net_1)?_add_map_x_14_data_org:10'b0)|
    ((_net_0)?_add_map_x_14_data_org_near:10'b0);
   assign  data_out_org65 = ((_net_1)?_add_map_x_15_data_org:10'b0)|
    ((_net_0)?_add_map_x_15_data_org_near:10'b0);
   assign  data_out_org66 = ((_net_1)?_add_map_x_15_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_15_data_org:10'b0);
   assign  data_out_org67 = ((_net_1)?_add_map_x_16_data_org:10'b0)|
    ((_net_0)?_add_map_x_16_data_org_near:10'b0);
   assign  data_out_org68 = ((_net_1)?_add_map_x_16_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_16_data_org:10'b0);
   assign  data_out_org69 = ((_net_1)?_add_map_x_17_data_org:10'b0)|
    ((_net_0)?_add_map_x_17_data_org_near:10'b0);
   assign  data_out_org70 = ((_net_1)?_add_map_x_17_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_17_data_org:10'b0);
   assign  data_out_org71 = ((_net_1)?_add_map_x_18_data_org:10'b0)|
    ((_net_0)?_add_map_x_18_data_org_near:10'b0);
   assign  data_out_org72 = ((_net_1)?_add_map_x_18_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_18_data_org:10'b0);
   assign  data_out_org73 = ((_net_1)?_add_map_x_19_data_org:10'b0)|
    ((_net_0)?_add_map_x_19_data_org_near:10'b0);
   assign  data_out_org74 = ((_net_1)?_add_map_x_19_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_19_data_org:10'b0);
   assign  data_out_org75 = ((_net_1)?_add_map_x_20_data_org:10'b0)|
    ((_net_0)?_add_map_x_20_data_org_near:10'b0);
   assign  data_out_org76 = ((_net_1)?_add_map_x_20_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_20_data_org:10'b0);
   assign  data_out_org77 = ((_net_1)?_add_map_x_21_data_org:10'b0)|
    ((_net_0)?_add_map_x_21_data_org_near:10'b0);
   assign  data_out_org78 = ((_net_1)?_add_map_x_21_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_21_data_org:10'b0);
   assign  data_out_org79 = ((_net_1)?_add_map_x_22_data_org:10'b0)|
    ((_net_0)?_add_map_x_22_data_org_near:10'b0);
   assign  data_out_org80 = ((_net_1)?_add_map_x_22_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_22_data_org:10'b0);
   assign  data_out_org81 = ((_net_1)?_add_map_x_23_data_org:10'b0)|
    ((_net_0)?_add_map_x_23_data_org_near:10'b0);
   assign  data_out_org82 = ((_net_1)?_add_map_x_23_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_23_data_org:10'b0);
   assign  data_out_org83 = ((_net_1)?_add_map_x_24_data_org:10'b0)|
    ((_net_0)?_add_map_x_24_data_org_near:10'b0);
   assign  data_out_org84 = ((_net_1)?_add_map_x_24_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_24_data_org:10'b0);
   assign  data_out_org85 = ((_net_1)?_add_map_x_25_data_org:10'b0)|
    ((_net_0)?_add_map_x_25_data_org_near:10'b0);
   assign  data_out_org86 = ((_net_1)?_add_map_x_25_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_25_data_org:10'b0);
   assign  data_out_org87 = ((_net_1)?_add_map_x_26_data_org:10'b0)|
    ((_net_0)?_add_map_x_26_data_org_near:10'b0);
   assign  data_out_org88 = ((_net_1)?_add_map_x_26_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_26_data_org:10'b0);
   assign  data_out_org89 = ((_net_1)?_add_map_x_27_data_org:10'b0)|
    ((_net_0)?_add_map_x_27_data_org_near:10'b0);
   assign  data_out_org90 = ((_net_1)?_add_map_x_27_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_27_data_org:10'b0);
   assign  data_out_org91 = ((_net_1)?_add_map_x_28_data_org:10'b0)|
    ((_net_0)?_add_map_x_28_data_org_near:10'b0);
   assign  data_out_org92 = ((_net_1)?_add_map_x_28_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_28_data_org:10'b0);
   assign  data_out_org93 = ((_net_1)?_add_map_x_29_data_org:10'b0)|
    ((_net_0)?_add_map_x_29_data_org_near:10'b0);
   assign  data_out_org94 = ((_net_1)?_add_map_x_29_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_29_data_org:10'b0);
   assign  data_out_org97 = ((_net_1)?_add_map_x_30_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_30_data_org:10'b0);
   assign  data_out_org98 = ((_net_1)?_add_map_x_30_data_org:10'b0)|
    ((_net_0)?_add_map_x_30_data_org_near:10'b0);
   assign  data_out_org99 = ((_net_1)?_add_map_x_31_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_31_data_org:10'b0);
   assign  data_out_org100 = ((_net_1)?_add_map_x_31_data_org:10'b0)|
    ((_net_0)?_add_map_x_31_data_org_near:10'b0);
   assign  data_out_org101 = ((_net_1)?_add_map_x_32_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_32_data_org:10'b0);
   assign  data_out_org102 = ((_net_1)?_add_map_x_32_data_org:10'b0)|
    ((_net_0)?_add_map_x_32_data_org_near:10'b0);
   assign  data_out_org103 = ((_net_1)?_add_map_x_33_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_33_data_org:10'b0);
   assign  data_out_org104 = ((_net_1)?_add_map_x_33_data_org:10'b0)|
    ((_net_0)?_add_map_x_33_data_org_near:10'b0);
   assign  data_out_org105 = ((_net_1)?_add_map_x_34_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_34_data_org:10'b0);
   assign  data_out_org106 = ((_net_1)?_add_map_x_34_data_org:10'b0)|
    ((_net_0)?_add_map_x_34_data_org_near:10'b0);
   assign  data_out_org107 = ((_net_1)?_add_map_x_35_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_35_data_org:10'b0);
   assign  data_out_org108 = ((_net_1)?_add_map_x_35_data_org:10'b0)|
    ((_net_0)?_add_map_x_35_data_org_near:10'b0);
   assign  data_out_org109 = ((_net_1)?_add_map_x_36_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_36_data_org:10'b0);
   assign  data_out_org110 = ((_net_1)?_add_map_x_36_data_org:10'b0)|
    ((_net_0)?_add_map_x_36_data_org_near:10'b0);
   assign  data_out_org111 = ((_net_1)?_add_map_x_37_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_37_data_org:10'b0);
   assign  data_out_org112 = ((_net_1)?_add_map_x_37_data_org:10'b0)|
    ((_net_0)?_add_map_x_37_data_org_near:10'b0);
   assign  data_out_org113 = ((_net_1)?_add_map_x_38_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_38_data_org:10'b0);
   assign  data_out_org114 = ((_net_1)?_add_map_x_38_data_org:10'b0)|
    ((_net_0)?_add_map_x_38_data_org_near:10'b0);
   assign  data_out_org115 = ((_net_1)?_add_map_x_39_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_39_data_org:10'b0);
   assign  data_out_org116 = ((_net_1)?_add_map_x_39_data_org:10'b0)|
    ((_net_0)?_add_map_x_39_data_org_near:10'b0);
   assign  data_out_org117 = ((_net_1)?_add_map_x_40_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_40_data_org:10'b0);
   assign  data_out_org118 = ((_net_1)?_add_map_x_40_data_org:10'b0)|
    ((_net_0)?_add_map_x_40_data_org_near:10'b0);
   assign  data_out_org119 = ((_net_1)?_add_map_x_41_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_41_data_org:10'b0);
   assign  data_out_org120 = ((_net_1)?_add_map_x_41_data_org:10'b0)|
    ((_net_0)?_add_map_x_41_data_org_near:10'b0);
   assign  data_out_org121 = ((_net_1)?_add_map_x_42_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_42_data_org:10'b0);
   assign  data_out_org122 = ((_net_1)?_add_map_x_42_data_org:10'b0)|
    ((_net_0)?_add_map_x_42_data_org_near:10'b0);
   assign  data_out_org123 = ((_net_1)?_add_map_x_43_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_43_data_org:10'b0);
   assign  data_out_org124 = ((_net_1)?_add_map_x_43_data_org:10'b0)|
    ((_net_0)?_add_map_x_43_data_org_near:10'b0);
   assign  data_out_org125 = ((_net_1)?_add_map_x_44_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_44_data_org:10'b0);
   assign  data_out_org126 = ((_net_1)?_add_map_x_44_data_org:10'b0)|
    ((_net_0)?_add_map_x_44_data_org_near:10'b0);
   assign  data_out_org129 = ((_net_1)?_add_map_x_45_data_org:10'b0)|
    ((_net_0)?_add_map_x_45_data_org_near:10'b0);
   assign  data_out_org130 = ((_net_1)?_add_map_x_45_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_45_data_org:10'b0);
   assign  data_out_org131 = ((_net_1)?_add_map_x_46_data_org:10'b0)|
    ((_net_0)?_add_map_x_46_data_org_near:10'b0);
   assign  data_out_org132 = ((_net_1)?_add_map_x_46_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_46_data_org:10'b0);
   assign  data_out_org133 = ((_net_1)?_add_map_x_47_data_org:10'b0)|
    ((_net_0)?_add_map_x_47_data_org_near:10'b0);
   assign  data_out_org134 = ((_net_1)?_add_map_x_47_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_47_data_org:10'b0);
   assign  data_out_org135 = ((_net_1)?_add_map_x_48_data_org:10'b0)|
    ((_net_0)?_add_map_x_48_data_org_near:10'b0);
   assign  data_out_org136 = ((_net_1)?_add_map_x_48_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_48_data_org:10'b0);
   assign  data_out_org137 = ((_net_1)?_add_map_x_49_data_org:10'b0)|
    ((_net_0)?_add_map_x_49_data_org_near:10'b0);
   assign  data_out_org138 = ((_net_1)?_add_map_x_49_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_49_data_org:10'b0);
   assign  data_out_org139 = ((_net_1)?_add_map_x_50_data_org:10'b0)|
    ((_net_0)?_add_map_x_50_data_org_near:10'b0);
   assign  data_out_org140 = ((_net_1)?_add_map_x_50_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_50_data_org:10'b0);
   assign  data_out_org141 = ((_net_1)?_add_map_x_51_data_org:10'b0)|
    ((_net_0)?_add_map_x_51_data_org_near:10'b0);
   assign  data_out_org142 = ((_net_1)?_add_map_x_51_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_51_data_org:10'b0);
   assign  data_out_org143 = ((_net_1)?_add_map_x_52_data_org:10'b0)|
    ((_net_0)?_add_map_x_52_data_org_near:10'b0);
   assign  data_out_org144 = ((_net_1)?_add_map_x_52_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_52_data_org:10'b0);
   assign  data_out_org145 = ((_net_1)?_add_map_x_53_data_org:10'b0)|
    ((_net_0)?_add_map_x_53_data_org_near:10'b0);
   assign  data_out_org146 = ((_net_1)?_add_map_x_53_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_53_data_org:10'b0);
   assign  data_out_org147 = ((_net_1)?_add_map_x_54_data_org:10'b0)|
    ((_net_0)?_add_map_x_54_data_org_near:10'b0);
   assign  data_out_org148 = ((_net_1)?_add_map_x_54_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_54_data_org:10'b0);
   assign  data_out_org149 = ((_net_1)?_add_map_x_55_data_org:10'b0)|
    ((_net_0)?_add_map_x_55_data_org_near:10'b0);
   assign  data_out_org150 = ((_net_1)?_add_map_x_55_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_55_data_org:10'b0);
   assign  data_out_org151 = ((_net_1)?_add_map_x_56_data_org:10'b0)|
    ((_net_0)?_add_map_x_56_data_org_near:10'b0);
   assign  data_out_org152 = ((_net_1)?_add_map_x_56_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_56_data_org:10'b0);
   assign  data_out_org153 = ((_net_1)?_add_map_x_57_data_org:10'b0)|
    ((_net_0)?_add_map_x_57_data_org_near:10'b0);
   assign  data_out_org154 = ((_net_1)?_add_map_x_57_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_57_data_org:10'b0);
   assign  data_out_org155 = ((_net_1)?_add_map_x_58_data_org:10'b0)|
    ((_net_0)?_add_map_x_58_data_org_near:10'b0);
   assign  data_out_org156 = ((_net_1)?_add_map_x_58_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_58_data_org:10'b0);
   assign  data_out_org157 = ((_net_1)?_add_map_x_59_data_org:10'b0)|
    ((_net_0)?_add_map_x_59_data_org_near:10'b0);
   assign  data_out_org158 = ((_net_1)?_add_map_x_59_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_59_data_org:10'b0);
   assign  data_out_org161 = ((_net_1)?_add_map_x_60_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_60_data_org:10'b0);
   assign  data_out_org162 = ((_net_1)?_add_map_x_60_data_org:10'b0)|
    ((_net_0)?_add_map_x_60_data_org_near:10'b0);
   assign  data_out_org163 = ((_net_1)?_add_map_x_61_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_61_data_org:10'b0);
   assign  data_out_org164 = ((_net_1)?_add_map_x_61_data_org:10'b0)|
    ((_net_0)?_add_map_x_61_data_org_near:10'b0);
   assign  data_out_org165 = ((_net_1)?_add_map_x_62_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_62_data_org:10'b0);
   assign  data_out_org166 = ((_net_1)?_add_map_x_62_data_org:10'b0)|
    ((_net_0)?_add_map_x_62_data_org_near:10'b0);
   assign  data_out_org167 = ((_net_1)?_add_map_x_63_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_63_data_org:10'b0);
   assign  data_out_org168 = ((_net_1)?_add_map_x_63_data_org:10'b0)|
    ((_net_0)?_add_map_x_63_data_org_near:10'b0);
   assign  data_out_org169 = ((_net_1)?_add_map_x_64_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_64_data_org:10'b0);
   assign  data_out_org170 = ((_net_1)?_add_map_x_64_data_org:10'b0)|
    ((_net_0)?_add_map_x_64_data_org_near:10'b0);
   assign  data_out_org171 = ((_net_1)?_add_map_x_65_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_65_data_org:10'b0);
   assign  data_out_org172 = ((_net_1)?_add_map_x_65_data_org:10'b0)|
    ((_net_0)?_add_map_x_65_data_org_near:10'b0);
   assign  data_out_org173 = ((_net_1)?_add_map_x_66_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_66_data_org:10'b0);
   assign  data_out_org174 = ((_net_1)?_add_map_x_66_data_org:10'b0)|
    ((_net_0)?_add_map_x_66_data_org_near:10'b0);
   assign  data_out_org175 = ((_net_1)?_add_map_x_67_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_67_data_org:10'b0);
   assign  data_out_org176 = ((_net_1)?_add_map_x_67_data_org:10'b0)|
    ((_net_0)?_add_map_x_67_data_org_near:10'b0);
   assign  data_out_org177 = ((_net_1)?_add_map_x_68_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_68_data_org:10'b0);
   assign  data_out_org178 = ((_net_1)?_add_map_x_68_data_org:10'b0)|
    ((_net_0)?_add_map_x_68_data_org_near:10'b0);
   assign  data_out_org179 = ((_net_1)?_add_map_x_69_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_69_data_org:10'b0);
   assign  data_out_org180 = ((_net_1)?_add_map_x_69_data_org:10'b0)|
    ((_net_0)?_add_map_x_69_data_org_near:10'b0);
   assign  data_out_org181 = ((_net_1)?_add_map_x_70_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_70_data_org:10'b0);
   assign  data_out_org182 = ((_net_1)?_add_map_x_70_data_org:10'b0)|
    ((_net_0)?_add_map_x_70_data_org_near:10'b0);
   assign  data_out_org183 = ((_net_1)?_add_map_x_71_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_71_data_org:10'b0);
   assign  data_out_org184 = ((_net_1)?_add_map_x_71_data_org:10'b0)|
    ((_net_0)?_add_map_x_71_data_org_near:10'b0);
   assign  data_out_org185 = ((_net_1)?_add_map_x_72_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_72_data_org:10'b0);
   assign  data_out_org186 = ((_net_1)?_add_map_x_72_data_org:10'b0)|
    ((_net_0)?_add_map_x_72_data_org_near:10'b0);
   assign  data_out_org187 = ((_net_1)?_add_map_x_73_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_73_data_org:10'b0);
   assign  data_out_org188 = ((_net_1)?_add_map_x_73_data_org:10'b0)|
    ((_net_0)?_add_map_x_73_data_org_near:10'b0);
   assign  data_out_org189 = ((_net_1)?_add_map_x_74_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_74_data_org:10'b0);
   assign  data_out_org190 = ((_net_1)?_add_map_x_74_data_org:10'b0)|
    ((_net_0)?_add_map_x_74_data_org_near:10'b0);
   assign  data_out_org193 = ((_net_1)?_add_map_x_75_data_org:10'b0)|
    ((_net_0)?_add_map_x_75_data_org_near:10'b0);
   assign  data_out_org194 = ((_net_1)?_add_map_x_75_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_75_data_org:10'b0);
   assign  data_out_org195 = ((_net_1)?_add_map_x_76_data_org:10'b0)|
    ((_net_0)?_add_map_x_76_data_org_near:10'b0);
   assign  data_out_org196 = ((_net_1)?_add_map_x_76_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_76_data_org:10'b0);
   assign  data_out_org197 = ((_net_1)?_add_map_x_77_data_org:10'b0)|
    ((_net_0)?_add_map_x_77_data_org_near:10'b0);
   assign  data_out_org198 = ((_net_1)?_add_map_x_77_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_77_data_org:10'b0);
   assign  data_out_org199 = ((_net_1)?_add_map_x_78_data_org:10'b0)|
    ((_net_0)?_add_map_x_78_data_org_near:10'b0);
   assign  data_out_org200 = ((_net_1)?_add_map_x_78_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_78_data_org:10'b0);
   assign  data_out_org201 = ((_net_1)?_add_map_x_79_data_org:10'b0)|
    ((_net_0)?_add_map_x_79_data_org_near:10'b0);
   assign  data_out_org202 = ((_net_1)?_add_map_x_79_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_79_data_org:10'b0);
   assign  data_out_org203 = ((_net_1)?_add_map_x_80_data_org:10'b0)|
    ((_net_0)?_add_map_x_80_data_org_near:10'b0);
   assign  data_out_org204 = ((_net_1)?_add_map_x_80_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_80_data_org:10'b0);
   assign  data_out_org205 = ((_net_1)?_add_map_x_81_data_org:10'b0)|
    ((_net_0)?_add_map_x_81_data_org_near:10'b0);
   assign  data_out_org206 = ((_net_1)?_add_map_x_81_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_81_data_org:10'b0);
   assign  data_out_org207 = ((_net_1)?_add_map_x_82_data_org:10'b0)|
    ((_net_0)?_add_map_x_82_data_org_near:10'b0);
   assign  data_out_org208 = ((_net_1)?_add_map_x_82_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_82_data_org:10'b0);
   assign  data_out_org209 = ((_net_1)?_add_map_x_83_data_org:10'b0)|
    ((_net_0)?_add_map_x_83_data_org_near:10'b0);
   assign  data_out_org210 = ((_net_1)?_add_map_x_83_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_83_data_org:10'b0);
   assign  data_out_org211 = ((_net_1)?_add_map_x_84_data_org:10'b0)|
    ((_net_0)?_add_map_x_84_data_org_near:10'b0);
   assign  data_out_org212 = ((_net_1)?_add_map_x_84_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_84_data_org:10'b0);
   assign  data_out_org213 = ((_net_1)?_add_map_x_85_data_org:10'b0)|
    ((_net_0)?_add_map_x_85_data_org_near:10'b0);
   assign  data_out_org214 = ((_net_1)?_add_map_x_85_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_85_data_org:10'b0);
   assign  data_out_org215 = ((_net_1)?_add_map_x_86_data_org:10'b0)|
    ((_net_0)?_add_map_x_86_data_org_near:10'b0);
   assign  data_out_org216 = ((_net_1)?_add_map_x_86_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_86_data_org:10'b0);
   assign  data_out_org217 = ((_net_1)?_add_map_x_87_data_org:10'b0)|
    ((_net_0)?_add_map_x_87_data_org_near:10'b0);
   assign  data_out_org218 = ((_net_1)?_add_map_x_87_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_87_data_org:10'b0);
   assign  data_out_org219 = ((_net_1)?_add_map_x_88_data_org:10'b0)|
    ((_net_0)?_add_map_x_88_data_org_near:10'b0);
   assign  data_out_org220 = ((_net_1)?_add_map_x_88_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_88_data_org:10'b0);
   assign  data_out_org221 = ((_net_1)?_add_map_x_89_data_org:10'b0)|
    ((_net_0)?_add_map_x_89_data_org_near:10'b0);
   assign  data_out_org222 = ((_net_1)?_add_map_x_89_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_89_data_org:10'b0);
   assign  data_out_org225 = ((_net_1)?_add_map_x_90_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_90_data_org:10'b0);
   assign  data_out_org226 = ((_net_1)?_add_map_x_90_data_org:10'b0)|
    ((_net_0)?_add_map_x_90_data_org_near:10'b0);
   assign  data_out_org227 = ((_net_1)?_add_map_x_91_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_91_data_org:10'b0);
   assign  data_out_org228 = ((_net_1)?_add_map_x_91_data_org:10'b0)|
    ((_net_0)?_add_map_x_91_data_org_near:10'b0);
   assign  data_out_org229 = ((_net_1)?_add_map_x_92_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_92_data_org:10'b0);
   assign  data_out_org230 = ((_net_1)?_add_map_x_92_data_org:10'b0)|
    ((_net_0)?_add_map_x_92_data_org_near:10'b0);
   assign  data_out_org231 = ((_net_1)?_add_map_x_93_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_93_data_org:10'b0);
   assign  data_out_org232 = ((_net_1)?_add_map_x_93_data_org:10'b0)|
    ((_net_0)?_add_map_x_93_data_org_near:10'b0);
   assign  data_out_org233 = ((_net_1)?_add_map_x_94_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_94_data_org:10'b0);
   assign  data_out_org234 = ((_net_1)?_add_map_x_94_data_org:10'b0)|
    ((_net_0)?_add_map_x_94_data_org_near:10'b0);
   assign  data_out_org235 = ((_net_1)?_add_map_x_95_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_95_data_org:10'b0);
   assign  data_out_org236 = ((_net_1)?_add_map_x_95_data_org:10'b0)|
    ((_net_0)?_add_map_x_95_data_org_near:10'b0);
   assign  data_out_org237 = ((_net_1)?_add_map_x_96_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_96_data_org:10'b0);
   assign  data_out_org238 = ((_net_1)?_add_map_x_96_data_org:10'b0)|
    ((_net_0)?_add_map_x_96_data_org_near:10'b0);
   assign  data_out_org239 = ((_net_1)?_add_map_x_97_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_97_data_org:10'b0);
   assign  data_out_org240 = ((_net_1)?_add_map_x_97_data_org:10'b0)|
    ((_net_0)?_add_map_x_97_data_org_near:10'b0);
   assign  data_out_org241 = ((_net_1)?_add_map_x_98_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_98_data_org:10'b0);
   assign  data_out_org242 = ((_net_1)?_add_map_x_98_data_org:10'b0)|
    ((_net_0)?_add_map_x_98_data_org_near:10'b0);
   assign  data_out_org243 = ((_net_1)?_add_map_x_99_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_99_data_org:10'b0);
   assign  data_out_org244 = ((_net_1)?_add_map_x_99_data_org:10'b0)|
    ((_net_0)?_add_map_x_99_data_org_near:10'b0);
   assign  data_out_org245 = ((_net_1)?_add_map_x_100_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_100_data_org:10'b0);
   assign  data_out_org246 = ((_net_1)?_add_map_x_100_data_org:10'b0)|
    ((_net_0)?_add_map_x_100_data_org_near:10'b0);
   assign  data_out_org247 = ((_net_1)?_add_map_x_101_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_101_data_org:10'b0);
   assign  data_out_org248 = ((_net_1)?_add_map_x_101_data_org:10'b0)|
    ((_net_0)?_add_map_x_101_data_org_near:10'b0);
   assign  data_out_org249 = ((_net_1)?_add_map_x_102_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_102_data_org:10'b0);
   assign  data_out_org250 = ((_net_1)?_add_map_x_102_data_org:10'b0)|
    ((_net_0)?_add_map_x_102_data_org_near:10'b0);
   assign  data_out_org251 = ((_net_1)?_add_map_x_103_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_103_data_org:10'b0);
   assign  data_out_org252 = ((_net_1)?_add_map_x_103_data_org:10'b0)|
    ((_net_0)?_add_map_x_103_data_org_near:10'b0);
   assign  data_out_org253 = ((_net_1)?_add_map_x_104_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_104_data_org:10'b0);
   assign  data_out_org254 = ((_net_1)?_add_map_x_104_data_org:10'b0)|
    ((_net_0)?_add_map_x_104_data_org_near:10'b0);
   assign  data_out_org257 = ((_net_1)?_add_map_x_105_data_org:10'b0)|
    ((_net_0)?_add_map_x_105_data_org_near:10'b0);
   assign  data_out_org258 = ((_net_1)?_add_map_x_105_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_105_data_org:10'b0);
   assign  data_out_org259 = ((_net_1)?_add_map_x_106_data_org:10'b0)|
    ((_net_0)?_add_map_x_106_data_org_near:10'b0);
   assign  data_out_org260 = ((_net_1)?_add_map_x_106_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_106_data_org:10'b0);
   assign  data_out_org261 = ((_net_1)?_add_map_x_107_data_org:10'b0)|
    ((_net_0)?_add_map_x_107_data_org_near:10'b0);
   assign  data_out_org262 = ((_net_1)?_add_map_x_107_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_107_data_org:10'b0);
   assign  data_out_org263 = ((_net_1)?_add_map_x_108_data_org:10'b0)|
    ((_net_0)?_add_map_x_108_data_org_near:10'b0);
   assign  data_out_org264 = ((_net_1)?_add_map_x_108_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_108_data_org:10'b0);
   assign  data_out_org265 = ((_net_1)?_add_map_x_109_data_org:10'b0)|
    ((_net_0)?_add_map_x_109_data_org_near:10'b0);
   assign  data_out_org266 = ((_net_1)?_add_map_x_109_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_109_data_org:10'b0);
   assign  data_out_org267 = ((_net_1)?_add_map_x_110_data_org:10'b0)|
    ((_net_0)?_add_map_x_110_data_org_near:10'b0);
   assign  data_out_org268 = ((_net_1)?_add_map_x_110_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_110_data_org:10'b0);
   assign  data_out_org269 = ((_net_1)?_add_map_x_111_data_org:10'b0)|
    ((_net_0)?_add_map_x_111_data_org_near:10'b0);
   assign  data_out_org270 = ((_net_1)?_add_map_x_111_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_111_data_org:10'b0);
   assign  data_out_org271 = ((_net_1)?_add_map_x_112_data_org:10'b0)|
    ((_net_0)?_add_map_x_112_data_org_near:10'b0);
   assign  data_out_org272 = ((_net_1)?_add_map_x_112_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_112_data_org:10'b0);
   assign  data_out_org273 = ((_net_1)?_add_map_x_113_data_org:10'b0)|
    ((_net_0)?_add_map_x_113_data_org_near:10'b0);
   assign  data_out_org274 = ((_net_1)?_add_map_x_113_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_113_data_org:10'b0);
   assign  data_out_org275 = ((_net_1)?_add_map_x_114_data_org:10'b0)|
    ((_net_0)?_add_map_x_114_data_org_near:10'b0);
   assign  data_out_org276 = ((_net_1)?_add_map_x_114_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_114_data_org:10'b0);
   assign  data_out_org277 = ((_net_1)?_add_map_x_115_data_org:10'b0)|
    ((_net_0)?_add_map_x_115_data_org_near:10'b0);
   assign  data_out_org278 = ((_net_1)?_add_map_x_115_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_115_data_org:10'b0);
   assign  data_out_org279 = ((_net_1)?_add_map_x_116_data_org:10'b0)|
    ((_net_0)?_add_map_x_116_data_org_near:10'b0);
   assign  data_out_org280 = ((_net_1)?_add_map_x_116_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_116_data_org:10'b0);
   assign  data_out_org281 = ((_net_1)?_add_map_x_117_data_org:10'b0)|
    ((_net_0)?_add_map_x_117_data_org_near:10'b0);
   assign  data_out_org282 = ((_net_1)?_add_map_x_117_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_117_data_org:10'b0);
   assign  data_out_org283 = ((_net_1)?_add_map_x_118_data_org:10'b0)|
    ((_net_0)?_add_map_x_118_data_org_near:10'b0);
   assign  data_out_org284 = ((_net_1)?_add_map_x_118_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_118_data_org:10'b0);
   assign  data_out_org285 = ((_net_1)?_add_map_x_119_data_org:10'b0)|
    ((_net_0)?_add_map_x_119_data_org_near:10'b0);
   assign  data_out_org286 = ((_net_1)?_add_map_x_119_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_119_data_org:10'b0);
   assign  data_out_org289 = ((_net_1)?_add_map_x_120_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_120_data_org:10'b0);
   assign  data_out_org290 = ((_net_1)?_add_map_x_120_data_org:10'b0)|
    ((_net_0)?_add_map_x_120_data_org_near:10'b0);
   assign  data_out_org291 = ((_net_1)?_add_map_x_121_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_121_data_org:10'b0);
   assign  data_out_org292 = ((_net_1)?_add_map_x_121_data_org:10'b0)|
    ((_net_0)?_add_map_x_121_data_org_near:10'b0);
   assign  data_out_org293 = ((_net_1)?_add_map_x_122_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_122_data_org:10'b0);
   assign  data_out_org294 = ((_net_1)?_add_map_x_122_data_org:10'b0)|
    ((_net_0)?_add_map_x_122_data_org_near:10'b0);
   assign  data_out_org295 = ((_net_1)?_add_map_x_123_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_123_data_org:10'b0);
   assign  data_out_org296 = ((_net_1)?_add_map_x_123_data_org:10'b0)|
    ((_net_0)?_add_map_x_123_data_org_near:10'b0);
   assign  data_out_org297 = ((_net_1)?_add_map_x_124_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_124_data_org:10'b0);
   assign  data_out_org298 = ((_net_1)?_add_map_x_124_data_org:10'b0)|
    ((_net_0)?_add_map_x_124_data_org_near:10'b0);
   assign  data_out_org299 = ((_net_1)?_add_map_x_125_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_125_data_org:10'b0);
   assign  data_out_org300 = ((_net_1)?_add_map_x_125_data_org:10'b0)|
    ((_net_0)?_add_map_x_125_data_org_near:10'b0);
   assign  data_out_org301 = ((_net_1)?_add_map_x_126_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_126_data_org:10'b0);
   assign  data_out_org302 = ((_net_1)?_add_map_x_126_data_org:10'b0)|
    ((_net_0)?_add_map_x_126_data_org_near:10'b0);
   assign  data_out_org303 = ((_net_1)?_add_map_x_127_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_127_data_org:10'b0);
   assign  data_out_org304 = ((_net_1)?_add_map_x_127_data_org:10'b0)|
    ((_net_0)?_add_map_x_127_data_org_near:10'b0);
   assign  data_out_org305 = ((_net_1)?_add_map_x_128_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_128_data_org:10'b0);
   assign  data_out_org306 = ((_net_1)?_add_map_x_128_data_org:10'b0)|
    ((_net_0)?_add_map_x_128_data_org_near:10'b0);
   assign  data_out_org307 = ((_net_1)?_add_map_x_129_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_129_data_org:10'b0);
   assign  data_out_org308 = ((_net_1)?_add_map_x_129_data_org:10'b0)|
    ((_net_0)?_add_map_x_129_data_org_near:10'b0);
   assign  data_out_org309 = ((_net_1)?_add_map_x_130_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_130_data_org:10'b0);
   assign  data_out_org310 = ((_net_1)?_add_map_x_130_data_org:10'b0)|
    ((_net_0)?_add_map_x_130_data_org_near:10'b0);
   assign  data_out_org311 = ((_net_1)?_add_map_x_131_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_131_data_org:10'b0);
   assign  data_out_org312 = ((_net_1)?_add_map_x_131_data_org:10'b0)|
    ((_net_0)?_add_map_x_131_data_org_near:10'b0);
   assign  data_out_org313 = ((_net_1)?_add_map_x_132_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_132_data_org:10'b0);
   assign  data_out_org314 = ((_net_1)?_add_map_x_132_data_org:10'b0)|
    ((_net_0)?_add_map_x_132_data_org_near:10'b0);
   assign  data_out_org315 = ((_net_1)?_add_map_x_133_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_133_data_org:10'b0);
   assign  data_out_org316 = ((_net_1)?_add_map_x_133_data_org:10'b0)|
    ((_net_0)?_add_map_x_133_data_org_near:10'b0);
   assign  data_out_org317 = ((_net_1)?_add_map_x_134_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_134_data_org:10'b0);
   assign  data_out_org318 = ((_net_1)?_add_map_x_134_data_org:10'b0)|
    ((_net_0)?_add_map_x_134_data_org_near:10'b0);
   assign  data_out_org321 = ((_net_1)?_add_map_x_135_data_org:10'b0)|
    ((_net_0)?_add_map_x_135_data_org_near:10'b0);
   assign  data_out_org322 = ((_net_1)?_add_map_x_135_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_135_data_org:10'b0);
   assign  data_out_org323 = ((_net_1)?_add_map_x_136_data_org:10'b0)|
    ((_net_0)?_add_map_x_136_data_org_near:10'b0);
   assign  data_out_org324 = ((_net_1)?_add_map_x_136_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_136_data_org:10'b0);
   assign  data_out_org325 = ((_net_1)?_add_map_x_137_data_org:10'b0)|
    ((_net_0)?_add_map_x_137_data_org_near:10'b0);
   assign  data_out_org326 = ((_net_1)?_add_map_x_137_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_137_data_org:10'b0);
   assign  data_out_org327 = ((_net_1)?_add_map_x_138_data_org:10'b0)|
    ((_net_0)?_add_map_x_138_data_org_near:10'b0);
   assign  data_out_org328 = ((_net_1)?_add_map_x_138_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_138_data_org:10'b0);
   assign  data_out_org329 = ((_net_1)?_add_map_x_139_data_org:10'b0)|
    ((_net_0)?_add_map_x_139_data_org_near:10'b0);
   assign  data_out_org330 = ((_net_1)?_add_map_x_139_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_139_data_org:10'b0);
   assign  data_out_org331 = ((_net_1)?_add_map_x_140_data_org:10'b0)|
    ((_net_0)?_add_map_x_140_data_org_near:10'b0);
   assign  data_out_org332 = ((_net_1)?_add_map_x_140_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_140_data_org:10'b0);
   assign  data_out_org333 = ((_net_1)?_add_map_x_141_data_org:10'b0)|
    ((_net_0)?_add_map_x_141_data_org_near:10'b0);
   assign  data_out_org334 = ((_net_1)?_add_map_x_141_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_141_data_org:10'b0);
   assign  data_out_org335 = ((_net_1)?_add_map_x_142_data_org:10'b0)|
    ((_net_0)?_add_map_x_142_data_org_near:10'b0);
   assign  data_out_org336 = ((_net_1)?_add_map_x_142_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_142_data_org:10'b0);
   assign  data_out_org337 = ((_net_1)?_add_map_x_143_data_org:10'b0)|
    ((_net_0)?_add_map_x_143_data_org_near:10'b0);
   assign  data_out_org338 = ((_net_1)?_add_map_x_143_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_143_data_org:10'b0);
   assign  data_out_org339 = ((_net_1)?_add_map_x_144_data_org:10'b0)|
    ((_net_0)?_add_map_x_144_data_org_near:10'b0);
   assign  data_out_org340 = ((_net_1)?_add_map_x_144_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_144_data_org:10'b0);
   assign  data_out_org341 = ((_net_1)?_add_map_x_145_data_org:10'b0)|
    ((_net_0)?_add_map_x_145_data_org_near:10'b0);
   assign  data_out_org342 = ((_net_1)?_add_map_x_145_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_145_data_org:10'b0);
   assign  data_out_org343 = ((_net_1)?_add_map_x_146_data_org:10'b0)|
    ((_net_0)?_add_map_x_146_data_org_near:10'b0);
   assign  data_out_org344 = ((_net_1)?_add_map_x_146_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_146_data_org:10'b0);
   assign  data_out_org345 = ((_net_1)?_add_map_x_147_data_org:10'b0)|
    ((_net_0)?_add_map_x_147_data_org_near:10'b0);
   assign  data_out_org346 = ((_net_1)?_add_map_x_147_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_147_data_org:10'b0);
   assign  data_out_org347 = ((_net_1)?_add_map_x_148_data_org:10'b0)|
    ((_net_0)?_add_map_x_148_data_org_near:10'b0);
   assign  data_out_org348 = ((_net_1)?_add_map_x_148_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_148_data_org:10'b0);
   assign  data_out_org349 = ((_net_1)?_add_map_x_149_data_org:10'b0)|
    ((_net_0)?_add_map_x_149_data_org_near:10'b0);
   assign  data_out_org350 = ((_net_1)?_add_map_x_149_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_149_data_org:10'b0);
   assign  data_out_org353 = ((_net_1)?_add_map_x_150_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_150_data_org:10'b0);
   assign  data_out_org354 = ((_net_1)?_add_map_x_150_data_org:10'b0)|
    ((_net_0)?_add_map_x_150_data_org_near:10'b0);
   assign  data_out_org355 = ((_net_1)?_add_map_x_151_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_151_data_org:10'b0);
   assign  data_out_org356 = ((_net_1)?_add_map_x_151_data_org:10'b0)|
    ((_net_0)?_add_map_x_151_data_org_near:10'b0);
   assign  data_out_org357 = ((_net_1)?_add_map_x_152_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_152_data_org:10'b0);
   assign  data_out_org358 = ((_net_1)?_add_map_x_152_data_org:10'b0)|
    ((_net_0)?_add_map_x_152_data_org_near:10'b0);
   assign  data_out_org359 = ((_net_1)?_add_map_x_153_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_153_data_org:10'b0);
   assign  data_out_org360 = ((_net_1)?_add_map_x_153_data_org:10'b0)|
    ((_net_0)?_add_map_x_153_data_org_near:10'b0);
   assign  data_out_org361 = ((_net_1)?_add_map_x_154_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_154_data_org:10'b0);
   assign  data_out_org362 = ((_net_1)?_add_map_x_154_data_org:10'b0)|
    ((_net_0)?_add_map_x_154_data_org_near:10'b0);
   assign  data_out_org363 = ((_net_1)?_add_map_x_155_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_155_data_org:10'b0);
   assign  data_out_org364 = ((_net_1)?_add_map_x_155_data_org:10'b0)|
    ((_net_0)?_add_map_x_155_data_org_near:10'b0);
   assign  data_out_org365 = ((_net_1)?_add_map_x_156_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_156_data_org:10'b0);
   assign  data_out_org366 = ((_net_1)?_add_map_x_156_data_org:10'b0)|
    ((_net_0)?_add_map_x_156_data_org_near:10'b0);
   assign  data_out_org367 = ((_net_1)?_add_map_x_157_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_157_data_org:10'b0);
   assign  data_out_org368 = ((_net_1)?_add_map_x_157_data_org:10'b0)|
    ((_net_0)?_add_map_x_157_data_org_near:10'b0);
   assign  data_out_org369 = ((_net_1)?_add_map_x_158_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_158_data_org:10'b0);
   assign  data_out_org370 = ((_net_1)?_add_map_x_158_data_org:10'b0)|
    ((_net_0)?_add_map_x_158_data_org_near:10'b0);
   assign  data_out_org371 = ((_net_1)?_add_map_x_159_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_159_data_org:10'b0);
   assign  data_out_org372 = ((_net_1)?_add_map_x_159_data_org:10'b0)|
    ((_net_0)?_add_map_x_159_data_org_near:10'b0);
   assign  data_out_org373 = ((_net_1)?_add_map_x_160_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_160_data_org:10'b0);
   assign  data_out_org374 = ((_net_1)?_add_map_x_160_data_org:10'b0)|
    ((_net_0)?_add_map_x_160_data_org_near:10'b0);
   assign  data_out_org375 = ((_net_1)?_add_map_x_161_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_161_data_org:10'b0);
   assign  data_out_org376 = ((_net_1)?_add_map_x_161_data_org:10'b0)|
    ((_net_0)?_add_map_x_161_data_org_near:10'b0);
   assign  data_out_org377 = ((_net_1)?_add_map_x_162_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_162_data_org:10'b0);
   assign  data_out_org378 = ((_net_1)?_add_map_x_162_data_org:10'b0)|
    ((_net_0)?_add_map_x_162_data_org_near:10'b0);
   assign  data_out_org379 = ((_net_1)?_add_map_x_163_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_163_data_org:10'b0);
   assign  data_out_org380 = ((_net_1)?_add_map_x_163_data_org:10'b0)|
    ((_net_0)?_add_map_x_163_data_org_near:10'b0);
   assign  data_out_org381 = ((_net_1)?_add_map_x_164_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_164_data_org:10'b0);
   assign  data_out_org382 = ((_net_1)?_add_map_x_164_data_org:10'b0)|
    ((_net_0)?_add_map_x_164_data_org_near:10'b0);
   assign  data_out_org385 = ((_net_1)?_add_map_x_165_data_org:10'b0)|
    ((_net_0)?_add_map_x_165_data_org_near:10'b0);
   assign  data_out_org386 = ((_net_1)?_add_map_x_165_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_165_data_org:10'b0);
   assign  data_out_org387 = ((_net_1)?_add_map_x_166_data_org:10'b0)|
    ((_net_0)?_add_map_x_166_data_org_near:10'b0);
   assign  data_out_org388 = ((_net_1)?_add_map_x_166_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_166_data_org:10'b0);
   assign  data_out_org389 = ((_net_1)?_add_map_x_167_data_org:10'b0)|
    ((_net_0)?_add_map_x_167_data_org_near:10'b0);
   assign  data_out_org390 = ((_net_1)?_add_map_x_167_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_167_data_org:10'b0);
   assign  data_out_org391 = ((_net_1)?_add_map_x_168_data_org:10'b0)|
    ((_net_0)?_add_map_x_168_data_org_near:10'b0);
   assign  data_out_org392 = ((_net_1)?_add_map_x_168_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_168_data_org:10'b0);
   assign  data_out_org393 = ((_net_1)?_add_map_x_169_data_org:10'b0)|
    ((_net_0)?_add_map_x_169_data_org_near:10'b0);
   assign  data_out_org394 = ((_net_1)?_add_map_x_169_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_169_data_org:10'b0);
   assign  data_out_org395 = ((_net_1)?_add_map_x_170_data_org:10'b0)|
    ((_net_0)?_add_map_x_170_data_org_near:10'b0);
   assign  data_out_org396 = ((_net_1)?_add_map_x_170_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_170_data_org:10'b0);
   assign  data_out_org397 = ((_net_1)?_add_map_x_171_data_org:10'b0)|
    ((_net_0)?_add_map_x_171_data_org_near:10'b0);
   assign  data_out_org398 = ((_net_1)?_add_map_x_171_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_171_data_org:10'b0);
   assign  data_out_org399 = ((_net_1)?_add_map_x_172_data_org:10'b0)|
    ((_net_0)?_add_map_x_172_data_org_near:10'b0);
   assign  data_out_org400 = ((_net_1)?_add_map_x_172_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_172_data_org:10'b0);
   assign  data_out_org401 = ((_net_1)?_add_map_x_173_data_org:10'b0)|
    ((_net_0)?_add_map_x_173_data_org_near:10'b0);
   assign  data_out_org402 = ((_net_1)?_add_map_x_173_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_173_data_org:10'b0);
   assign  data_out_org403 = ((_net_1)?_add_map_x_174_data_org:10'b0)|
    ((_net_0)?_add_map_x_174_data_org_near:10'b0);
   assign  data_out_org404 = ((_net_1)?_add_map_x_174_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_174_data_org:10'b0);
   assign  data_out_org405 = ((_net_1)?_add_map_x_175_data_org:10'b0)|
    ((_net_0)?_add_map_x_175_data_org_near:10'b0);
   assign  data_out_org406 = ((_net_1)?_add_map_x_175_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_175_data_org:10'b0);
   assign  data_out_org407 = ((_net_1)?_add_map_x_176_data_org:10'b0)|
    ((_net_0)?_add_map_x_176_data_org_near:10'b0);
   assign  data_out_org408 = ((_net_1)?_add_map_x_176_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_176_data_org:10'b0);
   assign  data_out_org409 = ((_net_1)?_add_map_x_177_data_org:10'b0)|
    ((_net_0)?_add_map_x_177_data_org_near:10'b0);
   assign  data_out_org410 = ((_net_1)?_add_map_x_177_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_177_data_org:10'b0);
   assign  data_out_org411 = ((_net_1)?_add_map_x_178_data_org:10'b0)|
    ((_net_0)?_add_map_x_178_data_org_near:10'b0);
   assign  data_out_org412 = ((_net_1)?_add_map_x_178_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_178_data_org:10'b0);
   assign  data_out_org413 = ((_net_1)?_add_map_x_179_data_org:10'b0)|
    ((_net_0)?_add_map_x_179_data_org_near:10'b0);
   assign  data_out_org414 = ((_net_1)?_add_map_x_179_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_179_data_org:10'b0);
   assign  data_out_org417 = ((_net_1)?_add_map_x_180_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_180_data_org:10'b0);
   assign  data_out_org418 = ((_net_1)?_add_map_x_180_data_org:10'b0)|
    ((_net_0)?_add_map_x_180_data_org_near:10'b0);
   assign  data_out_org419 = ((_net_1)?_add_map_x_181_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_181_data_org:10'b0);
   assign  data_out_org420 = ((_net_1)?_add_map_x_181_data_org:10'b0)|
    ((_net_0)?_add_map_x_181_data_org_near:10'b0);
   assign  data_out_org421 = ((_net_1)?_add_map_x_182_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_182_data_org:10'b0);
   assign  data_out_org422 = ((_net_1)?_add_map_x_182_data_org:10'b0)|
    ((_net_0)?_add_map_x_182_data_org_near:10'b0);
   assign  data_out_org423 = ((_net_1)?_add_map_x_183_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_183_data_org:10'b0);
   assign  data_out_org424 = ((_net_1)?_add_map_x_183_data_org:10'b0)|
    ((_net_0)?_add_map_x_183_data_org_near:10'b0);
   assign  data_out_org425 = ((_net_1)?_add_map_x_184_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_184_data_org:10'b0);
   assign  data_out_org426 = ((_net_1)?_add_map_x_184_data_org:10'b0)|
    ((_net_0)?_add_map_x_184_data_org_near:10'b0);
   assign  data_out_org427 = ((_net_1)?_add_map_x_185_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_185_data_org:10'b0);
   assign  data_out_org428 = ((_net_1)?_add_map_x_185_data_org:10'b0)|
    ((_net_0)?_add_map_x_185_data_org_near:10'b0);
   assign  data_out_org429 = ((_net_1)?_add_map_x_186_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_186_data_org:10'b0);
   assign  data_out_org430 = ((_net_1)?_add_map_x_186_data_org:10'b0)|
    ((_net_0)?_add_map_x_186_data_org_near:10'b0);
   assign  data_out_org431 = ((_net_1)?_add_map_x_187_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_187_data_org:10'b0);
   assign  data_out_org432 = ((_net_1)?_add_map_x_187_data_org:10'b0)|
    ((_net_0)?_add_map_x_187_data_org_near:10'b0);
   assign  data_out_org433 = ((_net_1)?_add_map_x_188_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_188_data_org:10'b0);
   assign  data_out_org434 = ((_net_1)?_add_map_x_188_data_org:10'b0)|
    ((_net_0)?_add_map_x_188_data_org_near:10'b0);
   assign  data_out_org435 = ((_net_1)?_add_map_x_189_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_189_data_org:10'b0);
   assign  data_out_org436 = ((_net_1)?_add_map_x_189_data_org:10'b0)|
    ((_net_0)?_add_map_x_189_data_org_near:10'b0);
   assign  data_out_org437 = ((_net_1)?_add_map_x_190_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_190_data_org:10'b0);
   assign  data_out_org438 = ((_net_1)?_add_map_x_190_data_org:10'b0)|
    ((_net_0)?_add_map_x_190_data_org_near:10'b0);
   assign  data_out_org439 = ((_net_1)?_add_map_x_191_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_191_data_org:10'b0);
   assign  data_out_org440 = ((_net_1)?_add_map_x_191_data_org:10'b0)|
    ((_net_0)?_add_map_x_191_data_org_near:10'b0);
   assign  data_out_org441 = ((_net_1)?_add_map_x_192_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_192_data_org:10'b0);
   assign  data_out_org442 = ((_net_1)?_add_map_x_192_data_org:10'b0)|
    ((_net_0)?_add_map_x_192_data_org_near:10'b0);
   assign  data_out_org443 = ((_net_1)?_add_map_x_193_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_193_data_org:10'b0);
   assign  data_out_org444 = ((_net_1)?_add_map_x_193_data_org:10'b0)|
    ((_net_0)?_add_map_x_193_data_org_near:10'b0);
   assign  data_out_org445 = ((_net_1)?_add_map_x_194_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_194_data_org:10'b0);
   assign  data_out_org446 = ((_net_1)?_add_map_x_194_data_org:10'b0)|
    ((_net_0)?_add_map_x_194_data_org_near:10'b0);
   assign  data_out_org449 = ((_net_1)?_add_map_x_195_data_org:10'b0)|
    ((_net_0)?_add_map_x_195_data_org_near:10'b0);
   assign  data_out_org450 = ((_net_1)?_add_map_x_195_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_195_data_org:10'b0);
   assign  data_out_org451 = ((_net_1)?_add_map_x_196_data_org:10'b0)|
    ((_net_0)?_add_map_x_196_data_org_near:10'b0);
   assign  data_out_org452 = ((_net_1)?_add_map_x_196_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_196_data_org:10'b0);
   assign  data_out_org453 = ((_net_1)?_add_map_x_197_data_org:10'b0)|
    ((_net_0)?_add_map_x_197_data_org_near:10'b0);
   assign  data_out_org454 = ((_net_1)?_add_map_x_197_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_197_data_org:10'b0);
   assign  data_out_org455 = ((_net_1)?_add_map_x_198_data_org:10'b0)|
    ((_net_0)?_add_map_x_198_data_org_near:10'b0);
   assign  data_out_org456 = ((_net_1)?_add_map_x_198_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_198_data_org:10'b0);
   assign  data_out_org457 = ((_net_1)?_add_map_x_199_data_org:10'b0)|
    ((_net_0)?_add_map_x_199_data_org_near:10'b0);
   assign  data_out_org458 = ((_net_1)?_add_map_x_199_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_199_data_org:10'b0);
   assign  data_out_org459 = ((_net_1)?_add_map_x_200_data_org:10'b0)|
    ((_net_0)?_add_map_x_200_data_org_near:10'b0);
   assign  data_out_org460 = ((_net_1)?_add_map_x_200_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_200_data_org:10'b0);
   assign  data_out_org461 = ((_net_1)?_add_map_x_201_data_org:10'b0)|
    ((_net_0)?_add_map_x_201_data_org_near:10'b0);
   assign  data_out_org462 = ((_net_1)?_add_map_x_201_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_201_data_org:10'b0);
   assign  data_out_org463 = ((_net_1)?_add_map_x_202_data_org:10'b0)|
    ((_net_0)?_add_map_x_202_data_org_near:10'b0);
   assign  data_out_org464 = ((_net_1)?_add_map_x_202_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_202_data_org:10'b0);
   assign  data_out_org465 = ((_net_1)?_add_map_x_203_data_org:10'b0)|
    ((_net_0)?_add_map_x_203_data_org_near:10'b0);
   assign  data_out_org466 = ((_net_1)?_add_map_x_203_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_203_data_org:10'b0);
   assign  data_out_org467 = ((_net_1)?_add_map_x_204_data_org:10'b0)|
    ((_net_0)?_add_map_x_204_data_org_near:10'b0);
   assign  data_out_org468 = ((_net_1)?_add_map_x_204_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_204_data_org:10'b0);
   assign  data_out_org469 = ((_net_1)?_add_map_x_205_data_org:10'b0)|
    ((_net_0)?_add_map_x_205_data_org_near:10'b0);
   assign  data_out_org470 = ((_net_1)?_add_map_x_205_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_205_data_org:10'b0);
   assign  data_out_org471 = ((_net_1)?_add_map_x_206_data_org:10'b0)|
    ((_net_0)?_add_map_x_206_data_org_near:10'b0);
   assign  data_out_org472 = ((_net_1)?_add_map_x_206_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_206_data_org:10'b0);
   assign  data_out_org473 = ((_net_1)?_add_map_x_207_data_org:10'b0)|
    ((_net_0)?_add_map_x_207_data_org_near:10'b0);
   assign  data_out_org474 = ((_net_1)?_add_map_x_207_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_207_data_org:10'b0);
   assign  data_out_org475 = ((_net_1)?_add_map_x_208_data_org:10'b0)|
    ((_net_0)?_add_map_x_208_data_org_near:10'b0);
   assign  data_out_org476 = ((_net_1)?_add_map_x_208_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_208_data_org:10'b0);
   assign  data_out_org477 = ((_net_1)?_add_map_x_209_data_org:10'b0)|
    ((_net_0)?_add_map_x_209_data_org_near:10'b0);
   assign  data_out_org478 = ((_net_1)?_add_map_x_209_data_org_near:10'b0)|
    ((_net_0)?_add_map_x_209_data_org:10'b0);
   assign  data_out33 = ((_net_1)?_add_map_x_data_near:10'b0)|
    ((_net_0)?_add_map_x_data_out:10'b0);
   assign  data_out34 = ((_net_1)?_add_map_x_data_out:10'b0)|
    ((_net_0)?_add_map_x_data_near:10'b0);
   assign  data_out35 = ((_net_1)?_add_map_x_1_data_near:10'b0)|
    ((_net_0)?_add_map_x_1_data_out:10'b0);
   assign  data_out36 = ((_net_1)?_add_map_x_1_data_out:10'b0)|
    ((_net_0)?_add_map_x_1_data_near:10'b0);
   assign  data_out37 = ((_net_1)?_add_map_x_2_data_near:10'b0)|
    ((_net_0)?_add_map_x_2_data_out:10'b0);
   assign  data_out38 = ((_net_1)?_add_map_x_2_data_out:10'b0)|
    ((_net_0)?_add_map_x_2_data_near:10'b0);
   assign  data_out39 = ((_net_1)?_add_map_x_3_data_near:10'b0)|
    ((_net_0)?_add_map_x_3_data_out:10'b0);
   assign  data_out40 = ((_net_1)?_add_map_x_3_data_out:10'b0)|
    ((_net_0)?_add_map_x_3_data_near:10'b0);
   assign  data_out41 = ((_net_1)?_add_map_x_4_data_near:10'b0)|
    ((_net_0)?_add_map_x_4_data_out:10'b0);
   assign  data_out42 = ((_net_1)?_add_map_x_4_data_out:10'b0)|
    ((_net_0)?_add_map_x_4_data_near:10'b0);
   assign  data_out43 = ((_net_1)?_add_map_x_5_data_near:10'b0)|
    ((_net_0)?_add_map_x_5_data_out:10'b0);
   assign  data_out44 = ((_net_1)?_add_map_x_5_data_out:10'b0)|
    ((_net_0)?_add_map_x_5_data_near:10'b0);
   assign  data_out45 = ((_net_1)?_add_map_x_6_data_near:10'b0)|
    ((_net_0)?_add_map_x_6_data_out:10'b0);
   assign  data_out46 = ((_net_1)?_add_map_x_6_data_out:10'b0)|
    ((_net_0)?_add_map_x_6_data_near:10'b0);
   assign  data_out47 = ((_net_1)?_add_map_x_7_data_near:10'b0)|
    ((_net_0)?_add_map_x_7_data_out:10'b0);
   assign  data_out48 = ((_net_1)?_add_map_x_7_data_out:10'b0)|
    ((_net_0)?_add_map_x_7_data_near:10'b0);
   assign  data_out49 = ((_net_1)?_add_map_x_8_data_near:10'b0)|
    ((_net_0)?_add_map_x_8_data_out:10'b0);
   assign  data_out50 = ((_net_1)?_add_map_x_8_data_out:10'b0)|
    ((_net_0)?_add_map_x_8_data_near:10'b0);
   assign  data_out51 = ((_net_1)?_add_map_x_9_data_near:10'b0)|
    ((_net_0)?_add_map_x_9_data_out:10'b0);
   assign  data_out52 = ((_net_1)?_add_map_x_9_data_out:10'b0)|
    ((_net_0)?_add_map_x_9_data_near:10'b0);
   assign  data_out53 = ((_net_1)?_add_map_x_10_data_near:10'b0)|
    ((_net_0)?_add_map_x_10_data_out:10'b0);
   assign  data_out54 = ((_net_1)?_add_map_x_10_data_out:10'b0)|
    ((_net_0)?_add_map_x_10_data_near:10'b0);
   assign  data_out55 = ((_net_1)?_add_map_x_11_data_near:10'b0)|
    ((_net_0)?_add_map_x_11_data_out:10'b0);
   assign  data_out56 = ((_net_1)?_add_map_x_11_data_out:10'b0)|
    ((_net_0)?_add_map_x_11_data_near:10'b0);
   assign  data_out57 = ((_net_1)?_add_map_x_12_data_near:10'b0)|
    ((_net_0)?_add_map_x_12_data_out:10'b0);
   assign  data_out58 = ((_net_1)?_add_map_x_12_data_out:10'b0)|
    ((_net_0)?_add_map_x_12_data_near:10'b0);
   assign  data_out59 = ((_net_1)?_add_map_x_13_data_near:10'b0)|
    ((_net_0)?_add_map_x_13_data_out:10'b0);
   assign  data_out60 = ((_net_1)?_add_map_x_13_data_out:10'b0)|
    ((_net_0)?_add_map_x_13_data_near:10'b0);
   assign  data_out61 = ((_net_1)?_add_map_x_14_data_near:10'b0)|
    ((_net_0)?_add_map_x_14_data_out:10'b0);
   assign  data_out62 = ((_net_1)?_add_map_x_14_data_out:10'b0)|
    ((_net_0)?_add_map_x_14_data_near:10'b0);
   assign  data_out65 = ((_net_1)?_add_map_x_15_data_out:10'b0)|
    ((_net_0)?_add_map_x_15_data_near:10'b0);
   assign  data_out66 = ((_net_1)?_add_map_x_15_data_near:10'b0)|
    ((_net_0)?_add_map_x_15_data_out:10'b0);
   assign  data_out67 = ((_net_1)?_add_map_x_16_data_out:10'b0)|
    ((_net_0)?_add_map_x_16_data_near:10'b0);
   assign  data_out68 = ((_net_1)?_add_map_x_16_data_near:10'b0)|
    ((_net_0)?_add_map_x_16_data_out:10'b0);
   assign  data_out69 = ((_net_1)?_add_map_x_17_data_out:10'b0)|
    ((_net_0)?_add_map_x_17_data_near:10'b0);
   assign  data_out70 = ((_net_1)?_add_map_x_17_data_near:10'b0)|
    ((_net_0)?_add_map_x_17_data_out:10'b0);
   assign  data_out71 = ((_net_1)?_add_map_x_18_data_out:10'b0)|
    ((_net_0)?_add_map_x_18_data_near:10'b0);
   assign  data_out72 = ((_net_1)?_add_map_x_18_data_near:10'b0)|
    ((_net_0)?_add_map_x_18_data_out:10'b0);
   assign  data_out73 = ((_net_1)?_add_map_x_19_data_out:10'b0)|
    ((_net_0)?_add_map_x_19_data_near:10'b0);
   assign  data_out74 = ((_net_1)?_add_map_x_19_data_near:10'b0)|
    ((_net_0)?_add_map_x_19_data_out:10'b0);
   assign  data_out75 = ((_net_1)?_add_map_x_20_data_out:10'b0)|
    ((_net_0)?_add_map_x_20_data_near:10'b0);
   assign  data_out76 = ((_net_1)?_add_map_x_20_data_near:10'b0)|
    ((_net_0)?_add_map_x_20_data_out:10'b0);
   assign  data_out77 = ((_net_1)?_add_map_x_21_data_out:10'b0)|
    ((_net_0)?_add_map_x_21_data_near:10'b0);
   assign  data_out78 = ((_net_1)?_add_map_x_21_data_near:10'b0)|
    ((_net_0)?_add_map_x_21_data_out:10'b0);
   assign  data_out79 = ((_net_1)?_add_map_x_22_data_out:10'b0)|
    ((_net_0)?_add_map_x_22_data_near:10'b0);
   assign  data_out80 = ((_net_1)?_add_map_x_22_data_near:10'b0)|
    ((_net_0)?_add_map_x_22_data_out:10'b0);
   assign  data_out81 = ((_net_1)?_add_map_x_23_data_out:10'b0)|
    ((_net_0)?_add_map_x_23_data_near:10'b0);
   assign  data_out82 = ((_net_1)?_add_map_x_23_data_near:10'b0)|
    ((_net_0)?_add_map_x_23_data_out:10'b0);
   assign  data_out83 = ((_net_1)?_add_map_x_24_data_out:10'b0)|
    ((_net_0)?_add_map_x_24_data_near:10'b0);
   assign  data_out84 = ((_net_1)?_add_map_x_24_data_near:10'b0)|
    ((_net_0)?_add_map_x_24_data_out:10'b0);
   assign  data_out85 = ((_net_1)?_add_map_x_25_data_out:10'b0)|
    ((_net_0)?_add_map_x_25_data_near:10'b0);
   assign  data_out86 = ((_net_1)?_add_map_x_25_data_near:10'b0)|
    ((_net_0)?_add_map_x_25_data_out:10'b0);
   assign  data_out87 = ((_net_1)?_add_map_x_26_data_out:10'b0)|
    ((_net_0)?_add_map_x_26_data_near:10'b0);
   assign  data_out88 = ((_net_1)?_add_map_x_26_data_near:10'b0)|
    ((_net_0)?_add_map_x_26_data_out:10'b0);
   assign  data_out89 = ((_net_1)?_add_map_x_27_data_out:10'b0)|
    ((_net_0)?_add_map_x_27_data_near:10'b0);
   assign  data_out90 = ((_net_1)?_add_map_x_27_data_near:10'b0)|
    ((_net_0)?_add_map_x_27_data_out:10'b0);
   assign  data_out91 = ((_net_1)?_add_map_x_28_data_out:10'b0)|
    ((_net_0)?_add_map_x_28_data_near:10'b0);
   assign  data_out92 = ((_net_1)?_add_map_x_28_data_near:10'b0)|
    ((_net_0)?_add_map_x_28_data_out:10'b0);
   assign  data_out93 = ((_net_1)?_add_map_x_29_data_out:10'b0)|
    ((_net_0)?_add_map_x_29_data_near:10'b0);
   assign  data_out94 = ((_net_1)?_add_map_x_29_data_near:10'b0)|
    ((_net_0)?_add_map_x_29_data_out:10'b0);
   assign  data_out97 = ((_net_1)?_add_map_x_30_data_near:10'b0)|
    ((_net_0)?_add_map_x_30_data_out:10'b0);
   assign  data_out98 = ((_net_1)?_add_map_x_30_data_out:10'b0)|
    ((_net_0)?_add_map_x_30_data_near:10'b0);
   assign  data_out99 = ((_net_1)?_add_map_x_31_data_near:10'b0)|
    ((_net_0)?_add_map_x_31_data_out:10'b0);
   assign  data_out100 = ((_net_1)?_add_map_x_31_data_out:10'b0)|
    ((_net_0)?_add_map_x_31_data_near:10'b0);
   assign  data_out101 = ((_net_1)?_add_map_x_32_data_near:10'b0)|
    ((_net_0)?_add_map_x_32_data_out:10'b0);
   assign  data_out102 = ((_net_1)?_add_map_x_32_data_out:10'b0)|
    ((_net_0)?_add_map_x_32_data_near:10'b0);
   assign  data_out103 = ((_net_1)?_add_map_x_33_data_near:10'b0)|
    ((_net_0)?_add_map_x_33_data_out:10'b0);
   assign  data_out104 = ((_net_1)?_add_map_x_33_data_out:10'b0)|
    ((_net_0)?_add_map_x_33_data_near:10'b0);
   assign  data_out105 = ((_net_1)?_add_map_x_34_data_near:10'b0)|
    ((_net_0)?_add_map_x_34_data_out:10'b0);
   assign  data_out106 = ((_net_1)?_add_map_x_34_data_out:10'b0)|
    ((_net_0)?_add_map_x_34_data_near:10'b0);
   assign  data_out107 = ((_net_1)?_add_map_x_35_data_near:10'b0)|
    ((_net_0)?_add_map_x_35_data_out:10'b0);
   assign  data_out108 = ((_net_1)?_add_map_x_35_data_out:10'b0)|
    ((_net_0)?_add_map_x_35_data_near:10'b0);
   assign  data_out109 = ((_net_1)?_add_map_x_36_data_near:10'b0)|
    ((_net_0)?_add_map_x_36_data_out:10'b0);
   assign  data_out110 = ((_net_1)?_add_map_x_36_data_out:10'b0)|
    ((_net_0)?_add_map_x_36_data_near:10'b0);
   assign  data_out111 = ((_net_1)?_add_map_x_37_data_near:10'b0)|
    ((_net_0)?_add_map_x_37_data_out:10'b0);
   assign  data_out112 = ((_net_1)?_add_map_x_37_data_out:10'b0)|
    ((_net_0)?_add_map_x_37_data_near:10'b0);
   assign  data_out113 = ((_net_1)?_add_map_x_38_data_near:10'b0)|
    ((_net_0)?_add_map_x_38_data_out:10'b0);
   assign  data_out114 = ((_net_1)?_add_map_x_38_data_out:10'b0)|
    ((_net_0)?_add_map_x_38_data_near:10'b0);
   assign  data_out115 = ((_net_1)?_add_map_x_39_data_near:10'b0)|
    ((_net_0)?_add_map_x_39_data_out:10'b0);
   assign  data_out116 = ((_net_1)?_add_map_x_39_data_out:10'b0)|
    ((_net_0)?_add_map_x_39_data_near:10'b0);
   assign  data_out117 = ((_net_1)?_add_map_x_40_data_near:10'b0)|
    ((_net_0)?_add_map_x_40_data_out:10'b0);
   assign  data_out118 = ((_net_1)?_add_map_x_40_data_out:10'b0)|
    ((_net_0)?_add_map_x_40_data_near:10'b0);
   assign  data_out119 = ((_net_1)?_add_map_x_41_data_near:10'b0)|
    ((_net_0)?_add_map_x_41_data_out:10'b0);
   assign  data_out120 = ((_net_1)?_add_map_x_41_data_out:10'b0)|
    ((_net_0)?_add_map_x_41_data_near:10'b0);
   assign  data_out121 = ((_net_1)?_add_map_x_42_data_near:10'b0)|
    ((_net_0)?_add_map_x_42_data_out:10'b0);
   assign  data_out122 = ((_net_1)?_add_map_x_42_data_out:10'b0)|
    ((_net_0)?_add_map_x_42_data_near:10'b0);
   assign  data_out123 = ((_net_1)?_add_map_x_43_data_near:10'b0)|
    ((_net_0)?_add_map_x_43_data_out:10'b0);
   assign  data_out124 = ((_net_1)?_add_map_x_43_data_out:10'b0)|
    ((_net_0)?_add_map_x_43_data_near:10'b0);
   assign  data_out125 = ((_net_1)?_add_map_x_44_data_near:10'b0)|
    ((_net_0)?_add_map_x_44_data_out:10'b0);
   assign  data_out126 = ((_net_1)?_add_map_x_44_data_out:10'b0)|
    ((_net_0)?_add_map_x_44_data_near:10'b0);
   assign  data_out129 = ((_net_1)?_add_map_x_45_data_out:10'b0)|
    ((_net_0)?_add_map_x_45_data_near:10'b0);
   assign  data_out130 = ((_net_1)?_add_map_x_45_data_near:10'b0)|
    ((_net_0)?_add_map_x_45_data_out:10'b0);
   assign  data_out131 = ((_net_1)?_add_map_x_46_data_out:10'b0)|
    ((_net_0)?_add_map_x_46_data_near:10'b0);
   assign  data_out132 = ((_net_1)?_add_map_x_46_data_near:10'b0)|
    ((_net_0)?_add_map_x_46_data_out:10'b0);
   assign  data_out133 = ((_net_1)?_add_map_x_47_data_out:10'b0)|
    ((_net_0)?_add_map_x_47_data_near:10'b0);
   assign  data_out134 = ((_net_1)?_add_map_x_47_data_near:10'b0)|
    ((_net_0)?_add_map_x_47_data_out:10'b0);
   assign  data_out135 = ((_net_1)?_add_map_x_48_data_out:10'b0)|
    ((_net_0)?_add_map_x_48_data_near:10'b0);
   assign  data_out136 = ((_net_1)?_add_map_x_48_data_near:10'b0)|
    ((_net_0)?_add_map_x_48_data_out:10'b0);
   assign  data_out137 = ((_net_1)?_add_map_x_49_data_out:10'b0)|
    ((_net_0)?_add_map_x_49_data_near:10'b0);
   assign  data_out138 = ((_net_1)?_add_map_x_49_data_near:10'b0)|
    ((_net_0)?_add_map_x_49_data_out:10'b0);
   assign  data_out139 = ((_net_1)?_add_map_x_50_data_out:10'b0)|
    ((_net_0)?_add_map_x_50_data_near:10'b0);
   assign  data_out140 = ((_net_1)?_add_map_x_50_data_near:10'b0)|
    ((_net_0)?_add_map_x_50_data_out:10'b0);
   assign  data_out141 = ((_net_1)?_add_map_x_51_data_out:10'b0)|
    ((_net_0)?_add_map_x_51_data_near:10'b0);
   assign  data_out142 = ((_net_1)?_add_map_x_51_data_near:10'b0)|
    ((_net_0)?_add_map_x_51_data_out:10'b0);
   assign  data_out143 = ((_net_1)?_add_map_x_52_data_out:10'b0)|
    ((_net_0)?_add_map_x_52_data_near:10'b0);
   assign  data_out144 = ((_net_1)?_add_map_x_52_data_near:10'b0)|
    ((_net_0)?_add_map_x_52_data_out:10'b0);
   assign  data_out145 = ((_net_1)?_add_map_x_53_data_out:10'b0)|
    ((_net_0)?_add_map_x_53_data_near:10'b0);
   assign  data_out146 = ((_net_1)?_add_map_x_53_data_near:10'b0)|
    ((_net_0)?_add_map_x_53_data_out:10'b0);
   assign  data_out147 = ((_net_1)?_add_map_x_54_data_out:10'b0)|
    ((_net_0)?_add_map_x_54_data_near:10'b0);
   assign  data_out148 = ((_net_1)?_add_map_x_54_data_near:10'b0)|
    ((_net_0)?_add_map_x_54_data_out:10'b0);
   assign  data_out149 = ((_net_1)?_add_map_x_55_data_out:10'b0)|
    ((_net_0)?_add_map_x_55_data_near:10'b0);
   assign  data_out150 = ((_net_1)?_add_map_x_55_data_near:10'b0)|
    ((_net_0)?_add_map_x_55_data_out:10'b0);
   assign  data_out151 = ((_net_1)?_add_map_x_56_data_out:10'b0)|
    ((_net_0)?_add_map_x_56_data_near:10'b0);
   assign  data_out152 = ((_net_1)?_add_map_x_56_data_near:10'b0)|
    ((_net_0)?_add_map_x_56_data_out:10'b0);
   assign  data_out153 = ((_net_1)?_add_map_x_57_data_out:10'b0)|
    ((_net_0)?_add_map_x_57_data_near:10'b0);
   assign  data_out154 = ((_net_1)?_add_map_x_57_data_near:10'b0)|
    ((_net_0)?_add_map_x_57_data_out:10'b0);
   assign  data_out155 = ((_net_1)?_add_map_x_58_data_out:10'b0)|
    ((_net_0)?_add_map_x_58_data_near:10'b0);
   assign  data_out156 = ((_net_1)?_add_map_x_58_data_near:10'b0)|
    ((_net_0)?_add_map_x_58_data_out:10'b0);
   assign  data_out157 = ((_net_1)?_add_map_x_59_data_out:10'b0)|
    ((_net_0)?_add_map_x_59_data_near:10'b0);
   assign  data_out158 = ((_net_1)?_add_map_x_59_data_near:10'b0)|
    ((_net_0)?_add_map_x_59_data_out:10'b0);
   assign  data_out161 = ((_net_1)?_add_map_x_60_data_near:10'b0)|
    ((_net_0)?_add_map_x_60_data_out:10'b0);
   assign  data_out162 = ((_net_1)?_add_map_x_60_data_out:10'b0)|
    ((_net_0)?_add_map_x_60_data_near:10'b0);
   assign  data_out163 = ((_net_1)?_add_map_x_61_data_near:10'b0)|
    ((_net_0)?_add_map_x_61_data_out:10'b0);
   assign  data_out164 = ((_net_1)?_add_map_x_61_data_out:10'b0)|
    ((_net_0)?_add_map_x_61_data_near:10'b0);
   assign  data_out165 = ((_net_1)?_add_map_x_62_data_near:10'b0)|
    ((_net_0)?_add_map_x_62_data_out:10'b0);
   assign  data_out166 = ((_net_1)?_add_map_x_62_data_out:10'b0)|
    ((_net_0)?_add_map_x_62_data_near:10'b0);
   assign  data_out167 = ((_net_1)?_add_map_x_63_data_near:10'b0)|
    ((_net_0)?_add_map_x_63_data_out:10'b0);
   assign  data_out168 = ((_net_1)?_add_map_x_63_data_out:10'b0)|
    ((_net_0)?_add_map_x_63_data_near:10'b0);
   assign  data_out169 = ((_net_1)?_add_map_x_64_data_near:10'b0)|
    ((_net_0)?_add_map_x_64_data_out:10'b0);
   assign  data_out170 = ((_net_1)?_add_map_x_64_data_out:10'b0)|
    ((_net_0)?_add_map_x_64_data_near:10'b0);
   assign  data_out171 = ((_net_1)?_add_map_x_65_data_near:10'b0)|
    ((_net_0)?_add_map_x_65_data_out:10'b0);
   assign  data_out172 = ((_net_1)?_add_map_x_65_data_out:10'b0)|
    ((_net_0)?_add_map_x_65_data_near:10'b0);
   assign  data_out173 = ((_net_1)?_add_map_x_66_data_near:10'b0)|
    ((_net_0)?_add_map_x_66_data_out:10'b0);
   assign  data_out174 = ((_net_1)?_add_map_x_66_data_out:10'b0)|
    ((_net_0)?_add_map_x_66_data_near:10'b0);
   assign  data_out175 = ((_net_1)?_add_map_x_67_data_near:10'b0)|
    ((_net_0)?_add_map_x_67_data_out:10'b0);
   assign  data_out176 = ((_net_1)?_add_map_x_67_data_out:10'b0)|
    ((_net_0)?_add_map_x_67_data_near:10'b0);
   assign  data_out177 = ((_net_1)?_add_map_x_68_data_near:10'b0)|
    ((_net_0)?_add_map_x_68_data_out:10'b0);
   assign  data_out178 = ((_net_1)?_add_map_x_68_data_out:10'b0)|
    ((_net_0)?_add_map_x_68_data_near:10'b0);
   assign  data_out179 = ((_net_1)?_add_map_x_69_data_near:10'b0)|
    ((_net_0)?_add_map_x_69_data_out:10'b0);
   assign  data_out180 = ((_net_1)?_add_map_x_69_data_out:10'b0)|
    ((_net_0)?_add_map_x_69_data_near:10'b0);
   assign  data_out181 = ((_net_1)?_add_map_x_70_data_near:10'b0)|
    ((_net_0)?_add_map_x_70_data_out:10'b0);
   assign  data_out182 = ((_net_1)?_add_map_x_70_data_out:10'b0)|
    ((_net_0)?_add_map_x_70_data_near:10'b0);
   assign  data_out183 = ((_net_1)?_add_map_x_71_data_near:10'b0)|
    ((_net_0)?_add_map_x_71_data_out:10'b0);
   assign  data_out184 = ((_net_1)?_add_map_x_71_data_out:10'b0)|
    ((_net_0)?_add_map_x_71_data_near:10'b0);
   assign  data_out185 = ((_net_1)?_add_map_x_72_data_near:10'b0)|
    ((_net_0)?_add_map_x_72_data_out:10'b0);
   assign  data_out186 = ((_net_1)?_add_map_x_72_data_out:10'b0)|
    ((_net_0)?_add_map_x_72_data_near:10'b0);
   assign  data_out187 = ((_net_1)?_add_map_x_73_data_near:10'b0)|
    ((_net_0)?_add_map_x_73_data_out:10'b0);
   assign  data_out188 = ((_net_1)?_add_map_x_73_data_out:10'b0)|
    ((_net_0)?_add_map_x_73_data_near:10'b0);
   assign  data_out189 = ((_net_1)?_add_map_x_74_data_near:10'b0)|
    ((_net_0)?_add_map_x_74_data_out:10'b0);
   assign  data_out190 = ((_net_1)?_add_map_x_74_data_out:10'b0)|
    ((_net_0)?_add_map_x_74_data_near:10'b0);
   assign  data_out193 = ((_net_1)?_add_map_x_75_data_out:10'b0)|
    ((_net_0)?_add_map_x_75_data_near:10'b0);
   assign  data_out194 = ((_net_1)?_add_map_x_75_data_near:10'b0)|
    ((_net_0)?_add_map_x_75_data_out:10'b0);
   assign  data_out195 = ((_net_1)?_add_map_x_76_data_out:10'b0)|
    ((_net_0)?_add_map_x_76_data_near:10'b0);
   assign  data_out196 = ((_net_1)?_add_map_x_76_data_near:10'b0)|
    ((_net_0)?_add_map_x_76_data_out:10'b0);
   assign  data_out197 = ((_net_1)?_add_map_x_77_data_out:10'b0)|
    ((_net_0)?_add_map_x_77_data_near:10'b0);
   assign  data_out198 = ((_net_1)?_add_map_x_77_data_near:10'b0)|
    ((_net_0)?_add_map_x_77_data_out:10'b0);
   assign  data_out199 = ((_net_1)?_add_map_x_78_data_out:10'b0)|
    ((_net_0)?_add_map_x_78_data_near:10'b0);
   assign  data_out200 = ((_net_1)?_add_map_x_78_data_near:10'b0)|
    ((_net_0)?_add_map_x_78_data_out:10'b0);
   assign  data_out201 = ((_net_1)?_add_map_x_79_data_out:10'b0)|
    ((_net_0)?_add_map_x_79_data_near:10'b0);
   assign  data_out202 = ((_net_1)?_add_map_x_79_data_near:10'b0)|
    ((_net_0)?_add_map_x_79_data_out:10'b0);
   assign  data_out203 = ((_net_1)?_add_map_x_80_data_out:10'b0)|
    ((_net_0)?_add_map_x_80_data_near:10'b0);
   assign  data_out204 = ((_net_1)?_add_map_x_80_data_near:10'b0)|
    ((_net_0)?_add_map_x_80_data_out:10'b0);
   assign  data_out205 = ((_net_1)?_add_map_x_81_data_out:10'b0)|
    ((_net_0)?_add_map_x_81_data_near:10'b0);
   assign  data_out206 = ((_net_1)?_add_map_x_81_data_near:10'b0)|
    ((_net_0)?_add_map_x_81_data_out:10'b0);
   assign  data_out207 = ((_net_1)?_add_map_x_82_data_out:10'b0)|
    ((_net_0)?_add_map_x_82_data_near:10'b0);
   assign  data_out208 = ((_net_1)?_add_map_x_82_data_near:10'b0)|
    ((_net_0)?_add_map_x_82_data_out:10'b0);
   assign  data_out209 = ((_net_1)?_add_map_x_83_data_out:10'b0)|
    ((_net_0)?_add_map_x_83_data_near:10'b0);
   assign  data_out210 = ((_net_1)?_add_map_x_83_data_near:10'b0)|
    ((_net_0)?_add_map_x_83_data_out:10'b0);
   assign  data_out211 = ((_net_1)?_add_map_x_84_data_out:10'b0)|
    ((_net_0)?_add_map_x_84_data_near:10'b0);
   assign  data_out212 = ((_net_1)?_add_map_x_84_data_near:10'b0)|
    ((_net_0)?_add_map_x_84_data_out:10'b0);
   assign  data_out213 = ((_net_1)?_add_map_x_85_data_out:10'b0)|
    ((_net_0)?_add_map_x_85_data_near:10'b0);
   assign  data_out214 = ((_net_1)?_add_map_x_85_data_near:10'b0)|
    ((_net_0)?_add_map_x_85_data_out:10'b0);
   assign  data_out215 = ((_net_1)?_add_map_x_86_data_out:10'b0)|
    ((_net_0)?_add_map_x_86_data_near:10'b0);
   assign  data_out216 = ((_net_1)?_add_map_x_86_data_near:10'b0)|
    ((_net_0)?_add_map_x_86_data_out:10'b0);
   assign  data_out217 = ((_net_1)?_add_map_x_87_data_out:10'b0)|
    ((_net_0)?_add_map_x_87_data_near:10'b0);
   assign  data_out218 = ((_net_1)?_add_map_x_87_data_near:10'b0)|
    ((_net_0)?_add_map_x_87_data_out:10'b0);
   assign  data_out219 = ((_net_1)?_add_map_x_88_data_out:10'b0)|
    ((_net_0)?_add_map_x_88_data_near:10'b0);
   assign  data_out220 = ((_net_1)?_add_map_x_88_data_near:10'b0)|
    ((_net_0)?_add_map_x_88_data_out:10'b0);
   assign  data_out221 = ((_net_1)?_add_map_x_89_data_out:10'b0)|
    ((_net_0)?_add_map_x_89_data_near:10'b0);
   assign  data_out222 = ((_net_1)?_add_map_x_89_data_near:10'b0)|
    ((_net_0)?_add_map_x_89_data_out:10'b0);
   assign  data_out225 = ((_net_1)?_add_map_x_90_data_near:10'b0)|
    ((_net_0)?_add_map_x_90_data_out:10'b0);
   assign  data_out226 = ((_net_1)?_add_map_x_90_data_out:10'b0)|
    ((_net_0)?_add_map_x_90_data_near:10'b0);
   assign  data_out227 = ((_net_1)?_add_map_x_91_data_near:10'b0)|
    ((_net_0)?_add_map_x_91_data_out:10'b0);
   assign  data_out228 = ((_net_1)?_add_map_x_91_data_out:10'b0)|
    ((_net_0)?_add_map_x_91_data_near:10'b0);
   assign  data_out229 = ((_net_1)?_add_map_x_92_data_near:10'b0)|
    ((_net_0)?_add_map_x_92_data_out:10'b0);
   assign  data_out230 = ((_net_1)?_add_map_x_92_data_out:10'b0)|
    ((_net_0)?_add_map_x_92_data_near:10'b0);
   assign  data_out231 = ((_net_1)?_add_map_x_93_data_near:10'b0)|
    ((_net_0)?_add_map_x_93_data_out:10'b0);
   assign  data_out232 = ((_net_1)?_add_map_x_93_data_out:10'b0)|
    ((_net_0)?_add_map_x_93_data_near:10'b0);
   assign  data_out233 = ((_net_1)?_add_map_x_94_data_near:10'b0)|
    ((_net_0)?_add_map_x_94_data_out:10'b0);
   assign  data_out234 = ((_net_1)?_add_map_x_94_data_out:10'b0)|
    ((_net_0)?_add_map_x_94_data_near:10'b0);
   assign  data_out235 = ((_net_1)?_add_map_x_95_data_near:10'b0)|
    ((_net_0)?_add_map_x_95_data_out:10'b0);
   assign  data_out236 = ((_net_1)?_add_map_x_95_data_out:10'b0)|
    ((_net_0)?_add_map_x_95_data_near:10'b0);
   assign  data_out237 = ((_net_1)?_add_map_x_96_data_near:10'b0)|
    ((_net_0)?_add_map_x_96_data_out:10'b0);
   assign  data_out238 = ((_net_1)?_add_map_x_96_data_out:10'b0)|
    ((_net_0)?_add_map_x_96_data_near:10'b0);
   assign  data_out239 = ((_net_1)?_add_map_x_97_data_near:10'b0)|
    ((_net_0)?_add_map_x_97_data_out:10'b0);
   assign  data_out240 = ((_net_1)?_add_map_x_97_data_out:10'b0)|
    ((_net_0)?_add_map_x_97_data_near:10'b0);
   assign  data_out241 = ((_net_1)?_add_map_x_98_data_near:10'b0)|
    ((_net_0)?_add_map_x_98_data_out:10'b0);
   assign  data_out242 = ((_net_1)?_add_map_x_98_data_out:10'b0)|
    ((_net_0)?_add_map_x_98_data_near:10'b0);
   assign  data_out243 = ((_net_1)?_add_map_x_99_data_near:10'b0)|
    ((_net_0)?_add_map_x_99_data_out:10'b0);
   assign  data_out244 = ((_net_1)?_add_map_x_99_data_out:10'b0)|
    ((_net_0)?_add_map_x_99_data_near:10'b0);
   assign  data_out245 = ((_net_1)?_add_map_x_100_data_near:10'b0)|
    ((_net_0)?_add_map_x_100_data_out:10'b0);
   assign  data_out246 = ((_net_1)?_add_map_x_100_data_out:10'b0)|
    ((_net_0)?_add_map_x_100_data_near:10'b0);
   assign  data_out247 = ((_net_1)?_add_map_x_101_data_near:10'b0)|
    ((_net_0)?_add_map_x_101_data_out:10'b0);
   assign  data_out248 = ((_net_1)?_add_map_x_101_data_out:10'b0)|
    ((_net_0)?_add_map_x_101_data_near:10'b0);
   assign  data_out249 = ((_net_1)?_add_map_x_102_data_near:10'b0)|
    ((_net_0)?_add_map_x_102_data_out:10'b0);
   assign  data_out250 = ((_net_1)?_add_map_x_102_data_out:10'b0)|
    ((_net_0)?_add_map_x_102_data_near:10'b0);
   assign  data_out251 = ((_net_1)?_add_map_x_103_data_near:10'b0)|
    ((_net_0)?_add_map_x_103_data_out:10'b0);
   assign  data_out252 = ((_net_1)?_add_map_x_103_data_out:10'b0)|
    ((_net_0)?_add_map_x_103_data_near:10'b0);
   assign  data_out253 = ((_net_1)?_add_map_x_104_data_near:10'b0)|
    ((_net_0)?_add_map_x_104_data_out:10'b0);
   assign  data_out254 = ((_net_1)?_add_map_x_104_data_out:10'b0)|
    ((_net_0)?_add_map_x_104_data_near:10'b0);
   assign  data_out257 = ((_net_1)?_add_map_x_105_data_out:10'b0)|
    ((_net_0)?_add_map_x_105_data_near:10'b0);
   assign  data_out258 = ((_net_1)?_add_map_x_105_data_near:10'b0)|
    ((_net_0)?_add_map_x_105_data_out:10'b0);
   assign  data_out259 = ((_net_1)?_add_map_x_106_data_out:10'b0)|
    ((_net_0)?_add_map_x_106_data_near:10'b0);
   assign  data_out260 = ((_net_1)?_add_map_x_106_data_near:10'b0)|
    ((_net_0)?_add_map_x_106_data_out:10'b0);
   assign  data_out261 = ((_net_1)?_add_map_x_107_data_out:10'b0)|
    ((_net_0)?_add_map_x_107_data_near:10'b0);
   assign  data_out262 = ((_net_1)?_add_map_x_107_data_near:10'b0)|
    ((_net_0)?_add_map_x_107_data_out:10'b0);
   assign  data_out263 = ((_net_1)?_add_map_x_108_data_out:10'b0)|
    ((_net_0)?_add_map_x_108_data_near:10'b0);
   assign  data_out264 = ((_net_1)?_add_map_x_108_data_near:10'b0)|
    ((_net_0)?_add_map_x_108_data_out:10'b0);
   assign  data_out265 = ((_net_1)?_add_map_x_109_data_out:10'b0)|
    ((_net_0)?_add_map_x_109_data_near:10'b0);
   assign  data_out266 = ((_net_1)?_add_map_x_109_data_near:10'b0)|
    ((_net_0)?_add_map_x_109_data_out:10'b0);
   assign  data_out267 = ((_net_1)?_add_map_x_110_data_out:10'b0)|
    ((_net_0)?_add_map_x_110_data_near:10'b0);
   assign  data_out268 = ((_net_1)?_add_map_x_110_data_near:10'b0)|
    ((_net_0)?_add_map_x_110_data_out:10'b0);
   assign  data_out269 = ((_net_1)?_add_map_x_111_data_out:10'b0)|
    ((_net_0)?_add_map_x_111_data_near:10'b0);
   assign  data_out270 = ((_net_1)?_add_map_x_111_data_near:10'b0)|
    ((_net_0)?_add_map_x_111_data_out:10'b0);
   assign  data_out271 = ((_net_1)?_add_map_x_112_data_out:10'b0)|
    ((_net_0)?_add_map_x_112_data_near:10'b0);
   assign  data_out272 = ((_net_1)?_add_map_x_112_data_near:10'b0)|
    ((_net_0)?_add_map_x_112_data_out:10'b0);
   assign  data_out273 = ((_net_1)?_add_map_x_113_data_out:10'b0)|
    ((_net_0)?_add_map_x_113_data_near:10'b0);
   assign  data_out274 = ((_net_1)?_add_map_x_113_data_near:10'b0)|
    ((_net_0)?_add_map_x_113_data_out:10'b0);
   assign  data_out275 = ((_net_1)?_add_map_x_114_data_out:10'b0)|
    ((_net_0)?_add_map_x_114_data_near:10'b0);
   assign  data_out276 = ((_net_1)?_add_map_x_114_data_near:10'b0)|
    ((_net_0)?_add_map_x_114_data_out:10'b0);
   assign  data_out277 = ((_net_1)?_add_map_x_115_data_out:10'b0)|
    ((_net_0)?_add_map_x_115_data_near:10'b0);
   assign  data_out278 = ((_net_1)?_add_map_x_115_data_near:10'b0)|
    ((_net_0)?_add_map_x_115_data_out:10'b0);
   assign  data_out279 = ((_net_1)?_add_map_x_116_data_out:10'b0)|
    ((_net_0)?_add_map_x_116_data_near:10'b0);
   assign  data_out280 = ((_net_1)?_add_map_x_116_data_near:10'b0)|
    ((_net_0)?_add_map_x_116_data_out:10'b0);
   assign  data_out281 = ((_net_1)?_add_map_x_117_data_out:10'b0)|
    ((_net_0)?_add_map_x_117_data_near:10'b0);
   assign  data_out282 = ((_net_1)?_add_map_x_117_data_near:10'b0)|
    ((_net_0)?_add_map_x_117_data_out:10'b0);
   assign  data_out283 = ((_net_1)?_add_map_x_118_data_out:10'b0)|
    ((_net_0)?_add_map_x_118_data_near:10'b0);
   assign  data_out284 = ((_net_1)?_add_map_x_118_data_near:10'b0)|
    ((_net_0)?_add_map_x_118_data_out:10'b0);
   assign  data_out285 = ((_net_1)?_add_map_x_119_data_out:10'b0)|
    ((_net_0)?_add_map_x_119_data_near:10'b0);
   assign  data_out286 = ((_net_1)?_add_map_x_119_data_near:10'b0)|
    ((_net_0)?_add_map_x_119_data_out:10'b0);
   assign  data_out289 = ((_net_1)?_add_map_x_120_data_near:10'b0)|
    ((_net_0)?_add_map_x_120_data_out:10'b0);
   assign  data_out290 = ((_net_1)?_add_map_x_120_data_out:10'b0)|
    ((_net_0)?_add_map_x_120_data_near:10'b0);
   assign  data_out291 = ((_net_1)?_add_map_x_121_data_near:10'b0)|
    ((_net_0)?_add_map_x_121_data_out:10'b0);
   assign  data_out292 = ((_net_1)?_add_map_x_121_data_out:10'b0)|
    ((_net_0)?_add_map_x_121_data_near:10'b0);
   assign  data_out293 = ((_net_1)?_add_map_x_122_data_near:10'b0)|
    ((_net_0)?_add_map_x_122_data_out:10'b0);
   assign  data_out294 = ((_net_1)?_add_map_x_122_data_out:10'b0)|
    ((_net_0)?_add_map_x_122_data_near:10'b0);
   assign  data_out295 = ((_net_1)?_add_map_x_123_data_near:10'b0)|
    ((_net_0)?_add_map_x_123_data_out:10'b0);
   assign  data_out296 = ((_net_1)?_add_map_x_123_data_out:10'b0)|
    ((_net_0)?_add_map_x_123_data_near:10'b0);
   assign  data_out297 = ((_net_1)?_add_map_x_124_data_near:10'b0)|
    ((_net_0)?_add_map_x_124_data_out:10'b0);
   assign  data_out298 = ((_net_1)?_add_map_x_124_data_out:10'b0)|
    ((_net_0)?_add_map_x_124_data_near:10'b0);
   assign  data_out299 = ((_net_1)?_add_map_x_125_data_near:10'b0)|
    ((_net_0)?_add_map_x_125_data_out:10'b0);
   assign  data_out300 = ((_net_1)?_add_map_x_125_data_out:10'b0)|
    ((_net_0)?_add_map_x_125_data_near:10'b0);
   assign  data_out301 = ((_net_1)?_add_map_x_126_data_near:10'b0)|
    ((_net_0)?_add_map_x_126_data_out:10'b0);
   assign  data_out302 = ((_net_1)?_add_map_x_126_data_out:10'b0)|
    ((_net_0)?_add_map_x_126_data_near:10'b0);
   assign  data_out303 = ((_net_1)?_add_map_x_127_data_near:10'b0)|
    ((_net_0)?_add_map_x_127_data_out:10'b0);
   assign  data_out304 = ((_net_1)?_add_map_x_127_data_out:10'b0)|
    ((_net_0)?_add_map_x_127_data_near:10'b0);
   assign  data_out305 = ((_net_1)?_add_map_x_128_data_near:10'b0)|
    ((_net_0)?_add_map_x_128_data_out:10'b0);
   assign  data_out306 = ((_net_1)?_add_map_x_128_data_out:10'b0)|
    ((_net_0)?_add_map_x_128_data_near:10'b0);
   assign  data_out307 = ((_net_1)?_add_map_x_129_data_near:10'b0)|
    ((_net_0)?_add_map_x_129_data_out:10'b0);
   assign  data_out308 = ((_net_1)?_add_map_x_129_data_out:10'b0)|
    ((_net_0)?_add_map_x_129_data_near:10'b0);
   assign  data_out309 = ((_net_1)?_add_map_x_130_data_near:10'b0)|
    ((_net_0)?_add_map_x_130_data_out:10'b0);
   assign  data_out310 = ((_net_1)?_add_map_x_130_data_out:10'b0)|
    ((_net_0)?_add_map_x_130_data_near:10'b0);
   assign  data_out311 = ((_net_1)?_add_map_x_131_data_near:10'b0)|
    ((_net_0)?_add_map_x_131_data_out:10'b0);
   assign  data_out312 = ((_net_1)?_add_map_x_131_data_out:10'b0)|
    ((_net_0)?_add_map_x_131_data_near:10'b0);
   assign  data_out313 = ((_net_1)?_add_map_x_132_data_near:10'b0)|
    ((_net_0)?_add_map_x_132_data_out:10'b0);
   assign  data_out314 = ((_net_1)?_add_map_x_132_data_out:10'b0)|
    ((_net_0)?_add_map_x_132_data_near:10'b0);
   assign  data_out315 = ((_net_1)?_add_map_x_133_data_near:10'b0)|
    ((_net_0)?_add_map_x_133_data_out:10'b0);
   assign  data_out316 = ((_net_1)?_add_map_x_133_data_out:10'b0)|
    ((_net_0)?_add_map_x_133_data_near:10'b0);
   assign  data_out317 = ((_net_1)?_add_map_x_134_data_near:10'b0)|
    ((_net_0)?_add_map_x_134_data_out:10'b0);
   assign  data_out318 = ((_net_1)?_add_map_x_134_data_out:10'b0)|
    ((_net_0)?_add_map_x_134_data_near:10'b0);
   assign  data_out321 = ((_net_1)?_add_map_x_135_data_out:10'b0)|
    ((_net_0)?_add_map_x_135_data_near:10'b0);
   assign  data_out322 = ((_net_1)?_add_map_x_135_data_near:10'b0)|
    ((_net_0)?_add_map_x_135_data_out:10'b0);
   assign  data_out323 = ((_net_1)?_add_map_x_136_data_out:10'b0)|
    ((_net_0)?_add_map_x_136_data_near:10'b0);
   assign  data_out324 = ((_net_1)?_add_map_x_136_data_near:10'b0)|
    ((_net_0)?_add_map_x_136_data_out:10'b0);
   assign  data_out325 = ((_net_1)?_add_map_x_137_data_out:10'b0)|
    ((_net_0)?_add_map_x_137_data_near:10'b0);
   assign  data_out326 = ((_net_1)?_add_map_x_137_data_near:10'b0)|
    ((_net_0)?_add_map_x_137_data_out:10'b0);
   assign  data_out327 = ((_net_1)?_add_map_x_138_data_out:10'b0)|
    ((_net_0)?_add_map_x_138_data_near:10'b0);
   assign  data_out328 = ((_net_1)?_add_map_x_138_data_near:10'b0)|
    ((_net_0)?_add_map_x_138_data_out:10'b0);
   assign  data_out329 = ((_net_1)?_add_map_x_139_data_out:10'b0)|
    ((_net_0)?_add_map_x_139_data_near:10'b0);
   assign  data_out330 = ((_net_1)?_add_map_x_139_data_near:10'b0)|
    ((_net_0)?_add_map_x_139_data_out:10'b0);
   assign  data_out331 = ((_net_1)?_add_map_x_140_data_out:10'b0)|
    ((_net_0)?_add_map_x_140_data_near:10'b0);
   assign  data_out332 = ((_net_1)?_add_map_x_140_data_near:10'b0)|
    ((_net_0)?_add_map_x_140_data_out:10'b0);
   assign  data_out333 = ((_net_1)?_add_map_x_141_data_out:10'b0)|
    ((_net_0)?_add_map_x_141_data_near:10'b0);
   assign  data_out334 = ((_net_1)?_add_map_x_141_data_near:10'b0)|
    ((_net_0)?_add_map_x_141_data_out:10'b0);
   assign  data_out335 = ((_net_1)?_add_map_x_142_data_out:10'b0)|
    ((_net_0)?_add_map_x_142_data_near:10'b0);
   assign  data_out336 = ((_net_1)?_add_map_x_142_data_near:10'b0)|
    ((_net_0)?_add_map_x_142_data_out:10'b0);
   assign  data_out337 = ((_net_1)?_add_map_x_143_data_out:10'b0)|
    ((_net_0)?_add_map_x_143_data_near:10'b0);
   assign  data_out338 = ((_net_1)?_add_map_x_143_data_near:10'b0)|
    ((_net_0)?_add_map_x_143_data_out:10'b0);
   assign  data_out339 = ((_net_1)?_add_map_x_144_data_out:10'b0)|
    ((_net_0)?_add_map_x_144_data_near:10'b0);
   assign  data_out340 = ((_net_1)?_add_map_x_144_data_near:10'b0)|
    ((_net_0)?_add_map_x_144_data_out:10'b0);
   assign  data_out341 = ((_net_1)?_add_map_x_145_data_out:10'b0)|
    ((_net_0)?_add_map_x_145_data_near:10'b0);
   assign  data_out342 = ((_net_1)?_add_map_x_145_data_near:10'b0)|
    ((_net_0)?_add_map_x_145_data_out:10'b0);
   assign  data_out343 = ((_net_1)?_add_map_x_146_data_out:10'b0)|
    ((_net_0)?_add_map_x_146_data_near:10'b0);
   assign  data_out344 = ((_net_1)?_add_map_x_146_data_near:10'b0)|
    ((_net_0)?_add_map_x_146_data_out:10'b0);
   assign  data_out345 = ((_net_1)?_add_map_x_147_data_out:10'b0)|
    ((_net_0)?_add_map_x_147_data_near:10'b0);
   assign  data_out346 = ((_net_1)?_add_map_x_147_data_near:10'b0)|
    ((_net_0)?_add_map_x_147_data_out:10'b0);
   assign  data_out347 = ((_net_1)?_add_map_x_148_data_out:10'b0)|
    ((_net_0)?_add_map_x_148_data_near:10'b0);
   assign  data_out348 = ((_net_1)?_add_map_x_148_data_near:10'b0)|
    ((_net_0)?_add_map_x_148_data_out:10'b0);
   assign  data_out349 = ((_net_1)?_add_map_x_149_data_out:10'b0)|
    ((_net_0)?_add_map_x_149_data_near:10'b0);
   assign  data_out350 = ((_net_1)?_add_map_x_149_data_near:10'b0)|
    ((_net_0)?_add_map_x_149_data_out:10'b0);
   assign  data_out353 = ((_net_1)?_add_map_x_150_data_near:10'b0)|
    ((_net_0)?_add_map_x_150_data_out:10'b0);
   assign  data_out354 = ((_net_1)?_add_map_x_150_data_out:10'b0)|
    ((_net_0)?_add_map_x_150_data_near:10'b0);
   assign  data_out355 = ((_net_1)?_add_map_x_151_data_near:10'b0)|
    ((_net_0)?_add_map_x_151_data_out:10'b0);
   assign  data_out356 = ((_net_1)?_add_map_x_151_data_out:10'b0)|
    ((_net_0)?_add_map_x_151_data_near:10'b0);
   assign  data_out357 = ((_net_1)?_add_map_x_152_data_near:10'b0)|
    ((_net_0)?_add_map_x_152_data_out:10'b0);
   assign  data_out358 = ((_net_1)?_add_map_x_152_data_out:10'b0)|
    ((_net_0)?_add_map_x_152_data_near:10'b0);
   assign  data_out359 = ((_net_1)?_add_map_x_153_data_near:10'b0)|
    ((_net_0)?_add_map_x_153_data_out:10'b0);
   assign  data_out360 = ((_net_1)?_add_map_x_153_data_out:10'b0)|
    ((_net_0)?_add_map_x_153_data_near:10'b0);
   assign  data_out361 = ((_net_1)?_add_map_x_154_data_near:10'b0)|
    ((_net_0)?_add_map_x_154_data_out:10'b0);
   assign  data_out362 = ((_net_1)?_add_map_x_154_data_out:10'b0)|
    ((_net_0)?_add_map_x_154_data_near:10'b0);
   assign  data_out363 = ((_net_1)?_add_map_x_155_data_near:10'b0)|
    ((_net_0)?_add_map_x_155_data_out:10'b0);
   assign  data_out364 = ((_net_1)?_add_map_x_155_data_out:10'b0)|
    ((_net_0)?_add_map_x_155_data_near:10'b0);
   assign  data_out365 = ((_net_1)?_add_map_x_156_data_near:10'b0)|
    ((_net_0)?_add_map_x_156_data_out:10'b0);
   assign  data_out366 = ((_net_1)?_add_map_x_156_data_out:10'b0)|
    ((_net_0)?_add_map_x_156_data_near:10'b0);
   assign  data_out367 = ((_net_1)?_add_map_x_157_data_near:10'b0)|
    ((_net_0)?_add_map_x_157_data_out:10'b0);
   assign  data_out368 = ((_net_1)?_add_map_x_157_data_out:10'b0)|
    ((_net_0)?_add_map_x_157_data_near:10'b0);
   assign  data_out369 = ((_net_1)?_add_map_x_158_data_near:10'b0)|
    ((_net_0)?_add_map_x_158_data_out:10'b0);
   assign  data_out370 = ((_net_1)?_add_map_x_158_data_out:10'b0)|
    ((_net_0)?_add_map_x_158_data_near:10'b0);
   assign  data_out371 = ((_net_1)?_add_map_x_159_data_near:10'b0)|
    ((_net_0)?_add_map_x_159_data_out:10'b0);
   assign  data_out372 = ((_net_1)?_add_map_x_159_data_out:10'b0)|
    ((_net_0)?_add_map_x_159_data_near:10'b0);
   assign  data_out373 = ((_net_1)?_add_map_x_160_data_near:10'b0)|
    ((_net_0)?_add_map_x_160_data_out:10'b0);
   assign  data_out374 = ((_net_1)?_add_map_x_160_data_out:10'b0)|
    ((_net_0)?_add_map_x_160_data_near:10'b0);
   assign  data_out375 = ((_net_1)?_add_map_x_161_data_near:10'b0)|
    ((_net_0)?_add_map_x_161_data_out:10'b0);
   assign  data_out376 = ((_net_1)?_add_map_x_161_data_out:10'b0)|
    ((_net_0)?_add_map_x_161_data_near:10'b0);
   assign  data_out377 = ((_net_1)?_add_map_x_162_data_near:10'b0)|
    ((_net_0)?_add_map_x_162_data_out:10'b0);
   assign  data_out378 = ((_net_1)?_add_map_x_162_data_out:10'b0)|
    ((_net_0)?_add_map_x_162_data_near:10'b0);
   assign  data_out379 = ((_net_1)?_add_map_x_163_data_near:10'b0)|
    ((_net_0)?_add_map_x_163_data_out:10'b0);
   assign  data_out380 = ((_net_1)?_add_map_x_163_data_out:10'b0)|
    ((_net_0)?_add_map_x_163_data_near:10'b0);
   assign  data_out381 = ((_net_1)?_add_map_x_164_data_near:10'b0)|
    ((_net_0)?_add_map_x_164_data_out:10'b0);
   assign  data_out382 = ((_net_1)?_add_map_x_164_data_out:10'b0)|
    ((_net_0)?_add_map_x_164_data_near:10'b0);
   assign  data_out385 = ((_net_1)?_add_map_x_165_data_out:10'b0)|
    ((_net_0)?_add_map_x_165_data_near:10'b0);
   assign  data_out386 = ((_net_1)?_add_map_x_165_data_near:10'b0)|
    ((_net_0)?_add_map_x_165_data_out:10'b0);
   assign  data_out387 = ((_net_1)?_add_map_x_166_data_out:10'b0)|
    ((_net_0)?_add_map_x_166_data_near:10'b0);
   assign  data_out388 = ((_net_1)?_add_map_x_166_data_near:10'b0)|
    ((_net_0)?_add_map_x_166_data_out:10'b0);
   assign  data_out389 = ((_net_1)?_add_map_x_167_data_out:10'b0)|
    ((_net_0)?_add_map_x_167_data_near:10'b0);
   assign  data_out390 = ((_net_1)?_add_map_x_167_data_near:10'b0)|
    ((_net_0)?_add_map_x_167_data_out:10'b0);
   assign  data_out391 = ((_net_1)?_add_map_x_168_data_out:10'b0)|
    ((_net_0)?_add_map_x_168_data_near:10'b0);
   assign  data_out392 = ((_net_1)?_add_map_x_168_data_near:10'b0)|
    ((_net_0)?_add_map_x_168_data_out:10'b0);
   assign  data_out393 = ((_net_1)?_add_map_x_169_data_out:10'b0)|
    ((_net_0)?_add_map_x_169_data_near:10'b0);
   assign  data_out394 = ((_net_1)?_add_map_x_169_data_near:10'b0)|
    ((_net_0)?_add_map_x_169_data_out:10'b0);
   assign  data_out395 = ((_net_1)?_add_map_x_170_data_out:10'b0)|
    ((_net_0)?_add_map_x_170_data_near:10'b0);
   assign  data_out396 = ((_net_1)?_add_map_x_170_data_near:10'b0)|
    ((_net_0)?_add_map_x_170_data_out:10'b0);
   assign  data_out397 = ((_net_1)?_add_map_x_171_data_out:10'b0)|
    ((_net_0)?_add_map_x_171_data_near:10'b0);
   assign  data_out398 = ((_net_1)?_add_map_x_171_data_near:10'b0)|
    ((_net_0)?_add_map_x_171_data_out:10'b0);
   assign  data_out399 = ((_net_1)?_add_map_x_172_data_out:10'b0)|
    ((_net_0)?_add_map_x_172_data_near:10'b0);
   assign  data_out400 = ((_net_1)?_add_map_x_172_data_near:10'b0)|
    ((_net_0)?_add_map_x_172_data_out:10'b0);
   assign  data_out401 = ((_net_1)?_add_map_x_173_data_out:10'b0)|
    ((_net_0)?_add_map_x_173_data_near:10'b0);
   assign  data_out402 = ((_net_1)?_add_map_x_173_data_near:10'b0)|
    ((_net_0)?_add_map_x_173_data_out:10'b0);
   assign  data_out403 = ((_net_1)?_add_map_x_174_data_out:10'b0)|
    ((_net_0)?_add_map_x_174_data_near:10'b0);
   assign  data_out404 = ((_net_1)?_add_map_x_174_data_near:10'b0)|
    ((_net_0)?_add_map_x_174_data_out:10'b0);
   assign  data_out405 = ((_net_1)?_add_map_x_175_data_out:10'b0)|
    ((_net_0)?_add_map_x_175_data_near:10'b0);
   assign  data_out406 = ((_net_1)?_add_map_x_175_data_near:10'b0)|
    ((_net_0)?_add_map_x_175_data_out:10'b0);
   assign  data_out407 = ((_net_1)?_add_map_x_176_data_out:10'b0)|
    ((_net_0)?_add_map_x_176_data_near:10'b0);
   assign  data_out408 = ((_net_1)?_add_map_x_176_data_near:10'b0)|
    ((_net_0)?_add_map_x_176_data_out:10'b0);
   assign  data_out409 = ((_net_1)?_add_map_x_177_data_out:10'b0)|
    ((_net_0)?_add_map_x_177_data_near:10'b0);
   assign  data_out410 = ((_net_1)?_add_map_x_177_data_near:10'b0)|
    ((_net_0)?_add_map_x_177_data_out:10'b0);
   assign  data_out411 = ((_net_1)?_add_map_x_178_data_out:10'b0)|
    ((_net_0)?_add_map_x_178_data_near:10'b0);
   assign  data_out412 = ((_net_1)?_add_map_x_178_data_near:10'b0)|
    ((_net_0)?_add_map_x_178_data_out:10'b0);
   assign  data_out413 = ((_net_1)?_add_map_x_179_data_out:10'b0)|
    ((_net_0)?_add_map_x_179_data_near:10'b0);
   assign  data_out414 = ((_net_1)?_add_map_x_179_data_near:10'b0)|
    ((_net_0)?_add_map_x_179_data_out:10'b0);
   assign  data_out417 = ((_net_1)?_add_map_x_180_data_near:10'b0)|
    ((_net_0)?_add_map_x_180_data_out:10'b0);
   assign  data_out418 = ((_net_1)?_add_map_x_180_data_out:10'b0)|
    ((_net_0)?_add_map_x_180_data_near:10'b0);
   assign  data_out419 = ((_net_1)?_add_map_x_181_data_near:10'b0)|
    ((_net_0)?_add_map_x_181_data_out:10'b0);
   assign  data_out420 = ((_net_1)?_add_map_x_181_data_out:10'b0)|
    ((_net_0)?_add_map_x_181_data_near:10'b0);
   assign  data_out421 = ((_net_1)?_add_map_x_182_data_near:10'b0)|
    ((_net_0)?_add_map_x_182_data_out:10'b0);
   assign  data_out422 = ((_net_1)?_add_map_x_182_data_out:10'b0)|
    ((_net_0)?_add_map_x_182_data_near:10'b0);
   assign  data_out423 = ((_net_1)?_add_map_x_183_data_near:10'b0)|
    ((_net_0)?_add_map_x_183_data_out:10'b0);
   assign  data_out424 = ((_net_1)?_add_map_x_183_data_out:10'b0)|
    ((_net_0)?_add_map_x_183_data_near:10'b0);
   assign  data_out425 = ((_net_1)?_add_map_x_184_data_near:10'b0)|
    ((_net_0)?_add_map_x_184_data_out:10'b0);
   assign  data_out426 = ((_net_1)?_add_map_x_184_data_out:10'b0)|
    ((_net_0)?_add_map_x_184_data_near:10'b0);
   assign  data_out427 = ((_net_1)?_add_map_x_185_data_near:10'b0)|
    ((_net_0)?_add_map_x_185_data_out:10'b0);
   assign  data_out428 = ((_net_1)?_add_map_x_185_data_out:10'b0)|
    ((_net_0)?_add_map_x_185_data_near:10'b0);
   assign  data_out429 = ((_net_1)?_add_map_x_186_data_near:10'b0)|
    ((_net_0)?_add_map_x_186_data_out:10'b0);
   assign  data_out430 = ((_net_1)?_add_map_x_186_data_out:10'b0)|
    ((_net_0)?_add_map_x_186_data_near:10'b0);
   assign  data_out431 = ((_net_1)?_add_map_x_187_data_near:10'b0)|
    ((_net_0)?_add_map_x_187_data_out:10'b0);
   assign  data_out432 = ((_net_1)?_add_map_x_187_data_out:10'b0)|
    ((_net_0)?_add_map_x_187_data_near:10'b0);
   assign  data_out433 = ((_net_1)?_add_map_x_188_data_near:10'b0)|
    ((_net_0)?_add_map_x_188_data_out:10'b0);
   assign  data_out434 = ((_net_1)?_add_map_x_188_data_out:10'b0)|
    ((_net_0)?_add_map_x_188_data_near:10'b0);
   assign  data_out435 = ((_net_1)?_add_map_x_189_data_near:10'b0)|
    ((_net_0)?_add_map_x_189_data_out:10'b0);
   assign  data_out436 = ((_net_1)?_add_map_x_189_data_out:10'b0)|
    ((_net_0)?_add_map_x_189_data_near:10'b0);
   assign  data_out437 = ((_net_1)?_add_map_x_190_data_near:10'b0)|
    ((_net_0)?_add_map_x_190_data_out:10'b0);
   assign  data_out438 = ((_net_1)?_add_map_x_190_data_out:10'b0)|
    ((_net_0)?_add_map_x_190_data_near:10'b0);
   assign  data_out439 = ((_net_1)?_add_map_x_191_data_near:10'b0)|
    ((_net_0)?_add_map_x_191_data_out:10'b0);
   assign  data_out440 = ((_net_1)?_add_map_x_191_data_out:10'b0)|
    ((_net_0)?_add_map_x_191_data_near:10'b0);
   assign  data_out441 = ((_net_1)?_add_map_x_192_data_near:10'b0)|
    ((_net_0)?_add_map_x_192_data_out:10'b0);
   assign  data_out442 = ((_net_1)?_add_map_x_192_data_out:10'b0)|
    ((_net_0)?_add_map_x_192_data_near:10'b0);
   assign  data_out443 = ((_net_1)?_add_map_x_193_data_near:10'b0)|
    ((_net_0)?_add_map_x_193_data_out:10'b0);
   assign  data_out444 = ((_net_1)?_add_map_x_193_data_out:10'b0)|
    ((_net_0)?_add_map_x_193_data_near:10'b0);
   assign  data_out445 = ((_net_1)?_add_map_x_194_data_near:10'b0)|
    ((_net_0)?_add_map_x_194_data_out:10'b0);
   assign  data_out446 = ((_net_1)?_add_map_x_194_data_out:10'b0)|
    ((_net_0)?_add_map_x_194_data_near:10'b0);
   assign  data_out449 = ((_net_1)?_add_map_x_195_data_out:10'b0)|
    ((_net_0)?_add_map_x_195_data_near:10'b0);
   assign  data_out450 = ((_net_1)?_add_map_x_195_data_near:10'b0)|
    ((_net_0)?_add_map_x_195_data_out:10'b0);
   assign  data_out451 = ((_net_1)?_add_map_x_196_data_out:10'b0)|
    ((_net_0)?_add_map_x_196_data_near:10'b0);
   assign  data_out452 = ((_net_1)?_add_map_x_196_data_near:10'b0)|
    ((_net_0)?_add_map_x_196_data_out:10'b0);
   assign  data_out453 = ((_net_1)?_add_map_x_197_data_out:10'b0)|
    ((_net_0)?_add_map_x_197_data_near:10'b0);
   assign  data_out454 = ((_net_1)?_add_map_x_197_data_near:10'b0)|
    ((_net_0)?_add_map_x_197_data_out:10'b0);
   assign  data_out455 = ((_net_1)?_add_map_x_198_data_out:10'b0)|
    ((_net_0)?_add_map_x_198_data_near:10'b0);
   assign  data_out456 = ((_net_1)?_add_map_x_198_data_near:10'b0)|
    ((_net_0)?_add_map_x_198_data_out:10'b0);
   assign  data_out457 = ((_net_1)?_add_map_x_199_data_out:10'b0)|
    ((_net_0)?_add_map_x_199_data_near:10'b0);
   assign  data_out458 = ((_net_1)?_add_map_x_199_data_near:10'b0)|
    ((_net_0)?_add_map_x_199_data_out:10'b0);
   assign  data_out459 = ((_net_1)?_add_map_x_200_data_out:10'b0)|
    ((_net_0)?_add_map_x_200_data_near:10'b0);
   assign  data_out460 = ((_net_1)?_add_map_x_200_data_near:10'b0)|
    ((_net_0)?_add_map_x_200_data_out:10'b0);
   assign  data_out461 = ((_net_1)?_add_map_x_201_data_out:10'b0)|
    ((_net_0)?_add_map_x_201_data_near:10'b0);
   assign  data_out462 = ((_net_1)?_add_map_x_201_data_near:10'b0)|
    ((_net_0)?_add_map_x_201_data_out:10'b0);
   assign  data_out463 = ((_net_1)?_add_map_x_202_data_out:10'b0)|
    ((_net_0)?_add_map_x_202_data_near:10'b0);
   assign  data_out464 = ((_net_1)?_add_map_x_202_data_near:10'b0)|
    ((_net_0)?_add_map_x_202_data_out:10'b0);
   assign  data_out465 = ((_net_1)?_add_map_x_203_data_out:10'b0)|
    ((_net_0)?_add_map_x_203_data_near:10'b0);
   assign  data_out466 = ((_net_1)?_add_map_x_203_data_near:10'b0)|
    ((_net_0)?_add_map_x_203_data_out:10'b0);
   assign  data_out467 = ((_net_1)?_add_map_x_204_data_out:10'b0)|
    ((_net_0)?_add_map_x_204_data_near:10'b0);
   assign  data_out468 = ((_net_1)?_add_map_x_204_data_near:10'b0)|
    ((_net_0)?_add_map_x_204_data_out:10'b0);
   assign  data_out469 = ((_net_1)?_add_map_x_205_data_out:10'b0)|
    ((_net_0)?_add_map_x_205_data_near:10'b0);
   assign  data_out470 = ((_net_1)?_add_map_x_205_data_near:10'b0)|
    ((_net_0)?_add_map_x_205_data_out:10'b0);
   assign  data_out471 = ((_net_1)?_add_map_x_206_data_out:10'b0)|
    ((_net_0)?_add_map_x_206_data_near:10'b0);
   assign  data_out472 = ((_net_1)?_add_map_x_206_data_near:10'b0)|
    ((_net_0)?_add_map_x_206_data_out:10'b0);
   assign  data_out473 = ((_net_1)?_add_map_x_207_data_out:10'b0)|
    ((_net_0)?_add_map_x_207_data_near:10'b0);
   assign  data_out474 = ((_net_1)?_add_map_x_207_data_near:10'b0)|
    ((_net_0)?_add_map_x_207_data_out:10'b0);
   assign  data_out475 = ((_net_1)?_add_map_x_208_data_out:10'b0)|
    ((_net_0)?_add_map_x_208_data_near:10'b0);
   assign  data_out476 = ((_net_1)?_add_map_x_208_data_near:10'b0)|
    ((_net_0)?_add_map_x_208_data_out:10'b0);
   assign  data_out477 = ((_net_1)?_add_map_x_209_data_out:10'b0)|
    ((_net_0)?_add_map_x_209_data_near:10'b0);
   assign  data_out478 = ((_net_1)?_add_map_x_209_data_near:10'b0)|
    ((_net_0)?_add_map_x_209_data_out:10'b0);
   assign  data_out_index33 = ((_net_1)?_add_map_x_data_near:10'b0)|
    ((_net_0)?_add_map_x_data_out_index:10'b0);
   assign  data_out_index34 = ((_net_1)?_add_map_x_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_data_near:10'b0);
   assign  data_out_index35 = ((_net_1)?_add_map_x_1_data_near:10'b0)|
    ((_net_0)?_add_map_x_1_data_out_index:10'b0);
   assign  data_out_index36 = ((_net_1)?_add_map_x_1_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_1_data_near:10'b0);
   assign  data_out_index37 = ((_net_1)?_add_map_x_2_data_near:10'b0)|
    ((_net_0)?_add_map_x_2_data_out_index:10'b0);
   assign  data_out_index38 = ((_net_1)?_add_map_x_2_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_2_data_near:10'b0);
   assign  data_out_index39 = ((_net_1)?_add_map_x_3_data_near:10'b0)|
    ((_net_0)?_add_map_x_3_data_out_index:10'b0);
   assign  data_out_index40 = ((_net_1)?_add_map_x_3_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_3_data_near:10'b0);
   assign  data_out_index41 = ((_net_1)?_add_map_x_4_data_near:10'b0)|
    ((_net_0)?_add_map_x_4_data_out_index:10'b0);
   assign  data_out_index42 = ((_net_1)?_add_map_x_4_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_4_data_near:10'b0);
   assign  data_out_index43 = ((_net_1)?_add_map_x_5_data_near:10'b0)|
    ((_net_0)?_add_map_x_5_data_out_index:10'b0);
   assign  data_out_index44 = ((_net_1)?_add_map_x_5_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_5_data_near:10'b0);
   assign  data_out_index45 = ((_net_1)?_add_map_x_6_data_near:10'b0)|
    ((_net_0)?_add_map_x_6_data_out_index:10'b0);
   assign  data_out_index46 = ((_net_1)?_add_map_x_6_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_6_data_near:10'b0);
   assign  data_out_index47 = ((_net_1)?_add_map_x_7_data_near:10'b0)|
    ((_net_0)?_add_map_x_7_data_out_index:10'b0);
   assign  data_out_index48 = ((_net_1)?_add_map_x_7_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_7_data_near:10'b0);
   assign  data_out_index49 = ((_net_1)?_add_map_x_8_data_near:10'b0)|
    ((_net_0)?_add_map_x_8_data_out_index:10'b0);
   assign  data_out_index50 = ((_net_1)?_add_map_x_8_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_8_data_near:10'b0);
   assign  data_out_index51 = ((_net_1)?_add_map_x_9_data_near:10'b0)|
    ((_net_0)?_add_map_x_9_data_out_index:10'b0);
   assign  data_out_index52 = ((_net_1)?_add_map_x_9_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_9_data_near:10'b0);
   assign  data_out_index53 = ((_net_1)?_add_map_x_10_data_near:10'b0)|
    ((_net_0)?_add_map_x_10_data_out_index:10'b0);
   assign  data_out_index54 = ((_net_1)?_add_map_x_10_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_10_data_near:10'b0);
   assign  data_out_index55 = ((_net_1)?_add_map_x_11_data_near:10'b0)|
    ((_net_0)?_add_map_x_11_data_out_index:10'b0);
   assign  data_out_index56 = ((_net_1)?_add_map_x_11_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_11_data_near:10'b0);
   assign  data_out_index57 = ((_net_1)?_add_map_x_12_data_near:10'b0)|
    ((_net_0)?_add_map_x_12_data_out_index:10'b0);
   assign  data_out_index58 = ((_net_1)?_add_map_x_12_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_12_data_near:10'b0);
   assign  data_out_index59 = ((_net_1)?_add_map_x_13_data_near:10'b0)|
    ((_net_0)?_add_map_x_13_data_out_index:10'b0);
   assign  data_out_index60 = ((_net_1)?_add_map_x_13_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_13_data_near:10'b0);
   assign  data_out_index61 = ((_net_1)?_add_map_x_14_data_near:10'b0)|
    ((_net_0)?_add_map_x_14_data_out_index:10'b0);
   assign  data_out_index62 = ((_net_1)?_add_map_x_14_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_14_data_near:10'b0);
   assign  data_out_index65 = ((_net_1)?_add_map_x_15_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_15_data_near:10'b0);
   assign  data_out_index66 = ((_net_1)?_add_map_x_15_data_near:10'b0)|
    ((_net_0)?_add_map_x_15_data_out_index:10'b0);
   assign  data_out_index67 = ((_net_1)?_add_map_x_16_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_16_data_near:10'b0);
   assign  data_out_index68 = ((_net_1)?_add_map_x_16_data_near:10'b0)|
    ((_net_0)?_add_map_x_16_data_out_index:10'b0);
   assign  data_out_index69 = ((_net_1)?_add_map_x_17_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_17_data_near:10'b0);
   assign  data_out_index70 = ((_net_1)?_add_map_x_17_data_near:10'b0)|
    ((_net_0)?_add_map_x_17_data_out_index:10'b0);
   assign  data_out_index71 = ((_net_1)?_add_map_x_18_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_18_data_near:10'b0);
   assign  data_out_index72 = ((_net_1)?_add_map_x_18_data_near:10'b0)|
    ((_net_0)?_add_map_x_18_data_out_index:10'b0);
   assign  data_out_index73 = ((_net_1)?_add_map_x_19_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_19_data_near:10'b0);
   assign  data_out_index74 = ((_net_1)?_add_map_x_19_data_near:10'b0)|
    ((_net_0)?_add_map_x_19_data_out_index:10'b0);
   assign  data_out_index75 = ((_net_1)?_add_map_x_20_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_20_data_near:10'b0);
   assign  data_out_index76 = ((_net_1)?_add_map_x_20_data_near:10'b0)|
    ((_net_0)?_add_map_x_20_data_out_index:10'b0);
   assign  data_out_index77 = ((_net_1)?_add_map_x_21_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_21_data_near:10'b0);
   assign  data_out_index78 = ((_net_1)?_add_map_x_21_data_near:10'b0)|
    ((_net_0)?_add_map_x_21_data_out_index:10'b0);
   assign  data_out_index79 = ((_net_1)?_add_map_x_22_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_22_data_near:10'b0);
   assign  data_out_index80 = ((_net_1)?_add_map_x_22_data_near:10'b0)|
    ((_net_0)?_add_map_x_22_data_out_index:10'b0);
   assign  data_out_index81 = ((_net_1)?_add_map_x_23_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_23_data_near:10'b0);
   assign  data_out_index82 = ((_net_1)?_add_map_x_23_data_near:10'b0)|
    ((_net_0)?_add_map_x_23_data_out_index:10'b0);
   assign  data_out_index83 = ((_net_1)?_add_map_x_24_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_24_data_near:10'b0);
   assign  data_out_index84 = ((_net_1)?_add_map_x_24_data_near:10'b0)|
    ((_net_0)?_add_map_x_24_data_out_index:10'b0);
   assign  data_out_index85 = ((_net_1)?_add_map_x_25_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_25_data_near:10'b0);
   assign  data_out_index86 = ((_net_1)?_add_map_x_25_data_near:10'b0)|
    ((_net_0)?_add_map_x_25_data_out_index:10'b0);
   assign  data_out_index87 = ((_net_1)?_add_map_x_26_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_26_data_near:10'b0);
   assign  data_out_index88 = ((_net_1)?_add_map_x_26_data_near:10'b0)|
    ((_net_0)?_add_map_x_26_data_out_index:10'b0);
   assign  data_out_index89 = ((_net_1)?_add_map_x_27_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_27_data_near:10'b0);
   assign  data_out_index90 = ((_net_1)?_add_map_x_27_data_near:10'b0)|
    ((_net_0)?_add_map_x_27_data_out_index:10'b0);
   assign  data_out_index91 = ((_net_1)?_add_map_x_28_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_28_data_near:10'b0);
   assign  data_out_index92 = ((_net_1)?_add_map_x_28_data_near:10'b0)|
    ((_net_0)?_add_map_x_28_data_out_index:10'b0);
   assign  data_out_index93 = ((_net_1)?_add_map_x_29_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_29_data_near:10'b0);
   assign  data_out_index94 = ((_net_1)?_add_map_x_29_data_near:10'b0)|
    ((_net_0)?_add_map_x_29_data_out_index:10'b0);
   assign  data_out_index97 = ((_net_1)?_add_map_x_30_data_near:10'b0)|
    ((_net_0)?_add_map_x_30_data_out_index:10'b0);
   assign  data_out_index98 = ((_net_1)?_add_map_x_30_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_30_data_near:10'b0);
   assign  data_out_index99 = ((_net_1)?_add_map_x_31_data_near:10'b0)|
    ((_net_0)?_add_map_x_31_data_out_index:10'b0);
   assign  data_out_index100 = ((_net_1)?_add_map_x_31_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_31_data_near:10'b0);
   assign  data_out_index101 = ((_net_1)?_add_map_x_32_data_near:10'b0)|
    ((_net_0)?_add_map_x_32_data_out_index:10'b0);
   assign  data_out_index102 = ((_net_1)?_add_map_x_32_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_32_data_near:10'b0);
   assign  data_out_index103 = ((_net_1)?_add_map_x_33_data_near:10'b0)|
    ((_net_0)?_add_map_x_33_data_out_index:10'b0);
   assign  data_out_index104 = ((_net_1)?_add_map_x_33_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_33_data_near:10'b0);
   assign  data_out_index105 = ((_net_1)?_add_map_x_34_data_near:10'b0)|
    ((_net_0)?_add_map_x_34_data_out_index:10'b0);
   assign  data_out_index106 = ((_net_1)?_add_map_x_34_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_34_data_near:10'b0);
   assign  data_out_index107 = ((_net_1)?_add_map_x_35_data_near:10'b0)|
    ((_net_0)?_add_map_x_35_data_out_index:10'b0);
   assign  data_out_index108 = ((_net_1)?_add_map_x_35_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_35_data_near:10'b0);
   assign  data_out_index109 = ((_net_1)?_add_map_x_36_data_near:10'b0)|
    ((_net_0)?_add_map_x_36_data_out_index:10'b0);
   assign  data_out_index110 = ((_net_1)?_add_map_x_36_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_36_data_near:10'b0);
   assign  data_out_index111 = ((_net_1)?_add_map_x_37_data_near:10'b0)|
    ((_net_0)?_add_map_x_37_data_out_index:10'b0);
   assign  data_out_index112 = ((_net_1)?_add_map_x_37_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_37_data_near:10'b0);
   assign  data_out_index113 = ((_net_1)?_add_map_x_38_data_near:10'b0)|
    ((_net_0)?_add_map_x_38_data_out_index:10'b0);
   assign  data_out_index114 = ((_net_1)?_add_map_x_38_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_38_data_near:10'b0);
   assign  data_out_index115 = ((_net_1)?_add_map_x_39_data_near:10'b0)|
    ((_net_0)?_add_map_x_39_data_out_index:10'b0);
   assign  data_out_index116 = ((_net_1)?_add_map_x_39_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_39_data_near:10'b0);
   assign  data_out_index117 = ((_net_1)?_add_map_x_40_data_near:10'b0)|
    ((_net_0)?_add_map_x_40_data_out_index:10'b0);
   assign  data_out_index118 = ((_net_1)?_add_map_x_40_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_40_data_near:10'b0);
   assign  data_out_index119 = ((_net_1)?_add_map_x_41_data_near:10'b0)|
    ((_net_0)?_add_map_x_41_data_out_index:10'b0);
   assign  data_out_index120 = ((_net_1)?_add_map_x_41_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_41_data_near:10'b0);
   assign  data_out_index121 = ((_net_1)?_add_map_x_42_data_near:10'b0)|
    ((_net_0)?_add_map_x_42_data_out_index:10'b0);
   assign  data_out_index122 = ((_net_1)?_add_map_x_42_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_42_data_near:10'b0);
   assign  data_out_index123 = ((_net_1)?_add_map_x_43_data_near:10'b0)|
    ((_net_0)?_add_map_x_43_data_out_index:10'b0);
   assign  data_out_index124 = ((_net_1)?_add_map_x_43_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_43_data_near:10'b0);
   assign  data_out_index125 = ((_net_1)?_add_map_x_44_data_near:10'b0)|
    ((_net_0)?_add_map_x_44_data_out_index:10'b0);
   assign  data_out_index126 = ((_net_1)?_add_map_x_44_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_44_data_near:10'b0);
   assign  data_out_index129 = ((_net_1)?_add_map_x_45_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_45_data_near:10'b0);
   assign  data_out_index130 = ((_net_1)?_add_map_x_45_data_near:10'b0)|
    ((_net_0)?_add_map_x_45_data_out_index:10'b0);
   assign  data_out_index131 = ((_net_1)?_add_map_x_46_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_46_data_near:10'b0);
   assign  data_out_index132 = ((_net_1)?_add_map_x_46_data_near:10'b0)|
    ((_net_0)?_add_map_x_46_data_out_index:10'b0);
   assign  data_out_index133 = ((_net_1)?_add_map_x_47_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_47_data_near:10'b0);
   assign  data_out_index134 = ((_net_1)?_add_map_x_47_data_near:10'b0)|
    ((_net_0)?_add_map_x_47_data_out_index:10'b0);
   assign  data_out_index135 = ((_net_1)?_add_map_x_48_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_48_data_near:10'b0);
   assign  data_out_index136 = ((_net_1)?_add_map_x_48_data_near:10'b0)|
    ((_net_0)?_add_map_x_48_data_out_index:10'b0);
   assign  data_out_index137 = ((_net_1)?_add_map_x_49_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_49_data_near:10'b0);
   assign  data_out_index138 = ((_net_1)?_add_map_x_49_data_near:10'b0)|
    ((_net_0)?_add_map_x_49_data_out_index:10'b0);
   assign  data_out_index139 = ((_net_1)?_add_map_x_50_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_50_data_near:10'b0);
   assign  data_out_index140 = ((_net_1)?_add_map_x_50_data_near:10'b0)|
    ((_net_0)?_add_map_x_50_data_out_index:10'b0);
   assign  data_out_index141 = ((_net_1)?_add_map_x_51_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_51_data_near:10'b0);
   assign  data_out_index142 = ((_net_1)?_add_map_x_51_data_near:10'b0)|
    ((_net_0)?_add_map_x_51_data_out_index:10'b0);
   assign  data_out_index143 = ((_net_1)?_add_map_x_52_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_52_data_near:10'b0);
   assign  data_out_index144 = ((_net_1)?_add_map_x_52_data_near:10'b0)|
    ((_net_0)?_add_map_x_52_data_out_index:10'b0);
   assign  data_out_index145 = ((_net_1)?_add_map_x_53_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_53_data_near:10'b0);
   assign  data_out_index146 = ((_net_1)?_add_map_x_53_data_near:10'b0)|
    ((_net_0)?_add_map_x_53_data_out_index:10'b0);
   assign  data_out_index147 = ((_net_1)?_add_map_x_54_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_54_data_near:10'b0);
   assign  data_out_index148 = ((_net_1)?_add_map_x_54_data_near:10'b0)|
    ((_net_0)?_add_map_x_54_data_out_index:10'b0);
   assign  data_out_index149 = ((_net_1)?_add_map_x_55_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_55_data_near:10'b0);
   assign  data_out_index150 = ((_net_1)?_add_map_x_55_data_near:10'b0)|
    ((_net_0)?_add_map_x_55_data_out_index:10'b0);
   assign  data_out_index151 = ((_net_1)?_add_map_x_56_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_56_data_near:10'b0);
   assign  data_out_index152 = ((_net_1)?_add_map_x_56_data_near:10'b0)|
    ((_net_0)?_add_map_x_56_data_out_index:10'b0);
   assign  data_out_index153 = ((_net_1)?_add_map_x_57_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_57_data_near:10'b0);
   assign  data_out_index154 = ((_net_1)?_add_map_x_57_data_near:10'b0)|
    ((_net_0)?_add_map_x_57_data_out_index:10'b0);
   assign  data_out_index155 = ((_net_1)?_add_map_x_58_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_58_data_near:10'b0);
   assign  data_out_index156 = ((_net_1)?_add_map_x_58_data_near:10'b0)|
    ((_net_0)?_add_map_x_58_data_out_index:10'b0);
   assign  data_out_index157 = ((_net_1)?_add_map_x_59_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_59_data_near:10'b0);
   assign  data_out_index158 = ((_net_1)?_add_map_x_59_data_near:10'b0)|
    ((_net_0)?_add_map_x_59_data_out_index:10'b0);
   assign  data_out_index161 = ((_net_1)?_add_map_x_60_data_near:10'b0)|
    ((_net_0)?_add_map_x_60_data_out_index:10'b0);
   assign  data_out_index162 = ((_net_1)?_add_map_x_60_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_60_data_near:10'b0);
   assign  data_out_index163 = ((_net_1)?_add_map_x_61_data_near:10'b0)|
    ((_net_0)?_add_map_x_61_data_out_index:10'b0);
   assign  data_out_index164 = ((_net_1)?_add_map_x_61_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_61_data_near:10'b0);
   assign  data_out_index165 = ((_net_1)?_add_map_x_62_data_near:10'b0)|
    ((_net_0)?_add_map_x_62_data_out_index:10'b0);
   assign  data_out_index166 = ((_net_1)?_add_map_x_62_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_62_data_near:10'b0);
   assign  data_out_index167 = ((_net_1)?_add_map_x_63_data_near:10'b0)|
    ((_net_0)?_add_map_x_63_data_out_index:10'b0);
   assign  data_out_index168 = ((_net_1)?_add_map_x_63_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_63_data_near:10'b0);
   assign  data_out_index169 = ((_net_1)?_add_map_x_64_data_near:10'b0)|
    ((_net_0)?_add_map_x_64_data_out_index:10'b0);
   assign  data_out_index170 = ((_net_1)?_add_map_x_64_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_64_data_near:10'b0);
   assign  data_out_index171 = ((_net_1)?_add_map_x_65_data_near:10'b0)|
    ((_net_0)?_add_map_x_65_data_out_index:10'b0);
   assign  data_out_index172 = ((_net_1)?_add_map_x_65_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_65_data_near:10'b0);
   assign  data_out_index173 = ((_net_1)?_add_map_x_66_data_near:10'b0)|
    ((_net_0)?_add_map_x_66_data_out_index:10'b0);
   assign  data_out_index174 = ((_net_1)?_add_map_x_66_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_66_data_near:10'b0);
   assign  data_out_index175 = ((_net_1)?_add_map_x_67_data_near:10'b0)|
    ((_net_0)?_add_map_x_67_data_out_index:10'b0);
   assign  data_out_index176 = ((_net_1)?_add_map_x_67_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_67_data_near:10'b0);
   assign  data_out_index177 = ((_net_1)?_add_map_x_68_data_near:10'b0)|
    ((_net_0)?_add_map_x_68_data_out_index:10'b0);
   assign  data_out_index178 = ((_net_1)?_add_map_x_68_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_68_data_near:10'b0);
   assign  data_out_index179 = ((_net_1)?_add_map_x_69_data_near:10'b0)|
    ((_net_0)?_add_map_x_69_data_out_index:10'b0);
   assign  data_out_index180 = ((_net_1)?_add_map_x_69_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_69_data_near:10'b0);
   assign  data_out_index181 = ((_net_1)?_add_map_x_70_data_near:10'b0)|
    ((_net_0)?_add_map_x_70_data_out_index:10'b0);
   assign  data_out_index182 = ((_net_1)?_add_map_x_70_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_70_data_near:10'b0);
   assign  data_out_index183 = ((_net_1)?_add_map_x_71_data_near:10'b0)|
    ((_net_0)?_add_map_x_71_data_out_index:10'b0);
   assign  data_out_index184 = ((_net_1)?_add_map_x_71_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_71_data_near:10'b0);
   assign  data_out_index185 = ((_net_1)?_add_map_x_72_data_near:10'b0)|
    ((_net_0)?_add_map_x_72_data_out_index:10'b0);
   assign  data_out_index186 = ((_net_1)?_add_map_x_72_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_72_data_near:10'b0);
   assign  data_out_index187 = ((_net_1)?_add_map_x_73_data_near:10'b0)|
    ((_net_0)?_add_map_x_73_data_out_index:10'b0);
   assign  data_out_index188 = ((_net_1)?_add_map_x_73_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_73_data_near:10'b0);
   assign  data_out_index189 = ((_net_1)?_add_map_x_74_data_near:10'b0)|
    ((_net_0)?_add_map_x_74_data_out_index:10'b0);
   assign  data_out_index190 = ((_net_1)?_add_map_x_74_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_74_data_near:10'b0);
   assign  data_out_index193 = ((_net_1)?_add_map_x_75_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_75_data_near:10'b0);
   assign  data_out_index194 = ((_net_1)?_add_map_x_75_data_near:10'b0)|
    ((_net_0)?_add_map_x_75_data_out_index:10'b0);
   assign  data_out_index195 = ((_net_1)?_add_map_x_76_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_76_data_near:10'b0);
   assign  data_out_index196 = ((_net_1)?_add_map_x_76_data_near:10'b0)|
    ((_net_0)?_add_map_x_76_data_out_index:10'b0);
   assign  data_out_index197 = ((_net_1)?_add_map_x_77_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_77_data_near:10'b0);
   assign  data_out_index198 = ((_net_1)?_add_map_x_77_data_near:10'b0)|
    ((_net_0)?_add_map_x_77_data_out_index:10'b0);
   assign  data_out_index199 = ((_net_1)?_add_map_x_78_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_78_data_near:10'b0);
   assign  data_out_index200 = ((_net_1)?_add_map_x_78_data_near:10'b0)|
    ((_net_0)?_add_map_x_78_data_out_index:10'b0);
   assign  data_out_index201 = ((_net_1)?_add_map_x_79_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_79_data_near:10'b0);
   assign  data_out_index202 = ((_net_1)?_add_map_x_79_data_near:10'b0)|
    ((_net_0)?_add_map_x_79_data_out_index:10'b0);
   assign  data_out_index203 = ((_net_1)?_add_map_x_80_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_80_data_near:10'b0);
   assign  data_out_index204 = ((_net_1)?_add_map_x_80_data_near:10'b0)|
    ((_net_0)?_add_map_x_80_data_out_index:10'b0);
   assign  data_out_index205 = ((_net_1)?_add_map_x_81_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_81_data_near:10'b0);
   assign  data_out_index206 = ((_net_1)?_add_map_x_81_data_near:10'b0)|
    ((_net_0)?_add_map_x_81_data_out_index:10'b0);
   assign  data_out_index207 = ((_net_1)?_add_map_x_82_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_82_data_near:10'b0);
   assign  data_out_index208 = ((_net_1)?_add_map_x_82_data_near:10'b0)|
    ((_net_0)?_add_map_x_82_data_out_index:10'b0);
   assign  data_out_index209 = ((_net_1)?_add_map_x_83_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_83_data_near:10'b0);
   assign  data_out_index210 = ((_net_1)?_add_map_x_83_data_near:10'b0)|
    ((_net_0)?_add_map_x_83_data_out_index:10'b0);
   assign  data_out_index211 = ((_net_1)?_add_map_x_84_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_84_data_near:10'b0);
   assign  data_out_index212 = ((_net_1)?_add_map_x_84_data_near:10'b0)|
    ((_net_0)?_add_map_x_84_data_out_index:10'b0);
   assign  data_out_index213 = ((_net_1)?_add_map_x_85_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_85_data_near:10'b0);
   assign  data_out_index214 = ((_net_1)?_add_map_x_85_data_near:10'b0)|
    ((_net_0)?_add_map_x_85_data_out_index:10'b0);
   assign  data_out_index215 = ((_net_1)?_add_map_x_86_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_86_data_near:10'b0);
   assign  data_out_index216 = ((_net_1)?_add_map_x_86_data_near:10'b0)|
    ((_net_0)?_add_map_x_86_data_out_index:10'b0);
   assign  data_out_index217 = ((_net_1)?_add_map_x_87_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_87_data_near:10'b0);
   assign  data_out_index218 = ((_net_1)?_add_map_x_87_data_near:10'b0)|
    ((_net_0)?_add_map_x_87_data_out_index:10'b0);
   assign  data_out_index219 = ((_net_1)?_add_map_x_88_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_88_data_near:10'b0);
   assign  data_out_index220 = ((_net_1)?_add_map_x_88_data_near:10'b0)|
    ((_net_0)?_add_map_x_88_data_out_index:10'b0);
   assign  data_out_index221 = ((_net_1)?_add_map_x_89_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_89_data_near:10'b0);
   assign  data_out_index222 = ((_net_1)?_add_map_x_89_data_near:10'b0)|
    ((_net_0)?_add_map_x_89_data_out_index:10'b0);
   assign  data_out_index225 = ((_net_1)?_add_map_x_90_data_near:10'b0)|
    ((_net_0)?_add_map_x_90_data_out_index:10'b0);
   assign  data_out_index226 = ((_net_1)?_add_map_x_90_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_90_data_near:10'b0);
   assign  data_out_index227 = ((_net_1)?_add_map_x_91_data_near:10'b0)|
    ((_net_0)?_add_map_x_91_data_out_index:10'b0);
   assign  data_out_index228 = ((_net_1)?_add_map_x_91_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_91_data_near:10'b0);
   assign  data_out_index229 = ((_net_1)?_add_map_x_92_data_near:10'b0)|
    ((_net_0)?_add_map_x_92_data_out_index:10'b0);
   assign  data_out_index230 = ((_net_1)?_add_map_x_92_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_92_data_near:10'b0);
   assign  data_out_index231 = ((_net_1)?_add_map_x_93_data_near:10'b0)|
    ((_net_0)?_add_map_x_93_data_out_index:10'b0);
   assign  data_out_index232 = ((_net_1)?_add_map_x_93_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_93_data_near:10'b0);
   assign  data_out_index233 = ((_net_1)?_add_map_x_94_data_near:10'b0)|
    ((_net_0)?_add_map_x_94_data_out_index:10'b0);
   assign  data_out_index234 = ((_net_1)?_add_map_x_94_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_94_data_near:10'b0);
   assign  data_out_index235 = ((_net_1)?_add_map_x_95_data_near:10'b0)|
    ((_net_0)?_add_map_x_95_data_out_index:10'b0);
   assign  data_out_index236 = ((_net_1)?_add_map_x_95_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_95_data_near:10'b0);
   assign  data_out_index237 = ((_net_1)?_add_map_x_96_data_near:10'b0)|
    ((_net_0)?_add_map_x_96_data_out_index:10'b0);
   assign  data_out_index238 = ((_net_1)?_add_map_x_96_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_96_data_near:10'b0);
   assign  data_out_index239 = ((_net_1)?_add_map_x_97_data_near:10'b0)|
    ((_net_0)?_add_map_x_97_data_out_index:10'b0);
   assign  data_out_index240 = ((_net_1)?_add_map_x_97_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_97_data_near:10'b0);
   assign  data_out_index241 = ((_net_1)?_add_map_x_98_data_near:10'b0)|
    ((_net_0)?_add_map_x_98_data_out_index:10'b0);
   assign  data_out_index242 = ((_net_1)?_add_map_x_98_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_98_data_near:10'b0);
   assign  data_out_index243 = ((_net_1)?_add_map_x_99_data_near:10'b0)|
    ((_net_0)?_add_map_x_99_data_out_index:10'b0);
   assign  data_out_index244 = ((_net_1)?_add_map_x_99_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_99_data_near:10'b0);
   assign  data_out_index245 = ((_net_1)?_add_map_x_100_data_near:10'b0)|
    ((_net_0)?_add_map_x_100_data_out_index:10'b0);
   assign  data_out_index246 = ((_net_1)?_add_map_x_100_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_100_data_near:10'b0);
   assign  data_out_index247 = ((_net_1)?_add_map_x_101_data_near:10'b0)|
    ((_net_0)?_add_map_x_101_data_out_index:10'b0);
   assign  data_out_index248 = ((_net_1)?_add_map_x_101_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_101_data_near:10'b0);
   assign  data_out_index249 = ((_net_1)?_add_map_x_102_data_near:10'b0)|
    ((_net_0)?_add_map_x_102_data_out_index:10'b0);
   assign  data_out_index250 = ((_net_1)?_add_map_x_102_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_102_data_near:10'b0);
   assign  data_out_index251 = ((_net_1)?_add_map_x_103_data_near:10'b0)|
    ((_net_0)?_add_map_x_103_data_out_index:10'b0);
   assign  data_out_index252 = ((_net_1)?_add_map_x_103_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_103_data_near:10'b0);
   assign  data_out_index253 = ((_net_1)?_add_map_x_104_data_near:10'b0)|
    ((_net_0)?_add_map_x_104_data_out_index:10'b0);
   assign  data_out_index254 = ((_net_1)?_add_map_x_104_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_104_data_near:10'b0);
   assign  data_out_index257 = ((_net_1)?_add_map_x_105_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_105_data_near:10'b0);
   assign  data_out_index258 = ((_net_1)?_add_map_x_105_data_near:10'b0)|
    ((_net_0)?_add_map_x_105_data_out_index:10'b0);
   assign  data_out_index259 = ((_net_1)?_add_map_x_106_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_106_data_near:10'b0);
   assign  data_out_index260 = ((_net_1)?_add_map_x_106_data_near:10'b0)|
    ((_net_0)?_add_map_x_106_data_out_index:10'b0);
   assign  data_out_index261 = ((_net_1)?_add_map_x_107_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_107_data_near:10'b0);
   assign  data_out_index262 = ((_net_1)?_add_map_x_107_data_near:10'b0)|
    ((_net_0)?_add_map_x_107_data_out_index:10'b0);
   assign  data_out_index263 = ((_net_1)?_add_map_x_108_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_108_data_near:10'b0);
   assign  data_out_index264 = ((_net_1)?_add_map_x_108_data_near:10'b0)|
    ((_net_0)?_add_map_x_108_data_out_index:10'b0);
   assign  data_out_index265 = ((_net_1)?_add_map_x_109_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_109_data_near:10'b0);
   assign  data_out_index266 = ((_net_1)?_add_map_x_109_data_near:10'b0)|
    ((_net_0)?_add_map_x_109_data_out_index:10'b0);
   assign  data_out_index267 = ((_net_1)?_add_map_x_110_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_110_data_near:10'b0);
   assign  data_out_index268 = ((_net_1)?_add_map_x_110_data_near:10'b0)|
    ((_net_0)?_add_map_x_110_data_out_index:10'b0);
   assign  data_out_index269 = ((_net_1)?_add_map_x_111_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_111_data_near:10'b0);
   assign  data_out_index270 = ((_net_1)?_add_map_x_111_data_near:10'b0)|
    ((_net_0)?_add_map_x_111_data_out_index:10'b0);
   assign  data_out_index271 = ((_net_1)?_add_map_x_112_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_112_data_near:10'b0);
   assign  data_out_index272 = ((_net_1)?_add_map_x_112_data_near:10'b0)|
    ((_net_0)?_add_map_x_112_data_out_index:10'b0);
   assign  data_out_index273 = ((_net_1)?_add_map_x_113_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_113_data_near:10'b0);
   assign  data_out_index274 = ((_net_1)?_add_map_x_113_data_near:10'b0)|
    ((_net_0)?_add_map_x_113_data_out_index:10'b0);
   assign  data_out_index275 = ((_net_1)?_add_map_x_114_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_114_data_near:10'b0);
   assign  data_out_index276 = ((_net_1)?_add_map_x_114_data_near:10'b0)|
    ((_net_0)?_add_map_x_114_data_out_index:10'b0);
   assign  data_out_index277 = ((_net_1)?_add_map_x_115_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_115_data_near:10'b0);
   assign  data_out_index278 = ((_net_1)?_add_map_x_115_data_near:10'b0)|
    ((_net_0)?_add_map_x_115_data_out_index:10'b0);
   assign  data_out_index279 = ((_net_1)?_add_map_x_116_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_116_data_near:10'b0);
   assign  data_out_index280 = ((_net_1)?_add_map_x_116_data_near:10'b0)|
    ((_net_0)?_add_map_x_116_data_out_index:10'b0);
   assign  data_out_index281 = ((_net_1)?_add_map_x_117_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_117_data_near:10'b0);
   assign  data_out_index282 = ((_net_1)?_add_map_x_117_data_near:10'b0)|
    ((_net_0)?_add_map_x_117_data_out_index:10'b0);
   assign  data_out_index283 = ((_net_1)?_add_map_x_118_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_118_data_near:10'b0);
   assign  data_out_index284 = ((_net_1)?_add_map_x_118_data_near:10'b0)|
    ((_net_0)?_add_map_x_118_data_out_index:10'b0);
   assign  data_out_index285 = ((_net_1)?_add_map_x_119_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_119_data_near:10'b0);
   assign  data_out_index286 = ((_net_1)?_add_map_x_119_data_near:10'b0)|
    ((_net_0)?_add_map_x_119_data_out_index:10'b0);
   assign  data_out_index289 = ((_net_1)?_add_map_x_120_data_near:10'b0)|
    ((_net_0)?_add_map_x_120_data_out_index:10'b0);
   assign  data_out_index290 = ((_net_1)?_add_map_x_120_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_120_data_near:10'b0);
   assign  data_out_index291 = ((_net_1)?_add_map_x_121_data_near:10'b0)|
    ((_net_0)?_add_map_x_121_data_out_index:10'b0);
   assign  data_out_index292 = ((_net_1)?_add_map_x_121_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_121_data_near:10'b0);
   assign  data_out_index293 = ((_net_1)?_add_map_x_122_data_near:10'b0)|
    ((_net_0)?_add_map_x_122_data_out_index:10'b0);
   assign  data_out_index294 = ((_net_1)?_add_map_x_122_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_122_data_near:10'b0);
   assign  data_out_index295 = ((_net_1)?_add_map_x_123_data_near:10'b0)|
    ((_net_0)?_add_map_x_123_data_out_index:10'b0);
   assign  data_out_index296 = ((_net_1)?_add_map_x_123_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_123_data_near:10'b0);
   assign  data_out_index297 = ((_net_1)?_add_map_x_124_data_near:10'b0)|
    ((_net_0)?_add_map_x_124_data_out_index:10'b0);
   assign  data_out_index298 = ((_net_1)?_add_map_x_124_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_124_data_near:10'b0);
   assign  data_out_index299 = ((_net_1)?_add_map_x_125_data_near:10'b0)|
    ((_net_0)?_add_map_x_125_data_out_index:10'b0);
   assign  data_out_index300 = ((_net_1)?_add_map_x_125_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_125_data_near:10'b0);
   assign  data_out_index301 = ((_net_1)?_add_map_x_126_data_near:10'b0)|
    ((_net_0)?_add_map_x_126_data_out_index:10'b0);
   assign  data_out_index302 = ((_net_1)?_add_map_x_126_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_126_data_near:10'b0);
   assign  data_out_index303 = ((_net_1)?_add_map_x_127_data_near:10'b0)|
    ((_net_0)?_add_map_x_127_data_out_index:10'b0);
   assign  data_out_index304 = ((_net_1)?_add_map_x_127_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_127_data_near:10'b0);
   assign  data_out_index305 = ((_net_1)?_add_map_x_128_data_near:10'b0)|
    ((_net_0)?_add_map_x_128_data_out_index:10'b0);
   assign  data_out_index306 = ((_net_1)?_add_map_x_128_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_128_data_near:10'b0);
   assign  data_out_index307 = ((_net_1)?_add_map_x_129_data_near:10'b0)|
    ((_net_0)?_add_map_x_129_data_out_index:10'b0);
   assign  data_out_index308 = ((_net_1)?_add_map_x_129_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_129_data_near:10'b0);
   assign  data_out_index309 = ((_net_1)?_add_map_x_130_data_near:10'b0)|
    ((_net_0)?_add_map_x_130_data_out_index:10'b0);
   assign  data_out_index310 = ((_net_1)?_add_map_x_130_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_130_data_near:10'b0);
   assign  data_out_index311 = ((_net_1)?_add_map_x_131_data_near:10'b0)|
    ((_net_0)?_add_map_x_131_data_out_index:10'b0);
   assign  data_out_index312 = ((_net_1)?_add_map_x_131_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_131_data_near:10'b0);
   assign  data_out_index313 = ((_net_1)?_add_map_x_132_data_near:10'b0)|
    ((_net_0)?_add_map_x_132_data_out_index:10'b0);
   assign  data_out_index314 = ((_net_1)?_add_map_x_132_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_132_data_near:10'b0);
   assign  data_out_index315 = ((_net_1)?_add_map_x_133_data_near:10'b0)|
    ((_net_0)?_add_map_x_133_data_out_index:10'b0);
   assign  data_out_index316 = ((_net_1)?_add_map_x_133_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_133_data_near:10'b0);
   assign  data_out_index317 = ((_net_1)?_add_map_x_134_data_near:10'b0)|
    ((_net_0)?_add_map_x_134_data_out_index:10'b0);
   assign  data_out_index318 = ((_net_1)?_add_map_x_134_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_134_data_near:10'b0);
   assign  data_out_index321 = ((_net_1)?_add_map_x_135_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_135_data_near:10'b0);
   assign  data_out_index322 = ((_net_1)?_add_map_x_135_data_near:10'b0)|
    ((_net_0)?_add_map_x_135_data_out_index:10'b0);
   assign  data_out_index323 = ((_net_1)?_add_map_x_136_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_136_data_near:10'b0);
   assign  data_out_index324 = ((_net_1)?_add_map_x_136_data_near:10'b0)|
    ((_net_0)?_add_map_x_136_data_out_index:10'b0);
   assign  data_out_index325 = ((_net_1)?_add_map_x_137_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_137_data_near:10'b0);
   assign  data_out_index326 = ((_net_1)?_add_map_x_137_data_near:10'b0)|
    ((_net_0)?_add_map_x_137_data_out_index:10'b0);
   assign  data_out_index327 = ((_net_1)?_add_map_x_138_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_138_data_near:10'b0);
   assign  data_out_index328 = ((_net_1)?_add_map_x_138_data_near:10'b0)|
    ((_net_0)?_add_map_x_138_data_out_index:10'b0);
   assign  data_out_index329 = ((_net_1)?_add_map_x_139_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_139_data_near:10'b0);
   assign  data_out_index330 = ((_net_1)?_add_map_x_139_data_near:10'b0)|
    ((_net_0)?_add_map_x_139_data_out_index:10'b0);
   assign  data_out_index331 = ((_net_1)?_add_map_x_140_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_140_data_near:10'b0);
   assign  data_out_index332 = ((_net_1)?_add_map_x_140_data_near:10'b0)|
    ((_net_0)?_add_map_x_140_data_out_index:10'b0);
   assign  data_out_index333 = ((_net_1)?_add_map_x_141_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_141_data_near:10'b0);
   assign  data_out_index334 = ((_net_1)?_add_map_x_141_data_near:10'b0)|
    ((_net_0)?_add_map_x_141_data_out_index:10'b0);
   assign  data_out_index335 = ((_net_1)?_add_map_x_142_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_142_data_near:10'b0);
   assign  data_out_index336 = ((_net_1)?_add_map_x_142_data_near:10'b0)|
    ((_net_0)?_add_map_x_142_data_out_index:10'b0);
   assign  data_out_index337 = ((_net_1)?_add_map_x_143_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_143_data_near:10'b0);
   assign  data_out_index338 = ((_net_1)?_add_map_x_143_data_near:10'b0)|
    ((_net_0)?_add_map_x_143_data_out_index:10'b0);
   assign  data_out_index339 = ((_net_1)?_add_map_x_144_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_144_data_near:10'b0);
   assign  data_out_index340 = ((_net_1)?_add_map_x_144_data_near:10'b0)|
    ((_net_0)?_add_map_x_144_data_out_index:10'b0);
   assign  data_out_index341 = ((_net_1)?_add_map_x_145_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_145_data_near:10'b0);
   assign  data_out_index342 = ((_net_1)?_add_map_x_145_data_near:10'b0)|
    ((_net_0)?_add_map_x_145_data_out_index:10'b0);
   assign  data_out_index343 = ((_net_1)?_add_map_x_146_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_146_data_near:10'b0);
   assign  data_out_index344 = ((_net_1)?_add_map_x_146_data_near:10'b0)|
    ((_net_0)?_add_map_x_146_data_out_index:10'b0);
   assign  data_out_index345 = ((_net_1)?_add_map_x_147_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_147_data_near:10'b0);
   assign  data_out_index346 = ((_net_1)?_add_map_x_147_data_near:10'b0)|
    ((_net_0)?_add_map_x_147_data_out_index:10'b0);
   assign  data_out_index347 = ((_net_1)?_add_map_x_148_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_148_data_near:10'b0);
   assign  data_out_index348 = ((_net_1)?_add_map_x_148_data_near:10'b0)|
    ((_net_0)?_add_map_x_148_data_out_index:10'b0);
   assign  data_out_index349 = ((_net_1)?_add_map_x_149_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_149_data_near:10'b0);
   assign  data_out_index350 = ((_net_1)?_add_map_x_149_data_near:10'b0)|
    ((_net_0)?_add_map_x_149_data_out_index:10'b0);
   assign  data_out_index353 = ((_net_1)?_add_map_x_150_data_near:10'b0)|
    ((_net_0)?_add_map_x_150_data_out_index:10'b0);
   assign  data_out_index354 = ((_net_1)?_add_map_x_150_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_150_data_near:10'b0);
   assign  data_out_index355 = ((_net_1)?_add_map_x_151_data_near:10'b0)|
    ((_net_0)?_add_map_x_151_data_out_index:10'b0);
   assign  data_out_index356 = ((_net_1)?_add_map_x_151_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_151_data_near:10'b0);
   assign  data_out_index357 = ((_net_1)?_add_map_x_152_data_near:10'b0)|
    ((_net_0)?_add_map_x_152_data_out_index:10'b0);
   assign  data_out_index358 = ((_net_1)?_add_map_x_152_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_152_data_near:10'b0);
   assign  data_out_index359 = ((_net_1)?_add_map_x_153_data_near:10'b0)|
    ((_net_0)?_add_map_x_153_data_out_index:10'b0);
   assign  data_out_index360 = ((_net_1)?_add_map_x_153_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_153_data_near:10'b0);
   assign  data_out_index361 = ((_net_1)?_add_map_x_154_data_near:10'b0)|
    ((_net_0)?_add_map_x_154_data_out_index:10'b0);
   assign  data_out_index362 = ((_net_1)?_add_map_x_154_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_154_data_near:10'b0);
   assign  data_out_index363 = ((_net_1)?_add_map_x_155_data_near:10'b0)|
    ((_net_0)?_add_map_x_155_data_out_index:10'b0);
   assign  data_out_index364 = ((_net_1)?_add_map_x_155_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_155_data_near:10'b0);
   assign  data_out_index365 = ((_net_1)?_add_map_x_156_data_near:10'b0)|
    ((_net_0)?_add_map_x_156_data_out_index:10'b0);
   assign  data_out_index366 = ((_net_1)?_add_map_x_156_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_156_data_near:10'b0);
   assign  data_out_index367 = ((_net_1)?_add_map_x_157_data_near:10'b0)|
    ((_net_0)?_add_map_x_157_data_out_index:10'b0);
   assign  data_out_index368 = ((_net_1)?_add_map_x_157_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_157_data_near:10'b0);
   assign  data_out_index369 = ((_net_1)?_add_map_x_158_data_near:10'b0)|
    ((_net_0)?_add_map_x_158_data_out_index:10'b0);
   assign  data_out_index370 = ((_net_1)?_add_map_x_158_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_158_data_near:10'b0);
   assign  data_out_index371 = ((_net_1)?_add_map_x_159_data_near:10'b0)|
    ((_net_0)?_add_map_x_159_data_out_index:10'b0);
   assign  data_out_index372 = ((_net_1)?_add_map_x_159_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_159_data_near:10'b0);
   assign  data_out_index373 = ((_net_1)?_add_map_x_160_data_near:10'b0)|
    ((_net_0)?_add_map_x_160_data_out_index:10'b0);
   assign  data_out_index374 = ((_net_1)?_add_map_x_160_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_160_data_near:10'b0);
   assign  data_out_index375 = ((_net_1)?_add_map_x_161_data_near:10'b0)|
    ((_net_0)?_add_map_x_161_data_out_index:10'b0);
   assign  data_out_index376 = ((_net_1)?_add_map_x_161_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_161_data_near:10'b0);
   assign  data_out_index377 = ((_net_1)?_add_map_x_162_data_near:10'b0)|
    ((_net_0)?_add_map_x_162_data_out_index:10'b0);
   assign  data_out_index378 = ((_net_1)?_add_map_x_162_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_162_data_near:10'b0);
   assign  data_out_index379 = ((_net_1)?_add_map_x_163_data_near:10'b0)|
    ((_net_0)?_add_map_x_163_data_out_index:10'b0);
   assign  data_out_index380 = ((_net_1)?_add_map_x_163_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_163_data_near:10'b0);
   assign  data_out_index381 = ((_net_1)?_add_map_x_164_data_near:10'b0)|
    ((_net_0)?_add_map_x_164_data_out_index:10'b0);
   assign  data_out_index382 = ((_net_1)?_add_map_x_164_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_164_data_near:10'b0);
   assign  data_out_index385 = ((_net_1)?_add_map_x_165_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_165_data_near:10'b0);
   assign  data_out_index386 = ((_net_1)?_add_map_x_165_data_near:10'b0)|
    ((_net_0)?_add_map_x_165_data_out_index:10'b0);
   assign  data_out_index387 = ((_net_1)?_add_map_x_166_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_166_data_near:10'b0);
   assign  data_out_index388 = ((_net_1)?_add_map_x_166_data_near:10'b0)|
    ((_net_0)?_add_map_x_166_data_out_index:10'b0);
   assign  data_out_index389 = ((_net_1)?_add_map_x_167_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_167_data_near:10'b0);
   assign  data_out_index390 = ((_net_1)?_add_map_x_167_data_near:10'b0)|
    ((_net_0)?_add_map_x_167_data_out_index:10'b0);
   assign  data_out_index391 = ((_net_1)?_add_map_x_168_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_168_data_near:10'b0);
   assign  data_out_index392 = ((_net_1)?_add_map_x_168_data_near:10'b0)|
    ((_net_0)?_add_map_x_168_data_out_index:10'b0);
   assign  data_out_index393 = ((_net_1)?_add_map_x_169_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_169_data_near:10'b0);
   assign  data_out_index394 = ((_net_1)?_add_map_x_169_data_near:10'b0)|
    ((_net_0)?_add_map_x_169_data_out_index:10'b0);
   assign  data_out_index395 = ((_net_1)?_add_map_x_170_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_170_data_near:10'b0);
   assign  data_out_index396 = ((_net_1)?_add_map_x_170_data_near:10'b0)|
    ((_net_0)?_add_map_x_170_data_out_index:10'b0);
   assign  data_out_index397 = ((_net_1)?_add_map_x_171_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_171_data_near:10'b0);
   assign  data_out_index398 = ((_net_1)?_add_map_x_171_data_near:10'b0)|
    ((_net_0)?_add_map_x_171_data_out_index:10'b0);
   assign  data_out_index399 = ((_net_1)?_add_map_x_172_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_172_data_near:10'b0);
   assign  data_out_index400 = ((_net_1)?_add_map_x_172_data_near:10'b0)|
    ((_net_0)?_add_map_x_172_data_out_index:10'b0);
   assign  data_out_index401 = ((_net_1)?_add_map_x_173_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_173_data_near:10'b0);
   assign  data_out_index402 = ((_net_1)?_add_map_x_173_data_near:10'b0)|
    ((_net_0)?_add_map_x_173_data_out_index:10'b0);
   assign  data_out_index403 = ((_net_1)?_add_map_x_174_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_174_data_near:10'b0);
   assign  data_out_index404 = ((_net_1)?_add_map_x_174_data_near:10'b0)|
    ((_net_0)?_add_map_x_174_data_out_index:10'b0);
   assign  data_out_index405 = ((_net_1)?_add_map_x_175_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_175_data_near:10'b0);
   assign  data_out_index406 = ((_net_1)?_add_map_x_175_data_near:10'b0)|
    ((_net_0)?_add_map_x_175_data_out_index:10'b0);
   assign  data_out_index407 = ((_net_1)?_add_map_x_176_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_176_data_near:10'b0);
   assign  data_out_index408 = ((_net_1)?_add_map_x_176_data_near:10'b0)|
    ((_net_0)?_add_map_x_176_data_out_index:10'b0);
   assign  data_out_index409 = ((_net_1)?_add_map_x_177_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_177_data_near:10'b0);
   assign  data_out_index410 = ((_net_1)?_add_map_x_177_data_near:10'b0)|
    ((_net_0)?_add_map_x_177_data_out_index:10'b0);
   assign  data_out_index411 = ((_net_1)?_add_map_x_178_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_178_data_near:10'b0);
   assign  data_out_index412 = ((_net_1)?_add_map_x_178_data_near:10'b0)|
    ((_net_0)?_add_map_x_178_data_out_index:10'b0);
   assign  data_out_index413 = ((_net_1)?_add_map_x_179_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_179_data_near:10'b0);
   assign  data_out_index414 = ((_net_1)?_add_map_x_179_data_near:10'b0)|
    ((_net_0)?_add_map_x_179_data_out_index:10'b0);
   assign  data_out_index417 = ((_net_1)?_add_map_x_180_data_near:10'b0)|
    ((_net_0)?_add_map_x_180_data_out_index:10'b0);
   assign  data_out_index418 = ((_net_1)?_add_map_x_180_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_180_data_near:10'b0);
   assign  data_out_index419 = ((_net_1)?_add_map_x_181_data_near:10'b0)|
    ((_net_0)?_add_map_x_181_data_out_index:10'b0);
   assign  data_out_index420 = ((_net_1)?_add_map_x_181_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_181_data_near:10'b0);
   assign  data_out_index421 = ((_net_1)?_add_map_x_182_data_near:10'b0)|
    ((_net_0)?_add_map_x_182_data_out_index:10'b0);
   assign  data_out_index422 = ((_net_1)?_add_map_x_182_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_182_data_near:10'b0);
   assign  data_out_index423 = ((_net_1)?_add_map_x_183_data_near:10'b0)|
    ((_net_0)?_add_map_x_183_data_out_index:10'b0);
   assign  data_out_index424 = ((_net_1)?_add_map_x_183_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_183_data_near:10'b0);
   assign  data_out_index425 = ((_net_1)?_add_map_x_184_data_near:10'b0)|
    ((_net_0)?_add_map_x_184_data_out_index:10'b0);
   assign  data_out_index426 = ((_net_1)?_add_map_x_184_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_184_data_near:10'b0);
   assign  data_out_index427 = ((_net_1)?_add_map_x_185_data_near:10'b0)|
    ((_net_0)?_add_map_x_185_data_out_index:10'b0);
   assign  data_out_index428 = ((_net_1)?_add_map_x_185_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_185_data_near:10'b0);
   assign  data_out_index429 = ((_net_1)?_add_map_x_186_data_near:10'b0)|
    ((_net_0)?_add_map_x_186_data_out_index:10'b0);
   assign  data_out_index430 = ((_net_1)?_add_map_x_186_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_186_data_near:10'b0);
   assign  data_out_index431 = ((_net_1)?_add_map_x_187_data_near:10'b0)|
    ((_net_0)?_add_map_x_187_data_out_index:10'b0);
   assign  data_out_index432 = ((_net_1)?_add_map_x_187_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_187_data_near:10'b0);
   assign  data_out_index433 = ((_net_1)?_add_map_x_188_data_near:10'b0)|
    ((_net_0)?_add_map_x_188_data_out_index:10'b0);
   assign  data_out_index434 = ((_net_1)?_add_map_x_188_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_188_data_near:10'b0);
   assign  data_out_index435 = ((_net_1)?_add_map_x_189_data_near:10'b0)|
    ((_net_0)?_add_map_x_189_data_out_index:10'b0);
   assign  data_out_index436 = ((_net_1)?_add_map_x_189_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_189_data_near:10'b0);
   assign  data_out_index437 = ((_net_1)?_add_map_x_190_data_near:10'b0)|
    ((_net_0)?_add_map_x_190_data_out_index:10'b0);
   assign  data_out_index438 = ((_net_1)?_add_map_x_190_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_190_data_near:10'b0);
   assign  data_out_index439 = ((_net_1)?_add_map_x_191_data_near:10'b0)|
    ((_net_0)?_add_map_x_191_data_out_index:10'b0);
   assign  data_out_index440 = ((_net_1)?_add_map_x_191_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_191_data_near:10'b0);
   assign  data_out_index441 = ((_net_1)?_add_map_x_192_data_near:10'b0)|
    ((_net_0)?_add_map_x_192_data_out_index:10'b0);
   assign  data_out_index442 = ((_net_1)?_add_map_x_192_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_192_data_near:10'b0);
   assign  data_out_index443 = ((_net_1)?_add_map_x_193_data_near:10'b0)|
    ((_net_0)?_add_map_x_193_data_out_index:10'b0);
   assign  data_out_index444 = ((_net_1)?_add_map_x_193_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_193_data_near:10'b0);
   assign  data_out_index445 = ((_net_1)?_add_map_x_194_data_near:10'b0)|
    ((_net_0)?_add_map_x_194_data_out_index:10'b0);
   assign  data_out_index446 = ((_net_1)?_add_map_x_194_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_194_data_near:10'b0);
   assign  data_out_index449 = ((_net_1)?_add_map_x_195_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_195_data_near:10'b0);
   assign  data_out_index450 = ((_net_1)?_add_map_x_195_data_near:10'b0)|
    ((_net_0)?_add_map_x_195_data_out_index:10'b0);
   assign  data_out_index451 = ((_net_1)?_add_map_x_196_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_196_data_near:10'b0);
   assign  data_out_index452 = ((_net_1)?_add_map_x_196_data_near:10'b0)|
    ((_net_0)?_add_map_x_196_data_out_index:10'b0);
   assign  data_out_index453 = ((_net_1)?_add_map_x_197_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_197_data_near:10'b0);
   assign  data_out_index454 = ((_net_1)?_add_map_x_197_data_near:10'b0)|
    ((_net_0)?_add_map_x_197_data_out_index:10'b0);
   assign  data_out_index455 = ((_net_1)?_add_map_x_198_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_198_data_near:10'b0);
   assign  data_out_index456 = ((_net_1)?_add_map_x_198_data_near:10'b0)|
    ((_net_0)?_add_map_x_198_data_out_index:10'b0);
   assign  data_out_index457 = ((_net_1)?_add_map_x_199_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_199_data_near:10'b0);
   assign  data_out_index458 = ((_net_1)?_add_map_x_199_data_near:10'b0)|
    ((_net_0)?_add_map_x_199_data_out_index:10'b0);
   assign  data_out_index459 = ((_net_1)?_add_map_x_200_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_200_data_near:10'b0);
   assign  data_out_index460 = ((_net_1)?_add_map_x_200_data_near:10'b0)|
    ((_net_0)?_add_map_x_200_data_out_index:10'b0);
   assign  data_out_index461 = ((_net_1)?_add_map_x_201_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_201_data_near:10'b0);
   assign  data_out_index462 = ((_net_1)?_add_map_x_201_data_near:10'b0)|
    ((_net_0)?_add_map_x_201_data_out_index:10'b0);
   assign  data_out_index463 = ((_net_1)?_add_map_x_202_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_202_data_near:10'b0);
   assign  data_out_index464 = ((_net_1)?_add_map_x_202_data_near:10'b0)|
    ((_net_0)?_add_map_x_202_data_out_index:10'b0);
   assign  data_out_index465 = ((_net_1)?_add_map_x_203_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_203_data_near:10'b0);
   assign  data_out_index466 = ((_net_1)?_add_map_x_203_data_near:10'b0)|
    ((_net_0)?_add_map_x_203_data_out_index:10'b0);
   assign  data_out_index467 = ((_net_1)?_add_map_x_204_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_204_data_near:10'b0);
   assign  data_out_index468 = ((_net_1)?_add_map_x_204_data_near:10'b0)|
    ((_net_0)?_add_map_x_204_data_out_index:10'b0);
   assign  data_out_index469 = ((_net_1)?_add_map_x_205_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_205_data_near:10'b0);
   assign  data_out_index470 = ((_net_1)?_add_map_x_205_data_near:10'b0)|
    ((_net_0)?_add_map_x_205_data_out_index:10'b0);
   assign  data_out_index471 = ((_net_1)?_add_map_x_206_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_206_data_near:10'b0);
   assign  data_out_index472 = ((_net_1)?_add_map_x_206_data_near:10'b0)|
    ((_net_0)?_add_map_x_206_data_out_index:10'b0);
   assign  data_out_index473 = ((_net_1)?_add_map_x_207_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_207_data_near:10'b0);
   assign  data_out_index474 = ((_net_1)?_add_map_x_207_data_near:10'b0)|
    ((_net_0)?_add_map_x_207_data_out_index:10'b0);
   assign  data_out_index475 = ((_net_1)?_add_map_x_208_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_208_data_near:10'b0);
   assign  data_out_index476 = ((_net_1)?_add_map_x_208_data_near:10'b0)|
    ((_net_0)?_add_map_x_208_data_out_index:10'b0);
   assign  data_out_index477 = ((_net_1)?_add_map_x_209_data_out_index:10'b0)|
    ((_net_0)?_add_map_x_209_data_near:10'b0);
   assign  data_out_index478 = ((_net_1)?_add_map_x_209_data_near:10'b0)|
    ((_net_0)?_add_map_x_209_data_out_index:10'b0);
   assign  sg_out33 = ((_net_1)?_add_map_x_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_s_g:2'b0);
   assign  sg_out34 = ((_net_1)?_add_map_x_s_g:2'b0)|
    ((_net_0)?_add_map_x_s_g_near:2'b0);
   assign  sg_out35 = ((_net_1)?_add_map_x_1_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_1_s_g:2'b0);
   assign  sg_out36 = ((_net_1)?_add_map_x_1_s_g:2'b0)|
    ((_net_0)?_add_map_x_1_s_g_near:2'b0);
   assign  sg_out37 = ((_net_1)?_add_map_x_2_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_2_s_g:2'b0);
   assign  sg_out38 = ((_net_1)?_add_map_x_2_s_g:2'b0)|
    ((_net_0)?_add_map_x_2_s_g_near:2'b0);
   assign  sg_out39 = ((_net_1)?_add_map_x_3_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_3_s_g:2'b0);
   assign  sg_out40 = ((_net_1)?_add_map_x_3_s_g:2'b0)|
    ((_net_0)?_add_map_x_3_s_g_near:2'b0);
   assign  sg_out41 = ((_net_1)?_add_map_x_4_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_4_s_g:2'b0);
   assign  sg_out42 = ((_net_1)?_add_map_x_4_s_g:2'b0)|
    ((_net_0)?_add_map_x_4_s_g_near:2'b0);
   assign  sg_out43 = ((_net_1)?_add_map_x_5_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_5_s_g:2'b0);
   assign  sg_out44 = ((_net_1)?_add_map_x_5_s_g:2'b0)|
    ((_net_0)?_add_map_x_5_s_g_near:2'b0);
   assign  sg_out45 = ((_net_1)?_add_map_x_6_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_6_s_g:2'b0);
   assign  sg_out46 = ((_net_1)?_add_map_x_6_s_g:2'b0)|
    ((_net_0)?_add_map_x_6_s_g_near:2'b0);
   assign  sg_out47 = ((_net_1)?_add_map_x_7_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_7_s_g:2'b0);
   assign  sg_out48 = ((_net_1)?_add_map_x_7_s_g:2'b0)|
    ((_net_0)?_add_map_x_7_s_g_near:2'b0);
   assign  sg_out49 = ((_net_1)?_add_map_x_8_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_8_s_g:2'b0);
   assign  sg_out50 = ((_net_1)?_add_map_x_8_s_g:2'b0)|
    ((_net_0)?_add_map_x_8_s_g_near:2'b0);
   assign  sg_out51 = ((_net_1)?_add_map_x_9_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_9_s_g:2'b0);
   assign  sg_out52 = ((_net_1)?_add_map_x_9_s_g:2'b0)|
    ((_net_0)?_add_map_x_9_s_g_near:2'b0);
   assign  sg_out53 = ((_net_1)?_add_map_x_10_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_10_s_g:2'b0);
   assign  sg_out54 = ((_net_1)?_add_map_x_10_s_g:2'b0)|
    ((_net_0)?_add_map_x_10_s_g_near:2'b0);
   assign  sg_out55 = ((_net_1)?_add_map_x_11_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_11_s_g:2'b0);
   assign  sg_out56 = ((_net_1)?_add_map_x_11_s_g:2'b0)|
    ((_net_0)?_add_map_x_11_s_g_near:2'b0);
   assign  sg_out57 = ((_net_1)?_add_map_x_12_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_12_s_g:2'b0);
   assign  sg_out58 = ((_net_1)?_add_map_x_12_s_g:2'b0)|
    ((_net_0)?_add_map_x_12_s_g_near:2'b0);
   assign  sg_out59 = ((_net_1)?_add_map_x_13_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_13_s_g:2'b0);
   assign  sg_out60 = ((_net_1)?_add_map_x_13_s_g:2'b0)|
    ((_net_0)?_add_map_x_13_s_g_near:2'b0);
   assign  sg_out61 = ((_net_1)?_add_map_x_14_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_14_s_g:2'b0);
   assign  sg_out62 = ((_net_1)?_add_map_x_14_s_g:10'b0)|
    ((_net_0)?_add_map_x_14_s_g_near:10'b0);
   assign  sg_out65 = ((_net_1)?_add_map_x_15_s_g:2'b0)|
    ((_net_0)?_add_map_x_15_s_g_near:2'b0);
   assign  sg_out66 = ((_net_1)?_add_map_x_15_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_15_s_g:2'b0);
   assign  sg_out67 = ((_net_1)?_add_map_x_16_s_g:2'b0)|
    ((_net_0)?_add_map_x_16_s_g_near:2'b0);
   assign  sg_out68 = ((_net_1)?_add_map_x_16_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_16_s_g:2'b0);
   assign  sg_out69 = ((_net_1)?_add_map_x_17_s_g:2'b0)|
    ((_net_0)?_add_map_x_17_s_g_near:2'b0);
   assign  sg_out70 = ((_net_1)?_add_map_x_17_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_17_s_g:2'b0);
   assign  sg_out71 = ((_net_1)?_add_map_x_18_s_g:2'b0)|
    ((_net_0)?_add_map_x_18_s_g_near:2'b0);
   assign  sg_out72 = ((_net_1)?_add_map_x_18_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_18_s_g:2'b0);
   assign  sg_out73 = ((_net_1)?_add_map_x_19_s_g:2'b0)|
    ((_net_0)?_add_map_x_19_s_g_near:2'b0);
   assign  sg_out74 = ((_net_1)?_add_map_x_19_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_19_s_g:2'b0);
   assign  sg_out75 = ((_net_1)?_add_map_x_20_s_g:2'b0)|
    ((_net_0)?_add_map_x_20_s_g_near:2'b0);
   assign  sg_out76 = ((_net_1)?_add_map_x_20_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_20_s_g:2'b0);
   assign  sg_out77 = ((_net_1)?_add_map_x_21_s_g:2'b0)|
    ((_net_0)?_add_map_x_21_s_g_near:2'b0);
   assign  sg_out78 = ((_net_1)?_add_map_x_21_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_21_s_g:2'b0);
   assign  sg_out79 = ((_net_1)?_add_map_x_22_s_g:2'b0)|
    ((_net_0)?_add_map_x_22_s_g_near:2'b0);
   assign  sg_out80 = ((_net_1)?_add_map_x_22_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_22_s_g:2'b0);
   assign  sg_out81 = ((_net_1)?_add_map_x_23_s_g:2'b0)|
    ((_net_0)?_add_map_x_23_s_g_near:2'b0);
   assign  sg_out82 = ((_net_1)?_add_map_x_23_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_23_s_g:2'b0);
   assign  sg_out83 = ((_net_1)?_add_map_x_24_s_g:2'b0)|
    ((_net_0)?_add_map_x_24_s_g_near:2'b0);
   assign  sg_out84 = ((_net_1)?_add_map_x_24_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_24_s_g:2'b0);
   assign  sg_out85 = ((_net_1)?_add_map_x_25_s_g:2'b0)|
    ((_net_0)?_add_map_x_25_s_g_near:2'b0);
   assign  sg_out86 = ((_net_1)?_add_map_x_25_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_25_s_g:2'b0);
   assign  sg_out87 = ((_net_1)?_add_map_x_26_s_g:2'b0)|
    ((_net_0)?_add_map_x_26_s_g_near:2'b0);
   assign  sg_out88 = ((_net_1)?_add_map_x_26_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_26_s_g:2'b0);
   assign  sg_out89 = ((_net_1)?_add_map_x_27_s_g:2'b0)|
    ((_net_0)?_add_map_x_27_s_g_near:2'b0);
   assign  sg_out90 = ((_net_1)?_add_map_x_27_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_27_s_g:2'b0);
   assign  sg_out91 = ((_net_1)?_add_map_x_28_s_g:2'b0)|
    ((_net_0)?_add_map_x_28_s_g_near:2'b0);
   assign  sg_out92 = ((_net_1)?_add_map_x_28_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_28_s_g:2'b0);
   assign  sg_out93 = ((_net_1)?_add_map_x_29_s_g:2'b0)|
    ((_net_0)?_add_map_x_29_s_g_near:2'b0);
   assign  sg_out94 = ((_net_1)?_add_map_x_29_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_29_s_g:2'b0);
   assign  sg_out97 = ((_net_1)?_add_map_x_30_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_30_s_g:2'b0);
   assign  sg_out98 = ((_net_1)?_add_map_x_30_s_g:2'b0)|
    ((_net_0)?_add_map_x_30_s_g_near:2'b0);
   assign  sg_out99 = ((_net_1)?_add_map_x_31_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_31_s_g:2'b0);
   assign  sg_out100 = ((_net_1)?_add_map_x_31_s_g:2'b0)|
    ((_net_0)?_add_map_x_31_s_g_near:2'b0);
   assign  sg_out101 = ((_net_1)?_add_map_x_32_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_32_s_g:2'b0);
   assign  sg_out102 = ((_net_1)?_add_map_x_32_s_g:2'b0)|
    ((_net_0)?_add_map_x_32_s_g_near:2'b0);
   assign  sg_out103 = ((_net_1)?_add_map_x_33_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_33_s_g:2'b0);
   assign  sg_out104 = ((_net_1)?_add_map_x_33_s_g:2'b0)|
    ((_net_0)?_add_map_x_33_s_g_near:2'b0);
   assign  sg_out105 = ((_net_1)?_add_map_x_34_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_34_s_g:2'b0);
   assign  sg_out106 = ((_net_1)?_add_map_x_34_s_g:2'b0)|
    ((_net_0)?_add_map_x_34_s_g_near:2'b0);
   assign  sg_out107 = ((_net_1)?_add_map_x_35_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_35_s_g:2'b0);
   assign  sg_out108 = ((_net_1)?_add_map_x_35_s_g:2'b0)|
    ((_net_0)?_add_map_x_35_s_g_near:2'b0);
   assign  sg_out109 = ((_net_1)?_add_map_x_36_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_36_s_g:2'b0);
   assign  sg_out110 = ((_net_1)?_add_map_x_36_s_g:2'b0)|
    ((_net_0)?_add_map_x_36_s_g_near:2'b0);
   assign  sg_out111 = ((_net_1)?_add_map_x_37_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_37_s_g:2'b0);
   assign  sg_out112 = ((_net_1)?_add_map_x_37_s_g:2'b0)|
    ((_net_0)?_add_map_x_37_s_g_near:2'b0);
   assign  sg_out113 = ((_net_1)?_add_map_x_38_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_38_s_g:2'b0);
   assign  sg_out114 = ((_net_1)?_add_map_x_38_s_g:2'b0)|
    ((_net_0)?_add_map_x_38_s_g_near:2'b0);
   assign  sg_out115 = ((_net_1)?_add_map_x_39_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_39_s_g:2'b0);
   assign  sg_out116 = ((_net_1)?_add_map_x_39_s_g:2'b0)|
    ((_net_0)?_add_map_x_39_s_g_near:2'b0);
   assign  sg_out117 = ((_net_1)?_add_map_x_40_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_40_s_g:2'b0);
   assign  sg_out118 = ((_net_1)?_add_map_x_40_s_g:2'b0)|
    ((_net_0)?_add_map_x_40_s_g_near:2'b0);
   assign  sg_out119 = ((_net_1)?_add_map_x_41_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_41_s_g:2'b0);
   assign  sg_out120 = ((_net_1)?_add_map_x_41_s_g:2'b0)|
    ((_net_0)?_add_map_x_41_s_g_near:2'b0);
   assign  sg_out121 = ((_net_1)?_add_map_x_42_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_42_s_g:2'b0);
   assign  sg_out122 = ((_net_1)?_add_map_x_42_s_g:2'b0)|
    ((_net_0)?_add_map_x_42_s_g_near:2'b0);
   assign  sg_out123 = ((_net_1)?_add_map_x_43_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_43_s_g:2'b0);
   assign  sg_out124 = ((_net_1)?_add_map_x_43_s_g:2'b0)|
    ((_net_0)?_add_map_x_43_s_g_near:2'b0);
   assign  sg_out125 = ((_net_1)?_add_map_x_44_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_44_s_g:2'b0);
   assign  sg_out126 = ((_net_1)?_add_map_x_44_s_g:2'b0)|
    ((_net_0)?_add_map_x_44_s_g_near:2'b0);
   assign  sg_out129 = ((_net_1)?_add_map_x_45_s_g:2'b0)|
    ((_net_0)?_add_map_x_45_s_g_near:2'b0);
   assign  sg_out130 = ((_net_1)?_add_map_x_45_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_45_s_g:2'b0);
   assign  sg_out131 = ((_net_1)?_add_map_x_46_s_g:2'b0)|
    ((_net_0)?_add_map_x_46_s_g_near:2'b0);
   assign  sg_out132 = ((_net_1)?_add_map_x_46_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_46_s_g:2'b0);
   assign  sg_out133 = ((_net_1)?_add_map_x_47_s_g:2'b0)|
    ((_net_0)?_add_map_x_47_s_g_near:2'b0);
   assign  sg_out134 = ((_net_1)?_add_map_x_47_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_47_s_g:2'b0);
   assign  sg_out135 = ((_net_1)?_add_map_x_48_s_g:2'b0)|
    ((_net_0)?_add_map_x_48_s_g_near:2'b0);
   assign  sg_out136 = ((_net_1)?_add_map_x_48_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_48_s_g:2'b0);
   assign  sg_out137 = ((_net_1)?_add_map_x_49_s_g:2'b0)|
    ((_net_0)?_add_map_x_49_s_g_near:2'b0);
   assign  sg_out138 = ((_net_1)?_add_map_x_49_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_49_s_g:2'b0);
   assign  sg_out139 = ((_net_1)?_add_map_x_50_s_g:2'b0)|
    ((_net_0)?_add_map_x_50_s_g_near:2'b0);
   assign  sg_out140 = ((_net_1)?_add_map_x_50_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_50_s_g:2'b0);
   assign  sg_out141 = ((_net_1)?_add_map_x_51_s_g:2'b0)|
    ((_net_0)?_add_map_x_51_s_g_near:2'b0);
   assign  sg_out142 = ((_net_1)?_add_map_x_51_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_51_s_g:2'b0);
   assign  sg_out143 = ((_net_1)?_add_map_x_52_s_g:2'b0)|
    ((_net_0)?_add_map_x_52_s_g_near:2'b0);
   assign  sg_out144 = ((_net_1)?_add_map_x_52_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_52_s_g:2'b0);
   assign  sg_out145 = ((_net_1)?_add_map_x_53_s_g:2'b0)|
    ((_net_0)?_add_map_x_53_s_g_near:2'b0);
   assign  sg_out146 = ((_net_1)?_add_map_x_53_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_53_s_g:2'b0);
   assign  sg_out147 = ((_net_1)?_add_map_x_54_s_g:2'b0)|
    ((_net_0)?_add_map_x_54_s_g_near:2'b0);
   assign  sg_out148 = ((_net_1)?_add_map_x_54_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_54_s_g:2'b0);
   assign  sg_out149 = ((_net_1)?_add_map_x_55_s_g:2'b0)|
    ((_net_0)?_add_map_x_55_s_g_near:2'b0);
   assign  sg_out150 = ((_net_1)?_add_map_x_55_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_55_s_g:2'b0);
   assign  sg_out151 = ((_net_1)?_add_map_x_56_s_g:2'b0)|
    ((_net_0)?_add_map_x_56_s_g_near:2'b0);
   assign  sg_out152 = ((_net_1)?_add_map_x_56_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_56_s_g:2'b0);
   assign  sg_out153 = ((_net_1)?_add_map_x_57_s_g:2'b0)|
    ((_net_0)?_add_map_x_57_s_g_near:2'b0);
   assign  sg_out154 = ((_net_1)?_add_map_x_57_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_57_s_g:2'b0);
   assign  sg_out155 = ((_net_1)?_add_map_x_58_s_g:2'b0)|
    ((_net_0)?_add_map_x_58_s_g_near:2'b0);
   assign  sg_out156 = ((_net_1)?_add_map_x_58_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_58_s_g:2'b0);
   assign  sg_out157 = ((_net_1)?_add_map_x_59_s_g:2'b0)|
    ((_net_0)?_add_map_x_59_s_g_near:2'b0);
   assign  sg_out158 = ((_net_1)?_add_map_x_59_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_59_s_g:2'b0);
   assign  sg_out161 = ((_net_1)?_add_map_x_60_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_60_s_g:2'b0);
   assign  sg_out162 = ((_net_1)?_add_map_x_60_s_g:2'b0)|
    ((_net_0)?_add_map_x_60_s_g_near:2'b0);
   assign  sg_out163 = ((_net_1)?_add_map_x_61_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_61_s_g:2'b0);
   assign  sg_out164 = ((_net_1)?_add_map_x_61_s_g:2'b0)|
    ((_net_0)?_add_map_x_61_s_g_near:2'b0);
   assign  sg_out165 = ((_net_1)?_add_map_x_62_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_62_s_g:2'b0);
   assign  sg_out166 = ((_net_1)?_add_map_x_62_s_g:2'b0)|
    ((_net_0)?_add_map_x_62_s_g_near:2'b0);
   assign  sg_out167 = ((_net_1)?_add_map_x_63_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_63_s_g:2'b0);
   assign  sg_out168 = ((_net_1)?_add_map_x_63_s_g:2'b0)|
    ((_net_0)?_add_map_x_63_s_g_near:2'b0);
   assign  sg_out169 = ((_net_1)?_add_map_x_64_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_64_s_g:2'b0);
   assign  sg_out170 = ((_net_1)?_add_map_x_64_s_g:2'b0)|
    ((_net_0)?_add_map_x_64_s_g_near:2'b0);
   assign  sg_out171 = ((_net_1)?_add_map_x_65_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_65_s_g:2'b0);
   assign  sg_out172 = ((_net_1)?_add_map_x_65_s_g:2'b0)|
    ((_net_0)?_add_map_x_65_s_g_near:2'b0);
   assign  sg_out173 = ((_net_1)?_add_map_x_66_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_66_s_g:2'b0);
   assign  sg_out174 = ((_net_1)?_add_map_x_66_s_g:2'b0)|
    ((_net_0)?_add_map_x_66_s_g_near:2'b0);
   assign  sg_out175 = ((_net_1)?_add_map_x_67_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_67_s_g:2'b0);
   assign  sg_out176 = ((_net_1)?_add_map_x_67_s_g:2'b0)|
    ((_net_0)?_add_map_x_67_s_g_near:2'b0);
   assign  sg_out177 = ((_net_1)?_add_map_x_68_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_68_s_g:2'b0);
   assign  sg_out178 = ((_net_1)?_add_map_x_68_s_g:2'b0)|
    ((_net_0)?_add_map_x_68_s_g_near:2'b0);
   assign  sg_out179 = ((_net_1)?_add_map_x_69_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_69_s_g:2'b0);
   assign  sg_out180 = ((_net_1)?_add_map_x_69_s_g:2'b0)|
    ((_net_0)?_add_map_x_69_s_g_near:2'b0);
   assign  sg_out181 = ((_net_1)?_add_map_x_70_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_70_s_g:2'b0);
   assign  sg_out182 = ((_net_1)?_add_map_x_70_s_g:2'b0)|
    ((_net_0)?_add_map_x_70_s_g_near:2'b0);
   assign  sg_out183 = ((_net_1)?_add_map_x_71_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_71_s_g:2'b0);
   assign  sg_out184 = ((_net_1)?_add_map_x_71_s_g:2'b0)|
    ((_net_0)?_add_map_x_71_s_g_near:2'b0);
   assign  sg_out185 = ((_net_1)?_add_map_x_72_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_72_s_g:2'b0);
   assign  sg_out186 = ((_net_1)?_add_map_x_72_s_g:2'b0)|
    ((_net_0)?_add_map_x_72_s_g_near:2'b0);
   assign  sg_out187 = ((_net_1)?_add_map_x_73_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_73_s_g:2'b0);
   assign  sg_out188 = ((_net_1)?_add_map_x_73_s_g:2'b0)|
    ((_net_0)?_add_map_x_73_s_g_near:2'b0);
   assign  sg_out189 = ((_net_1)?_add_map_x_74_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_74_s_g:2'b0);
   assign  sg_out190 = ((_net_1)?_add_map_x_74_s_g:2'b0)|
    ((_net_0)?_add_map_x_74_s_g_near:2'b0);
   assign  sg_out193 = ((_net_1)?_add_map_x_75_s_g:2'b0)|
    ((_net_0)?_add_map_x_75_s_g_near:2'b0);
   assign  sg_out194 = ((_net_1)?_add_map_x_75_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_75_s_g:2'b0);
   assign  sg_out195 = ((_net_1)?_add_map_x_76_s_g:2'b0)|
    ((_net_0)?_add_map_x_76_s_g_near:2'b0);
   assign  sg_out196 = ((_net_1)?_add_map_x_76_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_76_s_g:2'b0);
   assign  sg_out197 = ((_net_1)?_add_map_x_77_s_g:2'b0)|
    ((_net_0)?_add_map_x_77_s_g_near:2'b0);
   assign  sg_out198 = ((_net_1)?_add_map_x_77_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_77_s_g:2'b0);
   assign  sg_out199 = ((_net_1)?_add_map_x_78_s_g:2'b0)|
    ((_net_0)?_add_map_x_78_s_g_near:2'b0);
   assign  sg_out200 = ((_net_1)?_add_map_x_78_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_78_s_g:2'b0);
   assign  sg_out201 = ((_net_1)?_add_map_x_79_s_g:2'b0)|
    ((_net_0)?_add_map_x_79_s_g_near:2'b0);
   assign  sg_out202 = ((_net_1)?_add_map_x_79_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_79_s_g:2'b0);
   assign  sg_out203 = ((_net_1)?_add_map_x_80_s_g:2'b0)|
    ((_net_0)?_add_map_x_80_s_g_near:2'b0);
   assign  sg_out204 = ((_net_1)?_add_map_x_80_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_80_s_g:2'b0);
   assign  sg_out205 = ((_net_1)?_add_map_x_81_s_g:2'b0)|
    ((_net_0)?_add_map_x_81_s_g_near:2'b0);
   assign  sg_out206 = ((_net_1)?_add_map_x_81_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_81_s_g:2'b0);
   assign  sg_out207 = ((_net_1)?_add_map_x_82_s_g:2'b0)|
    ((_net_0)?_add_map_x_82_s_g_near:2'b0);
   assign  sg_out208 = ((_net_1)?_add_map_x_82_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_82_s_g:2'b0);
   assign  sg_out209 = ((_net_1)?_add_map_x_83_s_g:2'b0)|
    ((_net_0)?_add_map_x_83_s_g_near:2'b0);
   assign  sg_out210 = ((_net_1)?_add_map_x_83_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_83_s_g:2'b0);
   assign  sg_out211 = ((_net_1)?_add_map_x_84_s_g:2'b0)|
    ((_net_0)?_add_map_x_84_s_g_near:2'b0);
   assign  sg_out212 = ((_net_1)?_add_map_x_84_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_84_s_g:2'b0);
   assign  sg_out213 = ((_net_1)?_add_map_x_85_s_g:2'b0)|
    ((_net_0)?_add_map_x_85_s_g_near:2'b0);
   assign  sg_out214 = ((_net_1)?_add_map_x_85_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_85_s_g:2'b0);
   assign  sg_out215 = ((_net_1)?_add_map_x_86_s_g:2'b0)|
    ((_net_0)?_add_map_x_86_s_g_near:2'b0);
   assign  sg_out216 = ((_net_1)?_add_map_x_86_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_86_s_g:2'b0);
   assign  sg_out217 = ((_net_1)?_add_map_x_87_s_g:2'b0)|
    ((_net_0)?_add_map_x_87_s_g_near:2'b0);
   assign  sg_out218 = ((_net_1)?_add_map_x_87_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_87_s_g:2'b0);
   assign  sg_out219 = ((_net_1)?_add_map_x_88_s_g:2'b0)|
    ((_net_0)?_add_map_x_88_s_g_near:2'b0);
   assign  sg_out220 = ((_net_1)?_add_map_x_88_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_88_s_g:2'b0);
   assign  sg_out221 = ((_net_1)?_add_map_x_89_s_g:2'b0)|
    ((_net_0)?_add_map_x_89_s_g_near:2'b0);
   assign  sg_out222 = ((_net_1)?_add_map_x_89_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_89_s_g:2'b0);
   assign  sg_out225 = ((_net_1)?_add_map_x_90_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_90_s_g:2'b0);
   assign  sg_out226 = ((_net_1)?_add_map_x_90_s_g:2'b0)|
    ((_net_0)?_add_map_x_90_s_g_near:2'b0);
   assign  sg_out227 = ((_net_1)?_add_map_x_91_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_91_s_g:2'b0);
   assign  sg_out228 = ((_net_1)?_add_map_x_91_s_g:2'b0)|
    ((_net_0)?_add_map_x_91_s_g_near:2'b0);
   assign  sg_out229 = ((_net_1)?_add_map_x_92_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_92_s_g:2'b0);
   assign  sg_out230 = ((_net_1)?_add_map_x_92_s_g:2'b0)|
    ((_net_0)?_add_map_x_92_s_g_near:2'b0);
   assign  sg_out231 = ((_net_1)?_add_map_x_93_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_93_s_g:2'b0);
   assign  sg_out232 = ((_net_1)?_add_map_x_93_s_g:2'b0)|
    ((_net_0)?_add_map_x_93_s_g_near:2'b0);
   assign  sg_out233 = ((_net_1)?_add_map_x_94_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_94_s_g:2'b0);
   assign  sg_out234 = ((_net_1)?_add_map_x_94_s_g:2'b0)|
    ((_net_0)?_add_map_x_94_s_g_near:2'b0);
   assign  sg_out235 = ((_net_1)?_add_map_x_95_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_95_s_g:2'b0);
   assign  sg_out236 = ((_net_1)?_add_map_x_95_s_g:2'b0)|
    ((_net_0)?_add_map_x_95_s_g_near:2'b0);
   assign  sg_out237 = ((_net_1)?_add_map_x_96_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_96_s_g:2'b0);
   assign  sg_out238 = ((_net_1)?_add_map_x_96_s_g:2'b0)|
    ((_net_0)?_add_map_x_96_s_g_near:2'b0);
   assign  sg_out239 = ((_net_1)?_add_map_x_97_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_97_s_g:2'b0);
   assign  sg_out240 = ((_net_1)?_add_map_x_97_s_g:2'b0)|
    ((_net_0)?_add_map_x_97_s_g_near:2'b0);
   assign  sg_out241 = ((_net_1)?_add_map_x_98_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_98_s_g:2'b0);
   assign  sg_out242 = ((_net_1)?_add_map_x_98_s_g:2'b0)|
    ((_net_0)?_add_map_x_98_s_g_near:2'b0);
   assign  sg_out243 = ((_net_1)?_add_map_x_99_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_99_s_g:2'b0);
   assign  sg_out244 = ((_net_1)?_add_map_x_99_s_g:2'b0)|
    ((_net_0)?_add_map_x_99_s_g_near:2'b0);
   assign  sg_out245 = ((_net_1)?_add_map_x_100_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_100_s_g:2'b0);
   assign  sg_out246 = ((_net_1)?_add_map_x_100_s_g:2'b0)|
    ((_net_0)?_add_map_x_100_s_g_near:2'b0);
   assign  sg_out247 = ((_net_1)?_add_map_x_101_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_101_s_g:2'b0);
   assign  sg_out248 = ((_net_1)?_add_map_x_101_s_g:2'b0)|
    ((_net_0)?_add_map_x_101_s_g_near:2'b0);
   assign  sg_out249 = ((_net_1)?_add_map_x_102_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_102_s_g:2'b0);
   assign  sg_out250 = ((_net_1)?_add_map_x_102_s_g:2'b0)|
    ((_net_0)?_add_map_x_102_s_g_near:2'b0);
   assign  sg_out251 = ((_net_1)?_add_map_x_103_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_103_s_g:2'b0);
   assign  sg_out252 = ((_net_1)?_add_map_x_103_s_g:2'b0)|
    ((_net_0)?_add_map_x_103_s_g_near:2'b0);
   assign  sg_out253 = ((_net_1)?_add_map_x_104_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_104_s_g:2'b0);
   assign  sg_out254 = ((_net_1)?_add_map_x_104_s_g:2'b0)|
    ((_net_0)?_add_map_x_104_s_g_near:2'b0);
   assign  sg_out257 = ((_net_1)?_add_map_x_105_s_g:2'b0)|
    ((_net_0)?_add_map_x_105_s_g_near:2'b0);
   assign  sg_out258 = ((_net_1)?_add_map_x_105_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_105_s_g:2'b0);
   assign  sg_out259 = ((_net_1)?_add_map_x_106_s_g:2'b0)|
    ((_net_0)?_add_map_x_106_s_g_near:2'b0);
   assign  sg_out260 = ((_net_1)?_add_map_x_106_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_106_s_g:2'b0);
   assign  sg_out261 = ((_net_1)?_add_map_x_107_s_g:2'b0)|
    ((_net_0)?_add_map_x_107_s_g_near:2'b0);
   assign  sg_out262 = ((_net_1)?_add_map_x_107_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_107_s_g:2'b0);
   assign  sg_out263 = ((_net_1)?_add_map_x_108_s_g:2'b0)|
    ((_net_0)?_add_map_x_108_s_g_near:2'b0);
   assign  sg_out264 = ((_net_1)?_add_map_x_108_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_108_s_g:2'b0);
   assign  sg_out265 = ((_net_1)?_add_map_x_109_s_g:2'b0)|
    ((_net_0)?_add_map_x_109_s_g_near:2'b0);
   assign  sg_out266 = ((_net_1)?_add_map_x_109_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_109_s_g:2'b0);
   assign  sg_out267 = ((_net_1)?_add_map_x_110_s_g:2'b0)|
    ((_net_0)?_add_map_x_110_s_g_near:2'b0);
   assign  sg_out268 = ((_net_1)?_add_map_x_110_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_110_s_g:2'b0);
   assign  sg_out269 = ((_net_1)?_add_map_x_111_s_g:2'b0)|
    ((_net_0)?_add_map_x_111_s_g_near:2'b0);
   assign  sg_out270 = ((_net_1)?_add_map_x_111_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_111_s_g:2'b0);
   assign  sg_out271 = ((_net_1)?_add_map_x_112_s_g:2'b0)|
    ((_net_0)?_add_map_x_112_s_g_near:2'b0);
   assign  sg_out272 = ((_net_1)?_add_map_x_112_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_112_s_g:2'b0);
   assign  sg_out273 = ((_net_1)?_add_map_x_113_s_g:2'b0)|
    ((_net_0)?_add_map_x_113_s_g_near:2'b0);
   assign  sg_out274 = ((_net_1)?_add_map_x_113_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_113_s_g:2'b0);
   assign  sg_out275 = ((_net_1)?_add_map_x_114_s_g:2'b0)|
    ((_net_0)?_add_map_x_114_s_g_near:2'b0);
   assign  sg_out276 = ((_net_1)?_add_map_x_114_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_114_s_g:2'b0);
   assign  sg_out277 = ((_net_1)?_add_map_x_115_s_g:2'b0)|
    ((_net_0)?_add_map_x_115_s_g_near:2'b0);
   assign  sg_out278 = ((_net_1)?_add_map_x_115_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_115_s_g:2'b0);
   assign  sg_out279 = ((_net_1)?_add_map_x_116_s_g:2'b0)|
    ((_net_0)?_add_map_x_116_s_g_near:2'b0);
   assign  sg_out280 = ((_net_1)?_add_map_x_116_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_116_s_g:2'b0);
   assign  sg_out281 = ((_net_1)?_add_map_x_117_s_g:2'b0)|
    ((_net_0)?_add_map_x_117_s_g_near:2'b0);
   assign  sg_out282 = ((_net_1)?_add_map_x_117_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_117_s_g:2'b0);
   assign  sg_out283 = ((_net_1)?_add_map_x_118_s_g:2'b0)|
    ((_net_0)?_add_map_x_118_s_g_near:2'b0);
   assign  sg_out284 = ((_net_1)?_add_map_x_118_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_118_s_g:2'b0);
   assign  sg_out285 = ((_net_1)?_add_map_x_119_s_g:2'b0)|
    ((_net_0)?_add_map_x_119_s_g_near:2'b0);
   assign  sg_out286 = ((_net_1)?_add_map_x_119_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_119_s_g:2'b0);
   assign  sg_out289 = ((_net_1)?_add_map_x_120_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_120_s_g:2'b0);
   assign  sg_out290 = ((_net_1)?_add_map_x_120_s_g:2'b0)|
    ((_net_0)?_add_map_x_120_s_g_near:2'b0);
   assign  sg_out291 = ((_net_1)?_add_map_x_121_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_121_s_g:2'b0);
   assign  sg_out292 = ((_net_1)?_add_map_x_121_s_g:2'b0)|
    ((_net_0)?_add_map_x_121_s_g_near:2'b0);
   assign  sg_out293 = ((_net_1)?_add_map_x_122_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_122_s_g:2'b0);
   assign  sg_out294 = ((_net_1)?_add_map_x_122_s_g:2'b0)|
    ((_net_0)?_add_map_x_122_s_g_near:2'b0);
   assign  sg_out295 = ((_net_1)?_add_map_x_123_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_123_s_g:2'b0);
   assign  sg_out296 = ((_net_1)?_add_map_x_123_s_g:2'b0)|
    ((_net_0)?_add_map_x_123_s_g_near:2'b0);
   assign  sg_out297 = ((_net_1)?_add_map_x_124_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_124_s_g:2'b0);
   assign  sg_out298 = ((_net_1)?_add_map_x_124_s_g:2'b0)|
    ((_net_0)?_add_map_x_124_s_g_near:2'b0);
   assign  sg_out299 = ((_net_1)?_add_map_x_125_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_125_s_g:2'b0);
   assign  sg_out300 = ((_net_1)?_add_map_x_125_s_g:2'b0)|
    ((_net_0)?_add_map_x_125_s_g_near:2'b0);
   assign  sg_out301 = ((_net_1)?_add_map_x_126_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_126_s_g:2'b0);
   assign  sg_out302 = ((_net_1)?_add_map_x_126_s_g:2'b0)|
    ((_net_0)?_add_map_x_126_s_g_near:2'b0);
   assign  sg_out303 = ((_net_1)?_add_map_x_127_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_127_s_g:2'b0);
   assign  sg_out304 = ((_net_1)?_add_map_x_127_s_g:2'b0)|
    ((_net_0)?_add_map_x_127_s_g_near:2'b0);
   assign  sg_out305 = ((_net_1)?_add_map_x_128_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_128_s_g:2'b0);
   assign  sg_out306 = ((_net_1)?_add_map_x_128_s_g:2'b0)|
    ((_net_0)?_add_map_x_128_s_g_near:2'b0);
   assign  sg_out307 = ((_net_1)?_add_map_x_129_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_129_s_g:2'b0);
   assign  sg_out308 = ((_net_1)?_add_map_x_129_s_g:2'b0)|
    ((_net_0)?_add_map_x_129_s_g_near:2'b0);
   assign  sg_out309 = ((_net_1)?_add_map_x_130_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_130_s_g:2'b0);
   assign  sg_out310 = ((_net_1)?_add_map_x_130_s_g:2'b0)|
    ((_net_0)?_add_map_x_130_s_g_near:2'b0);
   assign  sg_out311 = ((_net_1)?_add_map_x_131_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_131_s_g:2'b0);
   assign  sg_out312 = ((_net_1)?_add_map_x_131_s_g:2'b0)|
    ((_net_0)?_add_map_x_131_s_g_near:2'b0);
   assign  sg_out313 = ((_net_1)?_add_map_x_132_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_132_s_g:2'b0);
   assign  sg_out314 = ((_net_1)?_add_map_x_132_s_g:2'b0)|
    ((_net_0)?_add_map_x_132_s_g_near:2'b0);
   assign  sg_out315 = ((_net_1)?_add_map_x_133_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_133_s_g:2'b0);
   assign  sg_out316 = ((_net_1)?_add_map_x_133_s_g:2'b0)|
    ((_net_0)?_add_map_x_133_s_g_near:2'b0);
   assign  sg_out317 = ((_net_1)?_add_map_x_134_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_134_s_g:2'b0);
   assign  sg_out318 = ((_net_1)?_add_map_x_134_s_g:2'b0)|
    ((_net_0)?_add_map_x_134_s_g_near:2'b0);
   assign  sg_out321 = ((_net_1)?_add_map_x_135_s_g:2'b0)|
    ((_net_0)?_add_map_x_135_s_g_near:2'b0);
   assign  sg_out322 = ((_net_1)?_add_map_x_135_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_135_s_g:2'b0);
   assign  sg_out323 = ((_net_1)?_add_map_x_136_s_g:2'b0)|
    ((_net_0)?_add_map_x_136_s_g_near:2'b0);
   assign  sg_out324 = ((_net_1)?_add_map_x_136_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_136_s_g:2'b0);
   assign  sg_out325 = ((_net_1)?_add_map_x_137_s_g:2'b0)|
    ((_net_0)?_add_map_x_137_s_g_near:2'b0);
   assign  sg_out326 = ((_net_1)?_add_map_x_137_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_137_s_g:2'b0);
   assign  sg_out327 = ((_net_1)?_add_map_x_138_s_g:2'b0)|
    ((_net_0)?_add_map_x_138_s_g_near:2'b0);
   assign  sg_out328 = ((_net_1)?_add_map_x_138_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_138_s_g:2'b0);
   assign  sg_out329 = ((_net_1)?_add_map_x_139_s_g:2'b0)|
    ((_net_0)?_add_map_x_139_s_g_near:2'b0);
   assign  sg_out330 = ((_net_1)?_add_map_x_139_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_139_s_g:2'b0);
   assign  sg_out331 = ((_net_1)?_add_map_x_140_s_g:2'b0)|
    ((_net_0)?_add_map_x_140_s_g_near:2'b0);
   assign  sg_out332 = ((_net_1)?_add_map_x_140_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_140_s_g:2'b0);
   assign  sg_out333 = ((_net_1)?_add_map_x_141_s_g:2'b0)|
    ((_net_0)?_add_map_x_141_s_g_near:2'b0);
   assign  sg_out334 = ((_net_1)?_add_map_x_141_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_141_s_g:2'b0);
   assign  sg_out335 = ((_net_1)?_add_map_x_142_s_g:2'b0)|
    ((_net_0)?_add_map_x_142_s_g_near:2'b0);
   assign  sg_out336 = ((_net_1)?_add_map_x_142_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_142_s_g:2'b0);
   assign  sg_out337 = ((_net_1)?_add_map_x_143_s_g:2'b0)|
    ((_net_0)?_add_map_x_143_s_g_near:2'b0);
   assign  sg_out338 = ((_net_1)?_add_map_x_143_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_143_s_g:2'b0);
   assign  sg_out339 = ((_net_1)?_add_map_x_144_s_g:2'b0)|
    ((_net_0)?_add_map_x_144_s_g_near:2'b0);
   assign  sg_out340 = ((_net_1)?_add_map_x_144_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_144_s_g:2'b0);
   assign  sg_out341 = ((_net_1)?_add_map_x_145_s_g:2'b0)|
    ((_net_0)?_add_map_x_145_s_g_near:2'b0);
   assign  sg_out342 = ((_net_1)?_add_map_x_145_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_145_s_g:2'b0);
   assign  sg_out343 = ((_net_1)?_add_map_x_146_s_g:2'b0)|
    ((_net_0)?_add_map_x_146_s_g_near:2'b0);
   assign  sg_out344 = ((_net_1)?_add_map_x_146_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_146_s_g:2'b0);
   assign  sg_out345 = ((_net_1)?_add_map_x_147_s_g:2'b0)|
    ((_net_0)?_add_map_x_147_s_g_near:2'b0);
   assign  sg_out346 = ((_net_1)?_add_map_x_147_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_147_s_g:2'b0);
   assign  sg_out347 = ((_net_1)?_add_map_x_148_s_g:2'b0)|
    ((_net_0)?_add_map_x_148_s_g_near:2'b0);
   assign  sg_out348 = ((_net_1)?_add_map_x_148_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_148_s_g:2'b0);
   assign  sg_out349 = ((_net_1)?_add_map_x_149_s_g:2'b0)|
    ((_net_0)?_add_map_x_149_s_g_near:2'b0);
   assign  sg_out350 = ((_net_1)?_add_map_x_149_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_149_s_g:2'b0);
   assign  sg_out353 = ((_net_1)?_add_map_x_150_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_150_s_g:2'b0);
   assign  sg_out354 = ((_net_1)?_add_map_x_150_s_g:2'b0)|
    ((_net_0)?_add_map_x_150_s_g_near:2'b0);
   assign  sg_out355 = ((_net_1)?_add_map_x_151_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_151_s_g:2'b0);
   assign  sg_out356 = ((_net_1)?_add_map_x_151_s_g:2'b0)|
    ((_net_0)?_add_map_x_151_s_g_near:2'b0);
   assign  sg_out357 = ((_net_1)?_add_map_x_152_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_152_s_g:2'b0);
   assign  sg_out358 = ((_net_1)?_add_map_x_152_s_g:2'b0)|
    ((_net_0)?_add_map_x_152_s_g_near:2'b0);
   assign  sg_out359 = ((_net_1)?_add_map_x_153_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_153_s_g:2'b0);
   assign  sg_out360 = ((_net_1)?_add_map_x_153_s_g:2'b0)|
    ((_net_0)?_add_map_x_153_s_g_near:2'b0);
   assign  sg_out361 = ((_net_1)?_add_map_x_154_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_154_s_g:2'b0);
   assign  sg_out362 = ((_net_1)?_add_map_x_154_s_g:2'b0)|
    ((_net_0)?_add_map_x_154_s_g_near:2'b0);
   assign  sg_out363 = ((_net_1)?_add_map_x_155_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_155_s_g:2'b0);
   assign  sg_out364 = ((_net_1)?_add_map_x_155_s_g:2'b0)|
    ((_net_0)?_add_map_x_155_s_g_near:2'b0);
   assign  sg_out365 = ((_net_1)?_add_map_x_156_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_156_s_g:2'b0);
   assign  sg_out366 = ((_net_1)?_add_map_x_156_s_g:2'b0)|
    ((_net_0)?_add_map_x_156_s_g_near:2'b0);
   assign  sg_out367 = ((_net_1)?_add_map_x_157_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_157_s_g:2'b0);
   assign  sg_out368 = ((_net_1)?_add_map_x_157_s_g:2'b0)|
    ((_net_0)?_add_map_x_157_s_g_near:2'b0);
   assign  sg_out369 = ((_net_1)?_add_map_x_158_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_158_s_g:2'b0);
   assign  sg_out370 = ((_net_1)?_add_map_x_158_s_g:2'b0)|
    ((_net_0)?_add_map_x_158_s_g_near:2'b0);
   assign  sg_out371 = ((_net_1)?_add_map_x_159_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_159_s_g:2'b0);
   assign  sg_out372 = ((_net_1)?_add_map_x_159_s_g:2'b0)|
    ((_net_0)?_add_map_x_159_s_g_near:2'b0);
   assign  sg_out373 = ((_net_1)?_add_map_x_160_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_160_s_g:2'b0);
   assign  sg_out374 = ((_net_1)?_add_map_x_160_s_g:2'b0)|
    ((_net_0)?_add_map_x_160_s_g_near:2'b0);
   assign  sg_out375 = ((_net_1)?_add_map_x_161_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_161_s_g:2'b0);
   assign  sg_out376 = ((_net_1)?_add_map_x_161_s_g:2'b0)|
    ((_net_0)?_add_map_x_161_s_g_near:2'b0);
   assign  sg_out377 = ((_net_1)?_add_map_x_162_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_162_s_g:2'b0);
   assign  sg_out378 = ((_net_1)?_add_map_x_162_s_g:2'b0)|
    ((_net_0)?_add_map_x_162_s_g_near:2'b0);
   assign  sg_out379 = ((_net_1)?_add_map_x_163_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_163_s_g:2'b0);
   assign  sg_out380 = ((_net_1)?_add_map_x_163_s_g:2'b0)|
    ((_net_0)?_add_map_x_163_s_g_near:2'b0);
   assign  sg_out381 = ((_net_1)?_add_map_x_164_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_164_s_g:2'b0);
   assign  sg_out382 = ((_net_1)?_add_map_x_164_s_g:2'b0)|
    ((_net_0)?_add_map_x_164_s_g_near:2'b0);
   assign  sg_out385 = ((_net_1)?_add_map_x_165_s_g:2'b0)|
    ((_net_0)?_add_map_x_165_s_g_near:2'b0);
   assign  sg_out386 = ((_net_1)?_add_map_x_165_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_165_s_g:2'b0);
   assign  sg_out387 = ((_net_1)?_add_map_x_166_s_g:2'b0)|
    ((_net_0)?_add_map_x_166_s_g_near:2'b0);
   assign  sg_out388 = ((_net_1)?_add_map_x_166_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_166_s_g:2'b0);
   assign  sg_out389 = ((_net_1)?_add_map_x_167_s_g:2'b0)|
    ((_net_0)?_add_map_x_167_s_g_near:2'b0);
   assign  sg_out390 = ((_net_1)?_add_map_x_167_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_167_s_g:2'b0);
   assign  sg_out391 = ((_net_1)?_add_map_x_168_s_g:2'b0)|
    ((_net_0)?_add_map_x_168_s_g_near:2'b0);
   assign  sg_out392 = ((_net_1)?_add_map_x_168_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_168_s_g:2'b0);
   assign  sg_out393 = ((_net_1)?_add_map_x_169_s_g:2'b0)|
    ((_net_0)?_add_map_x_169_s_g_near:2'b0);
   assign  sg_out394 = ((_net_1)?_add_map_x_169_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_169_s_g:2'b0);
   assign  sg_out395 = ((_net_1)?_add_map_x_170_s_g:2'b0)|
    ((_net_0)?_add_map_x_170_s_g_near:2'b0);
   assign  sg_out396 = ((_net_1)?_add_map_x_170_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_170_s_g:2'b0);
   assign  sg_out397 = ((_net_1)?_add_map_x_171_s_g:2'b0)|
    ((_net_0)?_add_map_x_171_s_g_near:2'b0);
   assign  sg_out398 = ((_net_1)?_add_map_x_171_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_171_s_g:2'b0);
   assign  sg_out399 = ((_net_1)?_add_map_x_172_s_g:2'b0)|
    ((_net_0)?_add_map_x_172_s_g_near:2'b0);
   assign  sg_out400 = ((_net_1)?_add_map_x_172_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_172_s_g:2'b0);
   assign  sg_out401 = ((_net_1)?_add_map_x_173_s_g:2'b0)|
    ((_net_0)?_add_map_x_173_s_g_near:2'b0);
   assign  sg_out402 = ((_net_1)?_add_map_x_173_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_173_s_g:2'b0);
   assign  sg_out403 = ((_net_1)?_add_map_x_174_s_g:2'b0)|
    ((_net_0)?_add_map_x_174_s_g_near:2'b0);
   assign  sg_out404 = ((_net_1)?_add_map_x_174_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_174_s_g:2'b0);
   assign  sg_out405 = ((_net_1)?_add_map_x_175_s_g:2'b0)|
    ((_net_0)?_add_map_x_175_s_g_near:2'b0);
   assign  sg_out406 = ((_net_1)?_add_map_x_175_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_175_s_g:2'b0);
   assign  sg_out407 = ((_net_1)?_add_map_x_176_s_g:2'b0)|
    ((_net_0)?_add_map_x_176_s_g_near:2'b0);
   assign  sg_out408 = ((_net_1)?_add_map_x_176_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_176_s_g:2'b0);
   assign  sg_out409 = ((_net_1)?_add_map_x_177_s_g:2'b0)|
    ((_net_0)?_add_map_x_177_s_g_near:2'b0);
   assign  sg_out410 = ((_net_1)?_add_map_x_177_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_177_s_g:2'b0);
   assign  sg_out411 = ((_net_1)?_add_map_x_178_s_g:2'b0)|
    ((_net_0)?_add_map_x_178_s_g_near:2'b0);
   assign  sg_out412 = ((_net_1)?_add_map_x_178_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_178_s_g:2'b0);
   assign  sg_out413 = ((_net_1)?_add_map_x_179_s_g:2'b0)|
    ((_net_0)?_add_map_x_179_s_g_near:2'b0);
   assign  sg_out414 = ((_net_1)?_add_map_x_179_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_179_s_g:2'b0);
   assign  sg_out417 = ((_net_1)?_add_map_x_180_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_180_s_g:2'b0);
   assign  sg_out418 = ((_net_1)?_add_map_x_180_s_g:2'b0)|
    ((_net_0)?_add_map_x_180_s_g_near:2'b0);
   assign  sg_out419 = ((_net_1)?_add_map_x_181_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_181_s_g:2'b0);
   assign  sg_out420 = ((_net_1)?_add_map_x_181_s_g:2'b0)|
    ((_net_0)?_add_map_x_181_s_g_near:2'b0);
   assign  sg_out421 = ((_net_1)?_add_map_x_182_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_182_s_g:2'b0);
   assign  sg_out422 = ((_net_1)?_add_map_x_182_s_g:2'b0)|
    ((_net_0)?_add_map_x_182_s_g_near:2'b0);
   assign  sg_out423 = ((_net_1)?_add_map_x_183_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_183_s_g:2'b0);
   assign  sg_out424 = ((_net_1)?_add_map_x_183_s_g:2'b0)|
    ((_net_0)?_add_map_x_183_s_g_near:2'b0);
   assign  sg_out425 = ((_net_1)?_add_map_x_184_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_184_s_g:2'b0);
   assign  sg_out426 = ((_net_1)?_add_map_x_184_s_g:2'b0)|
    ((_net_0)?_add_map_x_184_s_g_near:2'b0);
   assign  sg_out427 = ((_net_1)?_add_map_x_185_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_185_s_g:2'b0);
   assign  sg_out428 = ((_net_1)?_add_map_x_185_s_g:2'b0)|
    ((_net_0)?_add_map_x_185_s_g_near:2'b0);
   assign  sg_out429 = ((_net_1)?_add_map_x_186_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_186_s_g:2'b0);
   assign  sg_out430 = ((_net_1)?_add_map_x_186_s_g:2'b0)|
    ((_net_0)?_add_map_x_186_s_g_near:2'b0);
   assign  sg_out431 = ((_net_1)?_add_map_x_187_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_187_s_g:2'b0);
   assign  sg_out432 = ((_net_1)?_add_map_x_187_s_g:2'b0)|
    ((_net_0)?_add_map_x_187_s_g_near:2'b0);
   assign  sg_out433 = ((_net_1)?_add_map_x_188_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_188_s_g:2'b0);
   assign  sg_out434 = ((_net_1)?_add_map_x_188_s_g:2'b0)|
    ((_net_0)?_add_map_x_188_s_g_near:2'b0);
   assign  sg_out435 = ((_net_1)?_add_map_x_189_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_189_s_g:2'b0);
   assign  sg_out436 = ((_net_1)?_add_map_x_189_s_g:2'b0)|
    ((_net_0)?_add_map_x_189_s_g_near:2'b0);
   assign  sg_out437 = ((_net_1)?_add_map_x_190_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_190_s_g:2'b0);
   assign  sg_out438 = ((_net_1)?_add_map_x_190_s_g:2'b0)|
    ((_net_0)?_add_map_x_190_s_g_near:2'b0);
   assign  sg_out439 = ((_net_1)?_add_map_x_191_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_191_s_g:2'b0);
   assign  sg_out440 = ((_net_1)?_add_map_x_191_s_g:2'b0)|
    ((_net_0)?_add_map_x_191_s_g_near:2'b0);
   assign  sg_out441 = ((_net_1)?_add_map_x_192_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_192_s_g:2'b0);
   assign  sg_out442 = ((_net_1)?_add_map_x_192_s_g:2'b0)|
    ((_net_0)?_add_map_x_192_s_g_near:2'b0);
   assign  sg_out443 = ((_net_1)?_add_map_x_193_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_193_s_g:2'b0);
   assign  sg_out444 = ((_net_1)?_add_map_x_193_s_g:2'b0)|
    ((_net_0)?_add_map_x_193_s_g_near:2'b0);
   assign  sg_out445 = ((_net_1)?_add_map_x_194_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_194_s_g:2'b0);
   assign  sg_out446 = ((_net_1)?_add_map_x_194_s_g:2'b0)|
    ((_net_0)?_add_map_x_194_s_g_near:2'b0);
   assign  sg_out449 = ((_net_1)?_add_map_x_195_s_g:2'b0)|
    ((_net_0)?_add_map_x_195_s_g_near:2'b0);
   assign  sg_out450 = ((_net_1)?_add_map_x_195_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_195_s_g:2'b0);
   assign  sg_out451 = ((_net_1)?_add_map_x_196_s_g:2'b0)|
    ((_net_0)?_add_map_x_196_s_g_near:2'b0);
   assign  sg_out452 = ((_net_1)?_add_map_x_196_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_196_s_g:2'b0);
   assign  sg_out453 = ((_net_1)?_add_map_x_197_s_g:2'b0)|
    ((_net_0)?_add_map_x_197_s_g_near:2'b0);
   assign  sg_out454 = ((_net_1)?_add_map_x_197_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_197_s_g:2'b0);
   assign  sg_out455 = ((_net_1)?_add_map_x_198_s_g:2'b0)|
    ((_net_0)?_add_map_x_198_s_g_near:2'b0);
   assign  sg_out456 = ((_net_1)?_add_map_x_198_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_198_s_g:2'b0);
   assign  sg_out457 = ((_net_1)?_add_map_x_199_s_g:2'b0)|
    ((_net_0)?_add_map_x_199_s_g_near:2'b0);
   assign  sg_out458 = ((_net_1)?_add_map_x_199_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_199_s_g:2'b0);
   assign  sg_out459 = ((_net_1)?_add_map_x_200_s_g:2'b0)|
    ((_net_0)?_add_map_x_200_s_g_near:2'b0);
   assign  sg_out460 = ((_net_1)?_add_map_x_200_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_200_s_g:2'b0);
   assign  sg_out461 = ((_net_1)?_add_map_x_201_s_g:2'b0)|
    ((_net_0)?_add_map_x_201_s_g_near:2'b0);
   assign  sg_out462 = ((_net_1)?_add_map_x_201_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_201_s_g:2'b0);
   assign  sg_out463 = ((_net_1)?_add_map_x_202_s_g:2'b0)|
    ((_net_0)?_add_map_x_202_s_g_near:2'b0);
   assign  sg_out464 = ((_net_1)?_add_map_x_202_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_202_s_g:2'b0);
   assign  sg_out465 = ((_net_1)?_add_map_x_203_s_g:2'b0)|
    ((_net_0)?_add_map_x_203_s_g_near:2'b0);
   assign  sg_out466 = ((_net_1)?_add_map_x_203_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_203_s_g:2'b0);
   assign  sg_out467 = ((_net_1)?_add_map_x_204_s_g:2'b0)|
    ((_net_0)?_add_map_x_204_s_g_near:2'b0);
   assign  sg_out468 = ((_net_1)?_add_map_x_204_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_204_s_g:2'b0);
   assign  sg_out469 = ((_net_1)?_add_map_x_205_s_g:2'b0)|
    ((_net_0)?_add_map_x_205_s_g_near:2'b0);
   assign  sg_out470 = ((_net_1)?_add_map_x_205_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_205_s_g:2'b0);
   assign  sg_out471 = ((_net_1)?_add_map_x_206_s_g:2'b0)|
    ((_net_0)?_add_map_x_206_s_g_near:2'b0);
   assign  sg_out472 = ((_net_1)?_add_map_x_206_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_206_s_g:2'b0);
   assign  sg_out473 = ((_net_1)?_add_map_x_207_s_g:2'b0)|
    ((_net_0)?_add_map_x_207_s_g_near:2'b0);
   assign  sg_out474 = ((_net_1)?_add_map_x_207_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_207_s_g:2'b0);
   assign  sg_out475 = ((_net_1)?_add_map_x_208_s_g:2'b0)|
    ((_net_0)?_add_map_x_208_s_g_near:2'b0);
   assign  sg_out476 = ((_net_1)?_add_map_x_208_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_208_s_g:2'b0);
   assign  sg_out477 = ((_net_1)?_add_map_x_209_s_g:2'b0)|
    ((_net_0)?_add_map_x_209_s_g_near:2'b0);
   assign  sg_out478 = ((_net_1)?_add_map_x_209_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_209_s_g:2'b0);
   assign  dig_t0 = _add_map_x_wall_t_out;
   assign  dig_t1 = _add_map_x_1_wall_t_out;
   assign  dig_t2 = _add_map_x_2_wall_t_out;
   assign  dig_t3 = _add_map_x_3_wall_t_out;
   assign  dig_t4 = _add_map_x_4_wall_t_out;
   assign  dig_t5 = _add_map_x_5_wall_t_out;
   assign  dig_t6 = _add_map_x_6_wall_t_out;
   assign  dig_t7 = _add_map_x_7_wall_t_out;
   assign  dig_t8 = _add_map_x_8_wall_t_out;
   assign  dig_t9 = _add_map_x_9_wall_t_out;
   assign  dig_t10 = _add_map_x_10_wall_t_out;
   assign  dig_t11 = _add_map_x_11_wall_t_out;
   assign  dig_t12 = _add_map_x_12_wall_t_out;
   assign  dig_t13 = _add_map_x_13_wall_t_out;
   assign  dig_t14 = _add_map_x_14_wall_t_out;
   assign  dig_t15 = _add_map_x_15_wall_t_out;
   assign  dig_t16 = _add_map_x_16_wall_t_out;
   assign  dig_t17 = _add_map_x_17_wall_t_out;
   assign  dig_t18 = _add_map_x_18_wall_t_out;
   assign  dig_t19 = _add_map_x_19_wall_t_out;
   assign  dig_t20 = _add_map_x_20_wall_t_out;
   assign  dig_t21 = _add_map_x_21_wall_t_out;
   assign  dig_t22 = _add_map_x_22_wall_t_out;
   assign  dig_t23 = _add_map_x_23_wall_t_out;
   assign  dig_t24 = _add_map_x_24_wall_t_out;
   assign  dig_t25 = _add_map_x_25_wall_t_out;
   assign  dig_t26 = _add_map_x_26_wall_t_out;
   assign  dig_t27 = _add_map_x_27_wall_t_out;
   assign  dig_t28 = _add_map_x_28_wall_t_out;
   assign  dig_t29 = _add_map_x_29_wall_t_out;
   assign  dig_t30 = _add_map_x_30_wall_t_out;
   assign  dig_t31 = _add_map_x_31_wall_t_out;
   assign  dig_t32 = _add_map_x_32_wall_t_out;
   assign  dig_t33 = _add_map_x_33_wall_t_out;
   assign  dig_t34 = _add_map_x_34_wall_t_out;
   assign  dig_t35 = _add_map_x_35_wall_t_out;
   assign  dig_t36 = _add_map_x_36_wall_t_out;
   assign  dig_t37 = _add_map_x_37_wall_t_out;
   assign  dig_t38 = _add_map_x_38_wall_t_out;
   assign  dig_t39 = _add_map_x_39_wall_t_out;
   assign  dig_t40 = _add_map_x_40_wall_t_out;
   assign  dig_t41 = _add_map_x_41_wall_t_out;
   assign  dig_t42 = _add_map_x_42_wall_t_out;
   assign  dig_t43 = _add_map_x_43_wall_t_out;
   assign  dig_t44 = _add_map_x_44_wall_t_out;
   assign  dig_t45 = _add_map_x_45_wall_t_out;
   assign  dig_t46 = _add_map_x_46_wall_t_out;
   assign  dig_t47 = _add_map_x_47_wall_t_out;
   assign  dig_t48 = _add_map_x_48_wall_t_out;
   assign  dig_t49 = _add_map_x_49_wall_t_out;
   assign  dig_t50 = _add_map_x_50_wall_t_out;
   assign  dig_t51 = _add_map_x_51_wall_t_out;
   assign  dig_t52 = _add_map_x_52_wall_t_out;
   assign  dig_t53 = _add_map_x_53_wall_t_out;
   assign  dig_t54 = _add_map_x_54_wall_t_out;
   assign  dig_t55 = _add_map_x_55_wall_t_out;
   assign  dig_t56 = _add_map_x_56_wall_t_out;
   assign  dig_t57 = _add_map_x_57_wall_t_out;
   assign  dig_t58 = _add_map_x_58_wall_t_out;
   assign  dig_t59 = _add_map_x_59_wall_t_out;
   assign  dig_t60 = _add_map_x_60_wall_t_out;
   assign  dig_t61 = _add_map_x_61_wall_t_out;
   assign  dig_t62 = _add_map_x_62_wall_t_out;
   assign  dig_t63 = _add_map_x_63_wall_t_out;
   assign  dig_t64 = _add_map_x_64_wall_t_out;
   assign  dig_t65 = _add_map_x_65_wall_t_out;
   assign  dig_t66 = _add_map_x_66_wall_t_out;
   assign  dig_t67 = _add_map_x_67_wall_t_out;
   assign  dig_t68 = _add_map_x_68_wall_t_out;
   assign  dig_t69 = _add_map_x_69_wall_t_out;
   assign  dig_t70 = _add_map_x_70_wall_t_out;
   assign  dig_t71 = _add_map_x_71_wall_t_out;
   assign  dig_t72 = _add_map_x_72_wall_t_out;
   assign  dig_t73 = _add_map_x_73_wall_t_out;
   assign  dig_t74 = _add_map_x_74_wall_t_out;
   assign  dig_t75 = _add_map_x_75_wall_t_out;
   assign  dig_t76 = _add_map_x_76_wall_t_out;
   assign  dig_t77 = _add_map_x_77_wall_t_out;
   assign  dig_t78 = _add_map_x_78_wall_t_out;
   assign  dig_t79 = _add_map_x_79_wall_t_out;
   assign  dig_t80 = _add_map_x_80_wall_t_out;
   assign  dig_t81 = _add_map_x_81_wall_t_out;
   assign  dig_t82 = _add_map_x_82_wall_t_out;
   assign  dig_t83 = _add_map_x_83_wall_t_out;
   assign  dig_t84 = _add_map_x_84_wall_t_out;
   assign  dig_t85 = _add_map_x_85_wall_t_out;
   assign  dig_t86 = _add_map_x_86_wall_t_out;
   assign  dig_t87 = _add_map_x_87_wall_t_out;
   assign  dig_t88 = _add_map_x_88_wall_t_out;
   assign  dig_t89 = _add_map_x_89_wall_t_out;
   assign  dig_t90 = _add_map_x_90_wall_t_out;
   assign  dig_t91 = _add_map_x_91_wall_t_out;
   assign  dig_t92 = _add_map_x_92_wall_t_out;
   assign  dig_t93 = _add_map_x_93_wall_t_out;
   assign  dig_t94 = _add_map_x_94_wall_t_out;
   assign  dig_t95 = _add_map_x_95_wall_t_out;
   assign  dig_t96 = _add_map_x_96_wall_t_out;
   assign  dig_t97 = _add_map_x_97_wall_t_out;
   assign  dig_t98 = _add_map_x_98_wall_t_out;
   assign  dig_t99 = _add_map_x_99_wall_t_out;
   assign  dig_t100 = _add_map_x_100_wall_t_out;
   assign  dig_t101 = _add_map_x_101_wall_t_out;
   assign  dig_t102 = _add_map_x_102_wall_t_out;
   assign  dig_t103 = _add_map_x_103_wall_t_out;
   assign  dig_t104 = _add_map_x_104_wall_t_out;
   assign  dig_t105 = _add_map_x_105_wall_t_out;
   assign  dig_t106 = _add_map_x_106_wall_t_out;
   assign  dig_t107 = _add_map_x_107_wall_t_out;
   assign  dig_t108 = _add_map_x_108_wall_t_out;
   assign  dig_t109 = _add_map_x_109_wall_t_out;
   assign  dig_t110 = _add_map_x_110_wall_t_out;
   assign  dig_t111 = _add_map_x_111_wall_t_out;
   assign  dig_t112 = _add_map_x_112_wall_t_out;
   assign  dig_t113 = _add_map_x_113_wall_t_out;
   assign  dig_t114 = _add_map_x_114_wall_t_out;
   assign  dig_t115 = _add_map_x_115_wall_t_out;
   assign  dig_t116 = _add_map_x_116_wall_t_out;
   assign  dig_t117 = _add_map_x_117_wall_t_out;
   assign  dig_t118 = _add_map_x_118_wall_t_out;
   assign  dig_t119 = _add_map_x_119_wall_t_out;
   assign  dig_t120 = _add_map_x_120_wall_t_out;
   assign  dig_t121 = _add_map_x_121_wall_t_out;
   assign  dig_t122 = _add_map_x_122_wall_t_out;
   assign  dig_t123 = _add_map_x_123_wall_t_out;
   assign  dig_t124 = _add_map_x_124_wall_t_out;
   assign  dig_t125 = _add_map_x_125_wall_t_out;
   assign  dig_t126 = _add_map_x_126_wall_t_out;
   assign  dig_t127 = _add_map_x_127_wall_t_out;
   assign  dig_t128 = _add_map_x_128_wall_t_out;
   assign  dig_t129 = _add_map_x_129_wall_t_out;
   assign  dig_t130 = _add_map_x_130_wall_t_out;
   assign  dig_t131 = _add_map_x_131_wall_t_out;
   assign  dig_t132 = _add_map_x_132_wall_t_out;
   assign  dig_t133 = _add_map_x_133_wall_t_out;
   assign  dig_t134 = _add_map_x_134_wall_t_out;
   assign  dig_t135 = _add_map_x_135_wall_t_out;
   assign  dig_t136 = _add_map_x_136_wall_t_out;
   assign  dig_t137 = _add_map_x_137_wall_t_out;
   assign  dig_t138 = _add_map_x_138_wall_t_out;
   assign  dig_t139 = _add_map_x_139_wall_t_out;
   assign  dig_t140 = _add_map_x_140_wall_t_out;
   assign  dig_t141 = _add_map_x_141_wall_t_out;
   assign  dig_t142 = _add_map_x_142_wall_t_out;
   assign  dig_t143 = _add_map_x_143_wall_t_out;
   assign  dig_t144 = _add_map_x_144_wall_t_out;
   assign  dig_t145 = _add_map_x_145_wall_t_out;
   assign  dig_t146 = _add_map_x_146_wall_t_out;
   assign  dig_t147 = _add_map_x_147_wall_t_out;
   assign  dig_t148 = _add_map_x_148_wall_t_out;
   assign  dig_t149 = _add_map_x_149_wall_t_out;
   assign  dig_t150 = _add_map_x_150_wall_t_out;
   assign  dig_t151 = _add_map_x_151_wall_t_out;
   assign  dig_t152 = _add_map_x_152_wall_t_out;
   assign  dig_t153 = _add_map_x_153_wall_t_out;
   assign  dig_t154 = _add_map_x_154_wall_t_out;
   assign  dig_t155 = _add_map_x_155_wall_t_out;
   assign  dig_t156 = _add_map_x_156_wall_t_out;
   assign  dig_t157 = _add_map_x_157_wall_t_out;
   assign  dig_t158 = _add_map_x_158_wall_t_out;
   assign  dig_t159 = _add_map_x_159_wall_t_out;
   assign  dig_t160 = _add_map_x_160_wall_t_out;
   assign  dig_t161 = _add_map_x_161_wall_t_out;
   assign  dig_t162 = _add_map_x_162_wall_t_out;
   assign  dig_t163 = _add_map_x_163_wall_t_out;
   assign  dig_t164 = _add_map_x_164_wall_t_out;
   assign  dig_t165 = _add_map_x_165_wall_t_out;
   assign  dig_t166 = _add_map_x_166_wall_t_out;
   assign  dig_t167 = _add_map_x_167_wall_t_out;
   assign  dig_t168 = _add_map_x_168_wall_t_out;
   assign  dig_t169 = _add_map_x_169_wall_t_out;
   assign  dig_t170 = _add_map_x_170_wall_t_out;
   assign  dig_t171 = _add_map_x_171_wall_t_out;
   assign  dig_t172 = _add_map_x_172_wall_t_out;
   assign  dig_t173 = _add_map_x_173_wall_t_out;
   assign  dig_t174 = _add_map_x_174_wall_t_out;
   assign  dig_t175 = _add_map_x_175_wall_t_out;
   assign  dig_t176 = _add_map_x_176_wall_t_out;
   assign  dig_t177 = _add_map_x_177_wall_t_out;
   assign  dig_t178 = _add_map_x_178_wall_t_out;
   assign  dig_t179 = _add_map_x_179_wall_t_out;
   assign  dig_t180 = _add_map_x_180_wall_t_out;
   assign  dig_t181 = _add_map_x_181_wall_t_out;
   assign  dig_t182 = _add_map_x_182_wall_t_out;
   assign  dig_t183 = _add_map_x_183_wall_t_out;
   assign  dig_t184 = _add_map_x_184_wall_t_out;
   assign  dig_t185 = _add_map_x_185_wall_t_out;
   assign  dig_t186 = _add_map_x_186_wall_t_out;
   assign  dig_t187 = _add_map_x_187_wall_t_out;
   assign  dig_t188 = _add_map_x_188_wall_t_out;
   assign  dig_t189 = _add_map_x_189_wall_t_out;
   assign  dig_t190 = _add_map_x_190_wall_t_out;
   assign  dig_t191 = _add_map_x_191_wall_t_out;
   assign  dig_t192 = _add_map_x_192_wall_t_out;
   assign  dig_t193 = _add_map_x_193_wall_t_out;
   assign  dig_t194 = _add_map_x_194_wall_t_out;
   assign  dig_t195 = _add_map_x_195_wall_t_out;
   assign  dig_t196 = _add_map_x_196_wall_t_out;
   assign  dig_t197 = _add_map_x_197_wall_t_out;
   assign  dig_t198 = _add_map_x_198_wall_t_out;
   assign  dig_t199 = _add_map_x_199_wall_t_out;
   assign  dig_t200 = _add_map_x_200_wall_t_out;
   assign  dig_t201 = _add_map_x_201_wall_t_out;
   assign  dig_t202 = _add_map_x_202_wall_t_out;
   assign  dig_t203 = _add_map_x_203_wall_t_out;
   assign  dig_t204 = _add_map_x_204_wall_t_out;
   assign  dig_t205 = _add_map_x_205_wall_t_out;
   assign  dig_t206 = _add_map_x_206_wall_t_out;
   assign  dig_t207 = _add_map_x_207_wall_t_out;
   assign  dig_t208 = _add_map_x_208_wall_t_out;
   assign  dig_t209 = _add_map_x_209_wall_t_out;
   assign  out_do = (_net_7985|_net_3993);
   assign  out_data = (_net_1|_net_0);
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     sig_reg <= 1'b0;
else if ((in_do)) 
      sig_reg <= sig;
end
endmodule

/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 14:47:42 2023
 Licensed to :EVALUATION USER*/
