
/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 14:47:40 2023
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module seach ( p_reset , m_clock , data_in33 , data_in34 , data_in35 , data_in36 , data_in37 , data_in38 , data_in39 , data_in40 , data_in41 , data_in42 , data_in43 , data_in44 , data_in45 , data_in46 , data_in47 , data_in48 , data_in49 , data_in50 , data_in51 , data_in52 , data_in53 , data_in54 , data_in55 , data_in56 , data_in57 , data_in58 , data_in59 , data_in60 , data_in61 , data_in62 , data_in65 , data_in66 , data_in67 , data_in68 , data_in69 , data_in70 , data_in71 , data_in72 , data_in73 , data_in74 , data_in75 , data_in76 , data_in77 , data_in78 , data_in79 , data_in80 , data_in81 , data_in82 , data_in83 , data_in84 , data_in85 , data_in86 , data_in87 , data_in88 , data_in89 , data_in90 , data_in91 , data_in92 , data_in93 , data_in94 , data_in97 , data_in98 , data_in99 , data_in100 , data_in101 , data_in102 , data_in103 , data_in104 , data_in105 , data_in106 , data_in107 , data_in108 , data_in109 , data_in110 , data_in111 , data_in112 , data_in113 , data_in114 , data_in115 , data_in116 , data_in117 , data_in118 , data_in119 , data_in120 , data_in121 , data_in122 , data_in123 , data_in124 , data_in125 , data_in126 , data_in129 , data_in130 , data_in131 , data_in132 , data_in133 , data_in134 , data_in135 , data_in136 , data_in137 , data_in138 , data_in139 , data_in140 , data_in141 , data_in142 , data_in143 , data_in144 , data_in145 , data_in146 , data_in147 , data_in148 , data_in149 , data_in150 , data_in151 , data_in152 , data_in153 , data_in154 , data_in155 , data_in156 , data_in157 , data_in158 , data_in161 , data_in162 , data_in163 , data_in164 , data_in165 , data_in166 , data_in167 , data_in168 , data_in169 , data_in170 , data_in171 , data_in172 , data_in173 , data_in174 , data_in175 , data_in176 , data_in177 , data_in178 , data_in179 , data_in180 , data_in181 , data_in182 , data_in183 , data_in184 , data_in185 , data_in186 , data_in187 , data_in188 , data_in189 , data_in190 , data_in193 , data_in194 , data_in195 , data_in196 , data_in197 , data_in198 , data_in199 , data_in200 , data_in201 , data_in202 , data_in203 , data_in204 , data_in205 , data_in206 , data_in207 , data_in208 , data_in209 , data_in210 , data_in211 , data_in212 , data_in213 , data_in214 , data_in215 , data_in216 , data_in217 , data_in218 , data_in219 , data_in220 , data_in221 , data_in222 , data_in225 , data_in226 , data_in227 , data_in228 , data_in229 , data_in230 , data_in231 , data_in232 , data_in233 , data_in234 , data_in235 , data_in236 , data_in237 , data_in238 , data_in239 , data_in240 , data_in241 , data_in242 , data_in243 , data_in244 , data_in245 , data_in246 , data_in247 , data_in248 , data_in249 , data_in250 , data_in251 , data_in252 , data_in253 , data_in254 , data_in257 , data_in258 , data_in259 , data_in260 , data_in261 , data_in262 , data_in263 , data_in264 , data_in265 , data_in266 , data_in267 , data_in268 , data_in269 , data_in270 , data_in271 , data_in272 , data_in273 , data_in274 , data_in275 , data_in276 , data_in277 , data_in278 , data_in279 , data_in280 , data_in281 , data_in282 , data_in283 , data_in284 , data_in285 , data_in286 , data_in289 , data_in290 , data_in291 , data_in292 , data_in293 , data_in294 , data_in295 , data_in296 , data_in297 , data_in298 , data_in299 , data_in300 , data_in301 , data_in302 , data_in303 , data_in304 , data_in305 , data_in306 , data_in307 , data_in308 , data_in309 , data_in310 , data_in311 , data_in312 , data_in313 , data_in314 , data_in315 , data_in316 , data_in317 , data_in318 , data_in321 , data_in322 , data_in323 , data_in324 , data_in325 , data_in326 , data_in327 , data_in328 , data_in329 , data_in330 , data_in331 , data_in332 , data_in333 , data_in334 , data_in335 , data_in336 , data_in337 , data_in338 , data_in339 , data_in340 , data_in341 , data_in342 , data_in343 , data_in344 , data_in345 , data_in346 , data_in347 , data_in348 , data_in349 , data_in350 , data_in353 , data_in354 , data_in355 , data_in356 , data_in357 , data_in358 , data_in359 , data_in360 , data_in361 , data_in362 , data_in363 , data_in364 , data_in365 , data_in366 , data_in367 , data_in368 , data_in369 , data_in370 , data_in371 , data_in372 , data_in373 , data_in374 , data_in375 , data_in376 , data_in377 , data_in378 , data_in379 , data_in380 , data_in381 , data_in382 , data_in385 , data_in386 , data_in387 , data_in388 , data_in389 , data_in390 , data_in391 , data_in392 , data_in393 , data_in394 , data_in395 , data_in396 , data_in397 , data_in398 , data_in399 , data_in400 , data_in401 , data_in402 , data_in403 , data_in404 , data_in405 , data_in406 , data_in407 , data_in408 , data_in409 , data_in410 , data_in411 , data_in412 , data_in413 , data_in414 , data_in417 , data_in418 , data_in419 , data_in420 , data_in421 , data_in422 , data_in423 , data_in424 , data_in425 , data_in426 , data_in427 , data_in428 , data_in429 , data_in430 , data_in431 , data_in432 , data_in433 , data_in434 , data_in435 , data_in436 , data_in437 , data_in438 , data_in439 , data_in440 , data_in441 , data_in442 , data_in443 , data_in444 , data_in445 , data_in446 , data_in449 , data_in450 , data_in451 , data_in452 , data_in453 , data_in454 , data_in455 , data_in456 , data_in457 , data_in458 , data_in459 , data_in460 , data_in461 , data_in462 , data_in463 , data_in464 , data_in465 , data_in466 , data_in467 , data_in468 , data_in469 , data_in470 , data_in471 , data_in472 , data_in473 , data_in474 , data_in475 , data_in476 , data_in477 , data_in478 , data_out33 , data_out34 , data_out35 , data_out36 , data_out37 , data_out38 , data_out39 , data_out40 , data_out41 , data_out42 , data_out43 , data_out44 , data_out45 , data_out46 , data_out47 , data_out48 , data_out49 , data_out50 , data_out51 , data_out52 , data_out53 , data_out54 , data_out55 , data_out56 , data_out57 , data_out58 , data_out59 , data_out60 , data_out61 , data_out62 , data_out65 , data_out66 , data_out67 , data_out68 , data_out69 , data_out70 , data_out71 , data_out72 , data_out73 , data_out74 , data_out75 , data_out76 , data_out77 , data_out78 , data_out79 , data_out80 , data_out81 , data_out82 , data_out83 , data_out84 , data_out85 , data_out86 , data_out87 , data_out88 , data_out89 , data_out90 , data_out91 , data_out92 , data_out93 , data_out94 , data_out97 , data_out98 , data_out99 , data_out100 , data_out101 , data_out102 , data_out103 , data_out104 , data_out105 , data_out106 , data_out107 , data_out108 , data_out109 , data_out110 , data_out111 , data_out112 , data_out113 , data_out114 , data_out115 , data_out116 , data_out117 , data_out118 , data_out119 , data_out120 , data_out121 , data_out122 , data_out123 , data_out124 , data_out125 , data_out126 , data_out129 , data_out130 , data_out131 , data_out132 , data_out133 , data_out134 , data_out135 , data_out136 , data_out137 , data_out138 , data_out139 , data_out140 , data_out141 , data_out142 , data_out143 , data_out144 , data_out145 , data_out146 , data_out147 , data_out148 , data_out149 , data_out150 , data_out151 , data_out152 , data_out153 , data_out154 , data_out155 , data_out156 , data_out157 , data_out158 , data_out161 , data_out162 , data_out163 , data_out164 , data_out165 , data_out166 , data_out167 , data_out168 , data_out169 , data_out170 , data_out171 , data_out172 , data_out173 , data_out174 , data_out175 , data_out176 , data_out177 , data_out178 , data_out179 , data_out180 , data_out181 , data_out182 , data_out183 , data_out184 , data_out185 , data_out186 , data_out187 , data_out188 , data_out189 , data_out190 , data_out193 , data_out194 , data_out195 , data_out196 , data_out197 , data_out198 , data_out199 , data_out200 , data_out201 , data_out202 , data_out203 , data_out204 , data_out205 , data_out206 , data_out207 , data_out208 , data_out209 , data_out210 , data_out211 , data_out212 , data_out213 , data_out214 , data_out215 , data_out216 , data_out217 , data_out218 , data_out219 , data_out220 , data_out221 , data_out222 , data_out225 , data_out226 , data_out227 , data_out228 , data_out229 , data_out230 , data_out231 , data_out232 , data_out233 , data_out234 , data_out235 , data_out236 , data_out237 , data_out238 , data_out239 , data_out240 , data_out241 , data_out242 , data_out243 , data_out244 , data_out245 , data_out246 , data_out247 , data_out248 , data_out249 , data_out250 , data_out251 , data_out252 , data_out253 , data_out254 , data_out257 , data_out258 , data_out259 , data_out260 , data_out261 , data_out262 , data_out263 , data_out264 , data_out265 , data_out266 , data_out267 , data_out268 , data_out269 , data_out270 , data_out271 , data_out272 , data_out273 , data_out274 , data_out275 , data_out276 , data_out277 , data_out278 , data_out279 , data_out280 , data_out281 , data_out282 , data_out283 , data_out284 , data_out285 , data_out286 , data_out289 , data_out290 , data_out291 , data_out292 , data_out293 , data_out294 , data_out295 , data_out296 , data_out297 , data_out298 , data_out299 , data_out300 , data_out301 , data_out302 , data_out303 , data_out304 , data_out305 , data_out306 , data_out307 , data_out308 , data_out309 , data_out310 , data_out311 , data_out312 , data_out313 , data_out314 , data_out315 , data_out316 , data_out317 , data_out318 , data_out321 , data_out322 , data_out323 , data_out324 , data_out325 , data_out326 , data_out327 , data_out328 , data_out329 , data_out330 , data_out331 , data_out332 , data_out333 , data_out334 , data_out335 , data_out336 , data_out337 , data_out338 , data_out339 , data_out340 , data_out341 , data_out342 , data_out343 , data_out344 , data_out345 , data_out346 , data_out347 , data_out348 , data_out349 , data_out350 , data_out353 , data_out354 , data_out355 , data_out356 , data_out357 , data_out358 , data_out359 , data_out360 , data_out361 , data_out362 , data_out363 , data_out364 , data_out365 , data_out366 , data_out367 , data_out368 , data_out369 , data_out370 , data_out371 , data_out372 , data_out373 , data_out374 , data_out375 , data_out376 , data_out377 , data_out378 , data_out379 , data_out380 , data_out381 , data_out382 , data_out385 , data_out386 , data_out387 , data_out388 , data_out389 , data_out390 , data_out391 , data_out392 , data_out393 , data_out394 , data_out395 , data_out396 , data_out397 , data_out398 , data_out399 , data_out400 , data_out401 , data_out402 , data_out403 , data_out404 , data_out405 , data_out406 , data_out407 , data_out408 , data_out409 , data_out410 , data_out411 , data_out412 , data_out413 , data_out414 , data_out417 , data_out418 , data_out419 , data_out420 , data_out421 , data_out422 , data_out423 , data_out424 , data_out425 , data_out426 , data_out427 , data_out428 , data_out429 , data_out430 , data_out431 , data_out432 , data_out433 , data_out434 , data_out435 , data_out436 , data_out437 , data_out438 , data_out439 , data_out440 , data_out441 , data_out442 , data_out443 , data_out444 , data_out445 , data_out446 , data_out449 , data_out450 , data_out451 , data_out452 , data_out453 , data_out454 , data_out455 , data_out456 , data_out457 , data_out458 , data_out459 , data_out460 , data_out461 , data_out462 , data_out463 , data_out464 , data_out465 , data_out466 , data_out467 , data_out468 , data_out469 , data_out470 , data_out471 , data_out472 , data_out473 , data_out474 , data_out475 , data_out476 , data_out477 , data_out478 , startplot , goalplot , in_do , out_do , out_data );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input [9:0] data_in33;
  wire [9:0] data_in33;
  input [9:0] data_in34;
  wire [9:0] data_in34;
  input [9:0] data_in35;
  wire [9:0] data_in35;
  input [9:0] data_in36;
  wire [9:0] data_in36;
  input [9:0] data_in37;
  wire [9:0] data_in37;
  input [9:0] data_in38;
  wire [9:0] data_in38;
  input [9:0] data_in39;
  wire [9:0] data_in39;
  input [9:0] data_in40;
  wire [9:0] data_in40;
  input [9:0] data_in41;
  wire [9:0] data_in41;
  input [9:0] data_in42;
  wire [9:0] data_in42;
  input [9:0] data_in43;
  wire [9:0] data_in43;
  input [9:0] data_in44;
  wire [9:0] data_in44;
  input [9:0] data_in45;
  wire [9:0] data_in45;
  input [9:0] data_in46;
  wire [9:0] data_in46;
  input [9:0] data_in47;
  wire [9:0] data_in47;
  input [9:0] data_in48;
  wire [9:0] data_in48;
  input [9:0] data_in49;
  wire [9:0] data_in49;
  input [9:0] data_in50;
  wire [9:0] data_in50;
  input [9:0] data_in51;
  wire [9:0] data_in51;
  input [9:0] data_in52;
  wire [9:0] data_in52;
  input [9:0] data_in53;
  wire [9:0] data_in53;
  input [9:0] data_in54;
  wire [9:0] data_in54;
  input [9:0] data_in55;
  wire [9:0] data_in55;
  input [9:0] data_in56;
  wire [9:0] data_in56;
  input [9:0] data_in57;
  wire [9:0] data_in57;
  input [9:0] data_in58;
  wire [9:0] data_in58;
  input [9:0] data_in59;
  wire [9:0] data_in59;
  input [9:0] data_in60;
  wire [9:0] data_in60;
  input [9:0] data_in61;
  wire [9:0] data_in61;
  input [9:0] data_in62;
  wire [9:0] data_in62;
  input [9:0] data_in65;
  wire [9:0] data_in65;
  input [9:0] data_in66;
  wire [9:0] data_in66;
  input [9:0] data_in67;
  wire [9:0] data_in67;
  input [9:0] data_in68;
  wire [9:0] data_in68;
  input [9:0] data_in69;
  wire [9:0] data_in69;
  input [9:0] data_in70;
  wire [9:0] data_in70;
  input [9:0] data_in71;
  wire [9:0] data_in71;
  input [9:0] data_in72;
  wire [9:0] data_in72;
  input [9:0] data_in73;
  wire [9:0] data_in73;
  input [9:0] data_in74;
  wire [9:0] data_in74;
  input [9:0] data_in75;
  wire [9:0] data_in75;
  input [9:0] data_in76;
  wire [9:0] data_in76;
  input [9:0] data_in77;
  wire [9:0] data_in77;
  input [9:0] data_in78;
  wire [9:0] data_in78;
  input [9:0] data_in79;
  wire [9:0] data_in79;
  input [9:0] data_in80;
  wire [9:0] data_in80;
  input [9:0] data_in81;
  wire [9:0] data_in81;
  input [9:0] data_in82;
  wire [9:0] data_in82;
  input [9:0] data_in83;
  wire [9:0] data_in83;
  input [9:0] data_in84;
  wire [9:0] data_in84;
  input [9:0] data_in85;
  wire [9:0] data_in85;
  input [9:0] data_in86;
  wire [9:0] data_in86;
  input [9:0] data_in87;
  wire [9:0] data_in87;
  input [9:0] data_in88;
  wire [9:0] data_in88;
  input [9:0] data_in89;
  wire [9:0] data_in89;
  input [9:0] data_in90;
  wire [9:0] data_in90;
  input [9:0] data_in91;
  wire [9:0] data_in91;
  input [9:0] data_in92;
  wire [9:0] data_in92;
  input [9:0] data_in93;
  wire [9:0] data_in93;
  input [9:0] data_in94;
  wire [9:0] data_in94;
  input [9:0] data_in97;
  wire [9:0] data_in97;
  input [9:0] data_in98;
  wire [9:0] data_in98;
  input [9:0] data_in99;
  wire [9:0] data_in99;
  input [9:0] data_in100;
  wire [9:0] data_in100;
  input [9:0] data_in101;
  wire [9:0] data_in101;
  input [9:0] data_in102;
  wire [9:0] data_in102;
  input [9:0] data_in103;
  wire [9:0] data_in103;
  input [9:0] data_in104;
  wire [9:0] data_in104;
  input [9:0] data_in105;
  wire [9:0] data_in105;
  input [9:0] data_in106;
  wire [9:0] data_in106;
  input [9:0] data_in107;
  wire [9:0] data_in107;
  input [9:0] data_in108;
  wire [9:0] data_in108;
  input [9:0] data_in109;
  wire [9:0] data_in109;
  input [9:0] data_in110;
  wire [9:0] data_in110;
  input [9:0] data_in111;
  wire [9:0] data_in111;
  input [9:0] data_in112;
  wire [9:0] data_in112;
  input [9:0] data_in113;
  wire [9:0] data_in113;
  input [9:0] data_in114;
  wire [9:0] data_in114;
  input [9:0] data_in115;
  wire [9:0] data_in115;
  input [9:0] data_in116;
  wire [9:0] data_in116;
  input [9:0] data_in117;
  wire [9:0] data_in117;
  input [9:0] data_in118;
  wire [9:0] data_in118;
  input [9:0] data_in119;
  wire [9:0] data_in119;
  input [9:0] data_in120;
  wire [9:0] data_in120;
  input [9:0] data_in121;
  wire [9:0] data_in121;
  input [9:0] data_in122;
  wire [9:0] data_in122;
  input [9:0] data_in123;
  wire [9:0] data_in123;
  input [9:0] data_in124;
  wire [9:0] data_in124;
  input [9:0] data_in125;
  wire [9:0] data_in125;
  input [9:0] data_in126;
  wire [9:0] data_in126;
  input [9:0] data_in129;
  wire [9:0] data_in129;
  input [9:0] data_in130;
  wire [9:0] data_in130;
  input [9:0] data_in131;
  wire [9:0] data_in131;
  input [9:0] data_in132;
  wire [9:0] data_in132;
  input [9:0] data_in133;
  wire [9:0] data_in133;
  input [9:0] data_in134;
  wire [9:0] data_in134;
  input [9:0] data_in135;
  wire [9:0] data_in135;
  input [9:0] data_in136;
  wire [9:0] data_in136;
  input [9:0] data_in137;
  wire [9:0] data_in137;
  input [9:0] data_in138;
  wire [9:0] data_in138;
  input [9:0] data_in139;
  wire [9:0] data_in139;
  input [9:0] data_in140;
  wire [9:0] data_in140;
  input [9:0] data_in141;
  wire [9:0] data_in141;
  input [9:0] data_in142;
  wire [9:0] data_in142;
  input [9:0] data_in143;
  wire [9:0] data_in143;
  input [9:0] data_in144;
  wire [9:0] data_in144;
  input [9:0] data_in145;
  wire [9:0] data_in145;
  input [9:0] data_in146;
  wire [9:0] data_in146;
  input [9:0] data_in147;
  wire [9:0] data_in147;
  input [9:0] data_in148;
  wire [9:0] data_in148;
  input [9:0] data_in149;
  wire [9:0] data_in149;
  input [9:0] data_in150;
  wire [9:0] data_in150;
  input [9:0] data_in151;
  wire [9:0] data_in151;
  input [9:0] data_in152;
  wire [9:0] data_in152;
  input [9:0] data_in153;
  wire [9:0] data_in153;
  input [9:0] data_in154;
  wire [9:0] data_in154;
  input [9:0] data_in155;
  wire [9:0] data_in155;
  input [9:0] data_in156;
  wire [9:0] data_in156;
  input [9:0] data_in157;
  wire [9:0] data_in157;
  input [9:0] data_in158;
  wire [9:0] data_in158;
  input [9:0] data_in161;
  wire [9:0] data_in161;
  input [9:0] data_in162;
  wire [9:0] data_in162;
  input [9:0] data_in163;
  wire [9:0] data_in163;
  input [9:0] data_in164;
  wire [9:0] data_in164;
  input [9:0] data_in165;
  wire [9:0] data_in165;
  input [9:0] data_in166;
  wire [9:0] data_in166;
  input [9:0] data_in167;
  wire [9:0] data_in167;
  input [9:0] data_in168;
  wire [9:0] data_in168;
  input [9:0] data_in169;
  wire [9:0] data_in169;
  input [9:0] data_in170;
  wire [9:0] data_in170;
  input [9:0] data_in171;
  wire [9:0] data_in171;
  input [9:0] data_in172;
  wire [9:0] data_in172;
  input [9:0] data_in173;
  wire [9:0] data_in173;
  input [9:0] data_in174;
  wire [9:0] data_in174;
  input [9:0] data_in175;
  wire [9:0] data_in175;
  input [9:0] data_in176;
  wire [9:0] data_in176;
  input [9:0] data_in177;
  wire [9:0] data_in177;
  input [9:0] data_in178;
  wire [9:0] data_in178;
  input [9:0] data_in179;
  wire [9:0] data_in179;
  input [9:0] data_in180;
  wire [9:0] data_in180;
  input [9:0] data_in181;
  wire [9:0] data_in181;
  input [9:0] data_in182;
  wire [9:0] data_in182;
  input [9:0] data_in183;
  wire [9:0] data_in183;
  input [9:0] data_in184;
  wire [9:0] data_in184;
  input [9:0] data_in185;
  wire [9:0] data_in185;
  input [9:0] data_in186;
  wire [9:0] data_in186;
  input [9:0] data_in187;
  wire [9:0] data_in187;
  input [9:0] data_in188;
  wire [9:0] data_in188;
  input [9:0] data_in189;
  wire [9:0] data_in189;
  input [9:0] data_in190;
  wire [9:0] data_in190;
  input [9:0] data_in193;
  wire [9:0] data_in193;
  input [9:0] data_in194;
  wire [9:0] data_in194;
  input [9:0] data_in195;
  wire [9:0] data_in195;
  input [9:0] data_in196;
  wire [9:0] data_in196;
  input [9:0] data_in197;
  wire [9:0] data_in197;
  input [9:0] data_in198;
  wire [9:0] data_in198;
  input [9:0] data_in199;
  wire [9:0] data_in199;
  input [9:0] data_in200;
  wire [9:0] data_in200;
  input [9:0] data_in201;
  wire [9:0] data_in201;
  input [9:0] data_in202;
  wire [9:0] data_in202;
  input [9:0] data_in203;
  wire [9:0] data_in203;
  input [9:0] data_in204;
  wire [9:0] data_in204;
  input [9:0] data_in205;
  wire [9:0] data_in205;
  input [9:0] data_in206;
  wire [9:0] data_in206;
  input [9:0] data_in207;
  wire [9:0] data_in207;
  input [9:0] data_in208;
  wire [9:0] data_in208;
  input [9:0] data_in209;
  wire [9:0] data_in209;
  input [9:0] data_in210;
  wire [9:0] data_in210;
  input [9:0] data_in211;
  wire [9:0] data_in211;
  input [9:0] data_in212;
  wire [9:0] data_in212;
  input [9:0] data_in213;
  wire [9:0] data_in213;
  input [9:0] data_in214;
  wire [9:0] data_in214;
  input [9:0] data_in215;
  wire [9:0] data_in215;
  input [9:0] data_in216;
  wire [9:0] data_in216;
  input [9:0] data_in217;
  wire [9:0] data_in217;
  input [9:0] data_in218;
  wire [9:0] data_in218;
  input [9:0] data_in219;
  wire [9:0] data_in219;
  input [9:0] data_in220;
  wire [9:0] data_in220;
  input [9:0] data_in221;
  wire [9:0] data_in221;
  input [9:0] data_in222;
  wire [9:0] data_in222;
  input [9:0] data_in225;
  wire [9:0] data_in225;
  input [9:0] data_in226;
  wire [9:0] data_in226;
  input [9:0] data_in227;
  wire [9:0] data_in227;
  input [9:0] data_in228;
  wire [9:0] data_in228;
  input [9:0] data_in229;
  wire [9:0] data_in229;
  input [9:0] data_in230;
  wire [9:0] data_in230;
  input [9:0] data_in231;
  wire [9:0] data_in231;
  input [9:0] data_in232;
  wire [9:0] data_in232;
  input [9:0] data_in233;
  wire [9:0] data_in233;
  input [9:0] data_in234;
  wire [9:0] data_in234;
  input [9:0] data_in235;
  wire [9:0] data_in235;
  input [9:0] data_in236;
  wire [9:0] data_in236;
  input [9:0] data_in237;
  wire [9:0] data_in237;
  input [9:0] data_in238;
  wire [9:0] data_in238;
  input [9:0] data_in239;
  wire [9:0] data_in239;
  input [9:0] data_in240;
  wire [9:0] data_in240;
  input [9:0] data_in241;
  wire [9:0] data_in241;
  input [9:0] data_in242;
  wire [9:0] data_in242;
  input [9:0] data_in243;
  wire [9:0] data_in243;
  input [9:0] data_in244;
  wire [9:0] data_in244;
  input [9:0] data_in245;
  wire [9:0] data_in245;
  input [9:0] data_in246;
  wire [9:0] data_in246;
  input [9:0] data_in247;
  wire [9:0] data_in247;
  input [9:0] data_in248;
  wire [9:0] data_in248;
  input [9:0] data_in249;
  wire [9:0] data_in249;
  input [9:0] data_in250;
  wire [9:0] data_in250;
  input [9:0] data_in251;
  wire [9:0] data_in251;
  input [9:0] data_in252;
  wire [9:0] data_in252;
  input [9:0] data_in253;
  wire [9:0] data_in253;
  input [9:0] data_in254;
  wire [9:0] data_in254;
  input [9:0] data_in257;
  wire [9:0] data_in257;
  input [9:0] data_in258;
  wire [9:0] data_in258;
  input [9:0] data_in259;
  wire [9:0] data_in259;
  input [9:0] data_in260;
  wire [9:0] data_in260;
  input [9:0] data_in261;
  wire [9:0] data_in261;
  input [9:0] data_in262;
  wire [9:0] data_in262;
  input [9:0] data_in263;
  wire [9:0] data_in263;
  input [9:0] data_in264;
  wire [9:0] data_in264;
  input [9:0] data_in265;
  wire [9:0] data_in265;
  input [9:0] data_in266;
  wire [9:0] data_in266;
  input [9:0] data_in267;
  wire [9:0] data_in267;
  input [9:0] data_in268;
  wire [9:0] data_in268;
  input [9:0] data_in269;
  wire [9:0] data_in269;
  input [9:0] data_in270;
  wire [9:0] data_in270;
  input [9:0] data_in271;
  wire [9:0] data_in271;
  input [9:0] data_in272;
  wire [9:0] data_in272;
  input [9:0] data_in273;
  wire [9:0] data_in273;
  input [9:0] data_in274;
  wire [9:0] data_in274;
  input [9:0] data_in275;
  wire [9:0] data_in275;
  input [9:0] data_in276;
  wire [9:0] data_in276;
  input [9:0] data_in277;
  wire [9:0] data_in277;
  input [9:0] data_in278;
  wire [9:0] data_in278;
  input [9:0] data_in279;
  wire [9:0] data_in279;
  input [9:0] data_in280;
  wire [9:0] data_in280;
  input [9:0] data_in281;
  wire [9:0] data_in281;
  input [9:0] data_in282;
  wire [9:0] data_in282;
  input [9:0] data_in283;
  wire [9:0] data_in283;
  input [9:0] data_in284;
  wire [9:0] data_in284;
  input [9:0] data_in285;
  wire [9:0] data_in285;
  input [9:0] data_in286;
  wire [9:0] data_in286;
  input [9:0] data_in289;
  wire [9:0] data_in289;
  input [9:0] data_in290;
  wire [9:0] data_in290;
  input [9:0] data_in291;
  wire [9:0] data_in291;
  input [9:0] data_in292;
  wire [9:0] data_in292;
  input [9:0] data_in293;
  wire [9:0] data_in293;
  input [9:0] data_in294;
  wire [9:0] data_in294;
  input [9:0] data_in295;
  wire [9:0] data_in295;
  input [9:0] data_in296;
  wire [9:0] data_in296;
  input [9:0] data_in297;
  wire [9:0] data_in297;
  input [9:0] data_in298;
  wire [9:0] data_in298;
  input [9:0] data_in299;
  wire [9:0] data_in299;
  input [9:0] data_in300;
  wire [9:0] data_in300;
  input [9:0] data_in301;
  wire [9:0] data_in301;
  input [9:0] data_in302;
  wire [9:0] data_in302;
  input [9:0] data_in303;
  wire [9:0] data_in303;
  input [9:0] data_in304;
  wire [9:0] data_in304;
  input [9:0] data_in305;
  wire [9:0] data_in305;
  input [9:0] data_in306;
  wire [9:0] data_in306;
  input [9:0] data_in307;
  wire [9:0] data_in307;
  input [9:0] data_in308;
  wire [9:0] data_in308;
  input [9:0] data_in309;
  wire [9:0] data_in309;
  input [9:0] data_in310;
  wire [9:0] data_in310;
  input [9:0] data_in311;
  wire [9:0] data_in311;
  input [9:0] data_in312;
  wire [9:0] data_in312;
  input [9:0] data_in313;
  wire [9:0] data_in313;
  input [9:0] data_in314;
  wire [9:0] data_in314;
  input [9:0] data_in315;
  wire [9:0] data_in315;
  input [9:0] data_in316;
  wire [9:0] data_in316;
  input [9:0] data_in317;
  wire [9:0] data_in317;
  input [9:0] data_in318;
  wire [9:0] data_in318;
  input [9:0] data_in321;
  wire [9:0] data_in321;
  input [9:0] data_in322;
  wire [9:0] data_in322;
  input [9:0] data_in323;
  wire [9:0] data_in323;
  input [9:0] data_in324;
  wire [9:0] data_in324;
  input [9:0] data_in325;
  wire [9:0] data_in325;
  input [9:0] data_in326;
  wire [9:0] data_in326;
  input [9:0] data_in327;
  wire [9:0] data_in327;
  input [9:0] data_in328;
  wire [9:0] data_in328;
  input [9:0] data_in329;
  wire [9:0] data_in329;
  input [9:0] data_in330;
  wire [9:0] data_in330;
  input [9:0] data_in331;
  wire [9:0] data_in331;
  input [9:0] data_in332;
  wire [9:0] data_in332;
  input [9:0] data_in333;
  wire [9:0] data_in333;
  input [9:0] data_in334;
  wire [9:0] data_in334;
  input [9:0] data_in335;
  wire [9:0] data_in335;
  input [9:0] data_in336;
  wire [9:0] data_in336;
  input [9:0] data_in337;
  wire [9:0] data_in337;
  input [9:0] data_in338;
  wire [9:0] data_in338;
  input [9:0] data_in339;
  wire [9:0] data_in339;
  input [9:0] data_in340;
  wire [9:0] data_in340;
  input [9:0] data_in341;
  wire [9:0] data_in341;
  input [9:0] data_in342;
  wire [9:0] data_in342;
  input [9:0] data_in343;
  wire [9:0] data_in343;
  input [9:0] data_in344;
  wire [9:0] data_in344;
  input [9:0] data_in345;
  wire [9:0] data_in345;
  input [9:0] data_in346;
  wire [9:0] data_in346;
  input [9:0] data_in347;
  wire [9:0] data_in347;
  input [9:0] data_in348;
  wire [9:0] data_in348;
  input [9:0] data_in349;
  wire [9:0] data_in349;
  input [9:0] data_in350;
  wire [9:0] data_in350;
  input [9:0] data_in353;
  wire [9:0] data_in353;
  input [9:0] data_in354;
  wire [9:0] data_in354;
  input [9:0] data_in355;
  wire [9:0] data_in355;
  input [9:0] data_in356;
  wire [9:0] data_in356;
  input [9:0] data_in357;
  wire [9:0] data_in357;
  input [9:0] data_in358;
  wire [9:0] data_in358;
  input [9:0] data_in359;
  wire [9:0] data_in359;
  input [9:0] data_in360;
  wire [9:0] data_in360;
  input [9:0] data_in361;
  wire [9:0] data_in361;
  input [9:0] data_in362;
  wire [9:0] data_in362;
  input [9:0] data_in363;
  wire [9:0] data_in363;
  input [9:0] data_in364;
  wire [9:0] data_in364;
  input [9:0] data_in365;
  wire [9:0] data_in365;
  input [9:0] data_in366;
  wire [9:0] data_in366;
  input [9:0] data_in367;
  wire [9:0] data_in367;
  input [9:0] data_in368;
  wire [9:0] data_in368;
  input [9:0] data_in369;
  wire [9:0] data_in369;
  input [9:0] data_in370;
  wire [9:0] data_in370;
  input [9:0] data_in371;
  wire [9:0] data_in371;
  input [9:0] data_in372;
  wire [9:0] data_in372;
  input [9:0] data_in373;
  wire [9:0] data_in373;
  input [9:0] data_in374;
  wire [9:0] data_in374;
  input [9:0] data_in375;
  wire [9:0] data_in375;
  input [9:0] data_in376;
  wire [9:0] data_in376;
  input [9:0] data_in377;
  wire [9:0] data_in377;
  input [9:0] data_in378;
  wire [9:0] data_in378;
  input [9:0] data_in379;
  wire [9:0] data_in379;
  input [9:0] data_in380;
  wire [9:0] data_in380;
  input [9:0] data_in381;
  wire [9:0] data_in381;
  input [9:0] data_in382;
  wire [9:0] data_in382;
  input [9:0] data_in385;
  wire [9:0] data_in385;
  input [9:0] data_in386;
  wire [9:0] data_in386;
  input [9:0] data_in387;
  wire [9:0] data_in387;
  input [9:0] data_in388;
  wire [9:0] data_in388;
  input [9:0] data_in389;
  wire [9:0] data_in389;
  input [9:0] data_in390;
  wire [9:0] data_in390;
  input [9:0] data_in391;
  wire [9:0] data_in391;
  input [9:0] data_in392;
  wire [9:0] data_in392;
  input [9:0] data_in393;
  wire [9:0] data_in393;
  input [9:0] data_in394;
  wire [9:0] data_in394;
  input [9:0] data_in395;
  wire [9:0] data_in395;
  input [9:0] data_in396;
  wire [9:0] data_in396;
  input [9:0] data_in397;
  wire [9:0] data_in397;
  input [9:0] data_in398;
  wire [9:0] data_in398;
  input [9:0] data_in399;
  wire [9:0] data_in399;
  input [9:0] data_in400;
  wire [9:0] data_in400;
  input [9:0] data_in401;
  wire [9:0] data_in401;
  input [9:0] data_in402;
  wire [9:0] data_in402;
  input [9:0] data_in403;
  wire [9:0] data_in403;
  input [9:0] data_in404;
  wire [9:0] data_in404;
  input [9:0] data_in405;
  wire [9:0] data_in405;
  input [9:0] data_in406;
  wire [9:0] data_in406;
  input [9:0] data_in407;
  wire [9:0] data_in407;
  input [9:0] data_in408;
  wire [9:0] data_in408;
  input [9:0] data_in409;
  wire [9:0] data_in409;
  input [9:0] data_in410;
  wire [9:0] data_in410;
  input [9:0] data_in411;
  wire [9:0] data_in411;
  input [9:0] data_in412;
  wire [9:0] data_in412;
  input [9:0] data_in413;
  wire [9:0] data_in413;
  input [9:0] data_in414;
  wire [9:0] data_in414;
  input [9:0] data_in417;
  wire [9:0] data_in417;
  input [9:0] data_in418;
  wire [9:0] data_in418;
  input [9:0] data_in419;
  wire [9:0] data_in419;
  input [9:0] data_in420;
  wire [9:0] data_in420;
  input [9:0] data_in421;
  wire [9:0] data_in421;
  input [9:0] data_in422;
  wire [9:0] data_in422;
  input [9:0] data_in423;
  wire [9:0] data_in423;
  input [9:0] data_in424;
  wire [9:0] data_in424;
  input [9:0] data_in425;
  wire [9:0] data_in425;
  input [9:0] data_in426;
  wire [9:0] data_in426;
  input [9:0] data_in427;
  wire [9:0] data_in427;
  input [9:0] data_in428;
  wire [9:0] data_in428;
  input [9:0] data_in429;
  wire [9:0] data_in429;
  input [9:0] data_in430;
  wire [9:0] data_in430;
  input [9:0] data_in431;
  wire [9:0] data_in431;
  input [9:0] data_in432;
  wire [9:0] data_in432;
  input [9:0] data_in433;
  wire [9:0] data_in433;
  input [9:0] data_in434;
  wire [9:0] data_in434;
  input [9:0] data_in435;
  wire [9:0] data_in435;
  input [9:0] data_in436;
  wire [9:0] data_in436;
  input [9:0] data_in437;
  wire [9:0] data_in437;
  input [9:0] data_in438;
  wire [9:0] data_in438;
  input [9:0] data_in439;
  wire [9:0] data_in439;
  input [9:0] data_in440;
  wire [9:0] data_in440;
  input [9:0] data_in441;
  wire [9:0] data_in441;
  input [9:0] data_in442;
  wire [9:0] data_in442;
  input [9:0] data_in443;
  wire [9:0] data_in443;
  input [9:0] data_in444;
  wire [9:0] data_in444;
  input [9:0] data_in445;
  wire [9:0] data_in445;
  input [9:0] data_in446;
  wire [9:0] data_in446;
  input [9:0] data_in449;
  wire [9:0] data_in449;
  input [9:0] data_in450;
  wire [9:0] data_in450;
  input [9:0] data_in451;
  wire [9:0] data_in451;
  input [9:0] data_in452;
  wire [9:0] data_in452;
  input [9:0] data_in453;
  wire [9:0] data_in453;
  input [9:0] data_in454;
  wire [9:0] data_in454;
  input [9:0] data_in455;
  wire [9:0] data_in455;
  input [9:0] data_in456;
  wire [9:0] data_in456;
  input [9:0] data_in457;
  wire [9:0] data_in457;
  input [9:0] data_in458;
  wire [9:0] data_in458;
  input [9:0] data_in459;
  wire [9:0] data_in459;
  input [9:0] data_in460;
  wire [9:0] data_in460;
  input [9:0] data_in461;
  wire [9:0] data_in461;
  input [9:0] data_in462;
  wire [9:0] data_in462;
  input [9:0] data_in463;
  wire [9:0] data_in463;
  input [9:0] data_in464;
  wire [9:0] data_in464;
  input [9:0] data_in465;
  wire [9:0] data_in465;
  input [9:0] data_in466;
  wire [9:0] data_in466;
  input [9:0] data_in467;
  wire [9:0] data_in467;
  input [9:0] data_in468;
  wire [9:0] data_in468;
  input [9:0] data_in469;
  wire [9:0] data_in469;
  input [9:0] data_in470;
  wire [9:0] data_in470;
  input [9:0] data_in471;
  wire [9:0] data_in471;
  input [9:0] data_in472;
  wire [9:0] data_in472;
  input [9:0] data_in473;
  wire [9:0] data_in473;
  input [9:0] data_in474;
  wire [9:0] data_in474;
  input [9:0] data_in475;
  wire [9:0] data_in475;
  input [9:0] data_in476;
  wire [9:0] data_in476;
  input [9:0] data_in477;
  wire [9:0] data_in477;
  input [9:0] data_in478;
  wire [9:0] data_in478;
  output [9:0] data_out33;
  wire [9:0] data_out33;
  output [9:0] data_out34;
  wire [9:0] data_out34;
  output [9:0] data_out35;
  wire [9:0] data_out35;
  output [9:0] data_out36;
  wire [9:0] data_out36;
  output [9:0] data_out37;
  wire [9:0] data_out37;
  output [9:0] data_out38;
  wire [9:0] data_out38;
  output [9:0] data_out39;
  wire [9:0] data_out39;
  output [9:0] data_out40;
  wire [9:0] data_out40;
  output [9:0] data_out41;
  wire [9:0] data_out41;
  output [9:0] data_out42;
  wire [9:0] data_out42;
  output [9:0] data_out43;
  wire [9:0] data_out43;
  output [9:0] data_out44;
  wire [9:0] data_out44;
  output [9:0] data_out45;
  wire [9:0] data_out45;
  output [9:0] data_out46;
  wire [9:0] data_out46;
  output [9:0] data_out47;
  wire [9:0] data_out47;
  output [9:0] data_out48;
  wire [9:0] data_out48;
  output [9:0] data_out49;
  wire [9:0] data_out49;
  output [9:0] data_out50;
  wire [9:0] data_out50;
  output [9:0] data_out51;
  wire [9:0] data_out51;
  output [9:0] data_out52;
  wire [9:0] data_out52;
  output [9:0] data_out53;
  wire [9:0] data_out53;
  output [9:0] data_out54;
  wire [9:0] data_out54;
  output [9:0] data_out55;
  wire [9:0] data_out55;
  output [9:0] data_out56;
  wire [9:0] data_out56;
  output [9:0] data_out57;
  wire [9:0] data_out57;
  output [9:0] data_out58;
  wire [9:0] data_out58;
  output [9:0] data_out59;
  wire [9:0] data_out59;
  output [9:0] data_out60;
  wire [9:0] data_out60;
  output [9:0] data_out61;
  wire [9:0] data_out61;
  output [9:0] data_out62;
  wire [9:0] data_out62;
  output [9:0] data_out65;
  wire [9:0] data_out65;
  output [9:0] data_out66;
  wire [9:0] data_out66;
  output [9:0] data_out67;
  wire [9:0] data_out67;
  output [9:0] data_out68;
  wire [9:0] data_out68;
  output [9:0] data_out69;
  wire [9:0] data_out69;
  output [9:0] data_out70;
  wire [9:0] data_out70;
  output [9:0] data_out71;
  wire [9:0] data_out71;
  output [9:0] data_out72;
  wire [9:0] data_out72;
  output [9:0] data_out73;
  wire [9:0] data_out73;
  output [9:0] data_out74;
  wire [9:0] data_out74;
  output [9:0] data_out75;
  wire [9:0] data_out75;
  output [9:0] data_out76;
  wire [9:0] data_out76;
  output [9:0] data_out77;
  wire [9:0] data_out77;
  output [9:0] data_out78;
  wire [9:0] data_out78;
  output [9:0] data_out79;
  wire [9:0] data_out79;
  output [9:0] data_out80;
  wire [9:0] data_out80;
  output [9:0] data_out81;
  wire [9:0] data_out81;
  output [9:0] data_out82;
  wire [9:0] data_out82;
  output [9:0] data_out83;
  wire [9:0] data_out83;
  output [9:0] data_out84;
  wire [9:0] data_out84;
  output [9:0] data_out85;
  wire [9:0] data_out85;
  output [9:0] data_out86;
  wire [9:0] data_out86;
  output [9:0] data_out87;
  wire [9:0] data_out87;
  output [9:0] data_out88;
  wire [9:0] data_out88;
  output [9:0] data_out89;
  wire [9:0] data_out89;
  output [9:0] data_out90;
  wire [9:0] data_out90;
  output [9:0] data_out91;
  wire [9:0] data_out91;
  output [9:0] data_out92;
  wire [9:0] data_out92;
  output [9:0] data_out93;
  wire [9:0] data_out93;
  output [9:0] data_out94;
  wire [9:0] data_out94;
  output [9:0] data_out97;
  wire [9:0] data_out97;
  output [9:0] data_out98;
  wire [9:0] data_out98;
  output [9:0] data_out99;
  wire [9:0] data_out99;
  output [9:0] data_out100;
  wire [9:0] data_out100;
  output [9:0] data_out101;
  wire [9:0] data_out101;
  output [9:0] data_out102;
  wire [9:0] data_out102;
  output [9:0] data_out103;
  wire [9:0] data_out103;
  output [9:0] data_out104;
  wire [9:0] data_out104;
  output [9:0] data_out105;
  wire [9:0] data_out105;
  output [9:0] data_out106;
  wire [9:0] data_out106;
  output [9:0] data_out107;
  wire [9:0] data_out107;
  output [9:0] data_out108;
  wire [9:0] data_out108;
  output [9:0] data_out109;
  wire [9:0] data_out109;
  output [9:0] data_out110;
  wire [9:0] data_out110;
  output [9:0] data_out111;
  wire [9:0] data_out111;
  output [9:0] data_out112;
  wire [9:0] data_out112;
  output [9:0] data_out113;
  wire [9:0] data_out113;
  output [9:0] data_out114;
  wire [9:0] data_out114;
  output [9:0] data_out115;
  wire [9:0] data_out115;
  output [9:0] data_out116;
  wire [9:0] data_out116;
  output [9:0] data_out117;
  wire [9:0] data_out117;
  output [9:0] data_out118;
  wire [9:0] data_out118;
  output [9:0] data_out119;
  wire [9:0] data_out119;
  output [9:0] data_out120;
  wire [9:0] data_out120;
  output [9:0] data_out121;
  wire [9:0] data_out121;
  output [9:0] data_out122;
  wire [9:0] data_out122;
  output [9:0] data_out123;
  wire [9:0] data_out123;
  output [9:0] data_out124;
  wire [9:0] data_out124;
  output [9:0] data_out125;
  wire [9:0] data_out125;
  output [9:0] data_out126;
  wire [9:0] data_out126;
  output [9:0] data_out129;
  wire [9:0] data_out129;
  output [9:0] data_out130;
  wire [9:0] data_out130;
  output [9:0] data_out131;
  wire [9:0] data_out131;
  output [9:0] data_out132;
  wire [9:0] data_out132;
  output [9:0] data_out133;
  wire [9:0] data_out133;
  output [9:0] data_out134;
  wire [9:0] data_out134;
  output [9:0] data_out135;
  wire [9:0] data_out135;
  output [9:0] data_out136;
  wire [9:0] data_out136;
  output [9:0] data_out137;
  wire [9:0] data_out137;
  output [9:0] data_out138;
  wire [9:0] data_out138;
  output [9:0] data_out139;
  wire [9:0] data_out139;
  output [9:0] data_out140;
  wire [9:0] data_out140;
  output [9:0] data_out141;
  wire [9:0] data_out141;
  output [9:0] data_out142;
  wire [9:0] data_out142;
  output [9:0] data_out143;
  wire [9:0] data_out143;
  output [9:0] data_out144;
  wire [9:0] data_out144;
  output [9:0] data_out145;
  wire [9:0] data_out145;
  output [9:0] data_out146;
  wire [9:0] data_out146;
  output [9:0] data_out147;
  wire [9:0] data_out147;
  output [9:0] data_out148;
  wire [9:0] data_out148;
  output [9:0] data_out149;
  wire [9:0] data_out149;
  output [9:0] data_out150;
  wire [9:0] data_out150;
  output [9:0] data_out151;
  wire [9:0] data_out151;
  output [9:0] data_out152;
  wire [9:0] data_out152;
  output [9:0] data_out153;
  wire [9:0] data_out153;
  output [9:0] data_out154;
  wire [9:0] data_out154;
  output [9:0] data_out155;
  wire [9:0] data_out155;
  output [9:0] data_out156;
  wire [9:0] data_out156;
  output [9:0] data_out157;
  wire [9:0] data_out157;
  output [9:0] data_out158;
  wire [9:0] data_out158;
  output [9:0] data_out161;
  wire [9:0] data_out161;
  output [9:0] data_out162;
  wire [9:0] data_out162;
  output [9:0] data_out163;
  wire [9:0] data_out163;
  output [9:0] data_out164;
  wire [9:0] data_out164;
  output [9:0] data_out165;
  wire [9:0] data_out165;
  output [9:0] data_out166;
  wire [9:0] data_out166;
  output [9:0] data_out167;
  wire [9:0] data_out167;
  output [9:0] data_out168;
  wire [9:0] data_out168;
  output [9:0] data_out169;
  wire [9:0] data_out169;
  output [9:0] data_out170;
  wire [9:0] data_out170;
  output [9:0] data_out171;
  wire [9:0] data_out171;
  output [9:0] data_out172;
  wire [9:0] data_out172;
  output [9:0] data_out173;
  wire [9:0] data_out173;
  output [9:0] data_out174;
  wire [9:0] data_out174;
  output [9:0] data_out175;
  wire [9:0] data_out175;
  output [9:0] data_out176;
  wire [9:0] data_out176;
  output [9:0] data_out177;
  wire [9:0] data_out177;
  output [9:0] data_out178;
  wire [9:0] data_out178;
  output [9:0] data_out179;
  wire [9:0] data_out179;
  output [9:0] data_out180;
  wire [9:0] data_out180;
  output [9:0] data_out181;
  wire [9:0] data_out181;
  output [9:0] data_out182;
  wire [9:0] data_out182;
  output [9:0] data_out183;
  wire [9:0] data_out183;
  output [9:0] data_out184;
  wire [9:0] data_out184;
  output [9:0] data_out185;
  wire [9:0] data_out185;
  output [9:0] data_out186;
  wire [9:0] data_out186;
  output [9:0] data_out187;
  wire [9:0] data_out187;
  output [9:0] data_out188;
  wire [9:0] data_out188;
  output [9:0] data_out189;
  wire [9:0] data_out189;
  output [9:0] data_out190;
  wire [9:0] data_out190;
  output [9:0] data_out193;
  wire [9:0] data_out193;
  output [9:0] data_out194;
  wire [9:0] data_out194;
  output [9:0] data_out195;
  wire [9:0] data_out195;
  output [9:0] data_out196;
  wire [9:0] data_out196;
  output [9:0] data_out197;
  wire [9:0] data_out197;
  output [9:0] data_out198;
  wire [9:0] data_out198;
  output [9:0] data_out199;
  wire [9:0] data_out199;
  output [9:0] data_out200;
  wire [9:0] data_out200;
  output [9:0] data_out201;
  wire [9:0] data_out201;
  output [9:0] data_out202;
  wire [9:0] data_out202;
  output [9:0] data_out203;
  wire [9:0] data_out203;
  output [9:0] data_out204;
  wire [9:0] data_out204;
  output [9:0] data_out205;
  wire [9:0] data_out205;
  output [9:0] data_out206;
  wire [9:0] data_out206;
  output [9:0] data_out207;
  wire [9:0] data_out207;
  output [9:0] data_out208;
  wire [9:0] data_out208;
  output [9:0] data_out209;
  wire [9:0] data_out209;
  output [9:0] data_out210;
  wire [9:0] data_out210;
  output [9:0] data_out211;
  wire [9:0] data_out211;
  output [9:0] data_out212;
  wire [9:0] data_out212;
  output [9:0] data_out213;
  wire [9:0] data_out213;
  output [9:0] data_out214;
  wire [9:0] data_out214;
  output [9:0] data_out215;
  wire [9:0] data_out215;
  output [9:0] data_out216;
  wire [9:0] data_out216;
  output [9:0] data_out217;
  wire [9:0] data_out217;
  output [9:0] data_out218;
  wire [9:0] data_out218;
  output [9:0] data_out219;
  wire [9:0] data_out219;
  output [9:0] data_out220;
  wire [9:0] data_out220;
  output [9:0] data_out221;
  wire [9:0] data_out221;
  output [9:0] data_out222;
  wire [9:0] data_out222;
  output [9:0] data_out225;
  wire [9:0] data_out225;
  output [9:0] data_out226;
  wire [9:0] data_out226;
  output [9:0] data_out227;
  wire [9:0] data_out227;
  output [9:0] data_out228;
  wire [9:0] data_out228;
  output [9:0] data_out229;
  wire [9:0] data_out229;
  output [9:0] data_out230;
  wire [9:0] data_out230;
  output [9:0] data_out231;
  wire [9:0] data_out231;
  output [9:0] data_out232;
  wire [9:0] data_out232;
  output [9:0] data_out233;
  wire [9:0] data_out233;
  output [9:0] data_out234;
  wire [9:0] data_out234;
  output [9:0] data_out235;
  wire [9:0] data_out235;
  output [9:0] data_out236;
  wire [9:0] data_out236;
  output [9:0] data_out237;
  wire [9:0] data_out237;
  output [9:0] data_out238;
  wire [9:0] data_out238;
  output [9:0] data_out239;
  wire [9:0] data_out239;
  output [9:0] data_out240;
  wire [9:0] data_out240;
  output [9:0] data_out241;
  wire [9:0] data_out241;
  output [9:0] data_out242;
  wire [9:0] data_out242;
  output [9:0] data_out243;
  wire [9:0] data_out243;
  output [9:0] data_out244;
  wire [9:0] data_out244;
  output [9:0] data_out245;
  wire [9:0] data_out245;
  output [9:0] data_out246;
  wire [9:0] data_out246;
  output [9:0] data_out247;
  wire [9:0] data_out247;
  output [9:0] data_out248;
  wire [9:0] data_out248;
  output [9:0] data_out249;
  wire [9:0] data_out249;
  output [9:0] data_out250;
  wire [9:0] data_out250;
  output [9:0] data_out251;
  wire [9:0] data_out251;
  output [9:0] data_out252;
  wire [9:0] data_out252;
  output [9:0] data_out253;
  wire [9:0] data_out253;
  output [9:0] data_out254;
  wire [9:0] data_out254;
  output [9:0] data_out257;
  wire [9:0] data_out257;
  output [9:0] data_out258;
  wire [9:0] data_out258;
  output [9:0] data_out259;
  wire [9:0] data_out259;
  output [9:0] data_out260;
  wire [9:0] data_out260;
  output [9:0] data_out261;
  wire [9:0] data_out261;
  output [9:0] data_out262;
  wire [9:0] data_out262;
  output [9:0] data_out263;
  wire [9:0] data_out263;
  output [9:0] data_out264;
  wire [9:0] data_out264;
  output [9:0] data_out265;
  wire [9:0] data_out265;
  output [9:0] data_out266;
  wire [9:0] data_out266;
  output [9:0] data_out267;
  wire [9:0] data_out267;
  output [9:0] data_out268;
  wire [9:0] data_out268;
  output [9:0] data_out269;
  wire [9:0] data_out269;
  output [9:0] data_out270;
  wire [9:0] data_out270;
  output [9:0] data_out271;
  wire [9:0] data_out271;
  output [9:0] data_out272;
  wire [9:0] data_out272;
  output [9:0] data_out273;
  wire [9:0] data_out273;
  output [9:0] data_out274;
  wire [9:0] data_out274;
  output [9:0] data_out275;
  wire [9:0] data_out275;
  output [9:0] data_out276;
  wire [9:0] data_out276;
  output [9:0] data_out277;
  wire [9:0] data_out277;
  output [9:0] data_out278;
  wire [9:0] data_out278;
  output [9:0] data_out279;
  wire [9:0] data_out279;
  output [9:0] data_out280;
  wire [9:0] data_out280;
  output [9:0] data_out281;
  wire [9:0] data_out281;
  output [9:0] data_out282;
  wire [9:0] data_out282;
  output [9:0] data_out283;
  wire [9:0] data_out283;
  output [9:0] data_out284;
  wire [9:0] data_out284;
  output [9:0] data_out285;
  wire [9:0] data_out285;
  output [9:0] data_out286;
  wire [9:0] data_out286;
  output [9:0] data_out289;
  wire [9:0] data_out289;
  output [9:0] data_out290;
  wire [9:0] data_out290;
  output [9:0] data_out291;
  wire [9:0] data_out291;
  output [9:0] data_out292;
  wire [9:0] data_out292;
  output [9:0] data_out293;
  wire [9:0] data_out293;
  output [9:0] data_out294;
  wire [9:0] data_out294;
  output [9:0] data_out295;
  wire [9:0] data_out295;
  output [9:0] data_out296;
  wire [9:0] data_out296;
  output [9:0] data_out297;
  wire [9:0] data_out297;
  output [9:0] data_out298;
  wire [9:0] data_out298;
  output [9:0] data_out299;
  wire [9:0] data_out299;
  output [9:0] data_out300;
  wire [9:0] data_out300;
  output [9:0] data_out301;
  wire [9:0] data_out301;
  output [9:0] data_out302;
  wire [9:0] data_out302;
  output [9:0] data_out303;
  wire [9:0] data_out303;
  output [9:0] data_out304;
  wire [9:0] data_out304;
  output [9:0] data_out305;
  wire [9:0] data_out305;
  output [9:0] data_out306;
  wire [9:0] data_out306;
  output [9:0] data_out307;
  wire [9:0] data_out307;
  output [9:0] data_out308;
  wire [9:0] data_out308;
  output [9:0] data_out309;
  wire [9:0] data_out309;
  output [9:0] data_out310;
  wire [9:0] data_out310;
  output [9:0] data_out311;
  wire [9:0] data_out311;
  output [9:0] data_out312;
  wire [9:0] data_out312;
  output [9:0] data_out313;
  wire [9:0] data_out313;
  output [9:0] data_out314;
  wire [9:0] data_out314;
  output [9:0] data_out315;
  wire [9:0] data_out315;
  output [9:0] data_out316;
  wire [9:0] data_out316;
  output [9:0] data_out317;
  wire [9:0] data_out317;
  output [9:0] data_out318;
  wire [9:0] data_out318;
  output [9:0] data_out321;
  wire [9:0] data_out321;
  output [9:0] data_out322;
  wire [9:0] data_out322;
  output [9:0] data_out323;
  wire [9:0] data_out323;
  output [9:0] data_out324;
  wire [9:0] data_out324;
  output [9:0] data_out325;
  wire [9:0] data_out325;
  output [9:0] data_out326;
  wire [9:0] data_out326;
  output [9:0] data_out327;
  wire [9:0] data_out327;
  output [9:0] data_out328;
  wire [9:0] data_out328;
  output [9:0] data_out329;
  wire [9:0] data_out329;
  output [9:0] data_out330;
  wire [9:0] data_out330;
  output [9:0] data_out331;
  wire [9:0] data_out331;
  output [9:0] data_out332;
  wire [9:0] data_out332;
  output [9:0] data_out333;
  wire [9:0] data_out333;
  output [9:0] data_out334;
  wire [9:0] data_out334;
  output [9:0] data_out335;
  wire [9:0] data_out335;
  output [9:0] data_out336;
  wire [9:0] data_out336;
  output [9:0] data_out337;
  wire [9:0] data_out337;
  output [9:0] data_out338;
  wire [9:0] data_out338;
  output [9:0] data_out339;
  wire [9:0] data_out339;
  output [9:0] data_out340;
  wire [9:0] data_out340;
  output [9:0] data_out341;
  wire [9:0] data_out341;
  output [9:0] data_out342;
  wire [9:0] data_out342;
  output [9:0] data_out343;
  wire [9:0] data_out343;
  output [9:0] data_out344;
  wire [9:0] data_out344;
  output [9:0] data_out345;
  wire [9:0] data_out345;
  output [9:0] data_out346;
  wire [9:0] data_out346;
  output [9:0] data_out347;
  wire [9:0] data_out347;
  output [9:0] data_out348;
  wire [9:0] data_out348;
  output [9:0] data_out349;
  wire [9:0] data_out349;
  output [9:0] data_out350;
  wire [9:0] data_out350;
  output [9:0] data_out353;
  wire [9:0] data_out353;
  output [9:0] data_out354;
  wire [9:0] data_out354;
  output [9:0] data_out355;
  wire [9:0] data_out355;
  output [9:0] data_out356;
  wire [9:0] data_out356;
  output [9:0] data_out357;
  wire [9:0] data_out357;
  output [9:0] data_out358;
  wire [9:0] data_out358;
  output [9:0] data_out359;
  wire [9:0] data_out359;
  output [9:0] data_out360;
  wire [9:0] data_out360;
  output [9:0] data_out361;
  wire [9:0] data_out361;
  output [9:0] data_out362;
  wire [9:0] data_out362;
  output [9:0] data_out363;
  wire [9:0] data_out363;
  output [9:0] data_out364;
  wire [9:0] data_out364;
  output [9:0] data_out365;
  wire [9:0] data_out365;
  output [9:0] data_out366;
  wire [9:0] data_out366;
  output [9:0] data_out367;
  wire [9:0] data_out367;
  output [9:0] data_out368;
  wire [9:0] data_out368;
  output [9:0] data_out369;
  wire [9:0] data_out369;
  output [9:0] data_out370;
  wire [9:0] data_out370;
  output [9:0] data_out371;
  wire [9:0] data_out371;
  output [9:0] data_out372;
  wire [9:0] data_out372;
  output [9:0] data_out373;
  wire [9:0] data_out373;
  output [9:0] data_out374;
  wire [9:0] data_out374;
  output [9:0] data_out375;
  wire [9:0] data_out375;
  output [9:0] data_out376;
  wire [9:0] data_out376;
  output [9:0] data_out377;
  wire [9:0] data_out377;
  output [9:0] data_out378;
  wire [9:0] data_out378;
  output [9:0] data_out379;
  wire [9:0] data_out379;
  output [9:0] data_out380;
  wire [9:0] data_out380;
  output [9:0] data_out381;
  wire [9:0] data_out381;
  output [9:0] data_out382;
  wire [9:0] data_out382;
  output [9:0] data_out385;
  wire [9:0] data_out385;
  output [9:0] data_out386;
  wire [9:0] data_out386;
  output [9:0] data_out387;
  wire [9:0] data_out387;
  output [9:0] data_out388;
  wire [9:0] data_out388;
  output [9:0] data_out389;
  wire [9:0] data_out389;
  output [9:0] data_out390;
  wire [9:0] data_out390;
  output [9:0] data_out391;
  wire [9:0] data_out391;
  output [9:0] data_out392;
  wire [9:0] data_out392;
  output [9:0] data_out393;
  wire [9:0] data_out393;
  output [9:0] data_out394;
  wire [9:0] data_out394;
  output [9:0] data_out395;
  wire [9:0] data_out395;
  output [9:0] data_out396;
  wire [9:0] data_out396;
  output [9:0] data_out397;
  wire [9:0] data_out397;
  output [9:0] data_out398;
  wire [9:0] data_out398;
  output [9:0] data_out399;
  wire [9:0] data_out399;
  output [9:0] data_out400;
  wire [9:0] data_out400;
  output [9:0] data_out401;
  wire [9:0] data_out401;
  output [9:0] data_out402;
  wire [9:0] data_out402;
  output [9:0] data_out403;
  wire [9:0] data_out403;
  output [9:0] data_out404;
  wire [9:0] data_out404;
  output [9:0] data_out405;
  wire [9:0] data_out405;
  output [9:0] data_out406;
  wire [9:0] data_out406;
  output [9:0] data_out407;
  wire [9:0] data_out407;
  output [9:0] data_out408;
  wire [9:0] data_out408;
  output [9:0] data_out409;
  wire [9:0] data_out409;
  output [9:0] data_out410;
  wire [9:0] data_out410;
  output [9:0] data_out411;
  wire [9:0] data_out411;
  output [9:0] data_out412;
  wire [9:0] data_out412;
  output [9:0] data_out413;
  wire [9:0] data_out413;
  output [9:0] data_out414;
  wire [9:0] data_out414;
  output [9:0] data_out417;
  wire [9:0] data_out417;
  output [9:0] data_out418;
  wire [9:0] data_out418;
  output [9:0] data_out419;
  wire [9:0] data_out419;
  output [9:0] data_out420;
  wire [9:0] data_out420;
  output [9:0] data_out421;
  wire [9:0] data_out421;
  output [9:0] data_out422;
  wire [9:0] data_out422;
  output [9:0] data_out423;
  wire [9:0] data_out423;
  output [9:0] data_out424;
  wire [9:0] data_out424;
  output [9:0] data_out425;
  wire [9:0] data_out425;
  output [9:0] data_out426;
  wire [9:0] data_out426;
  output [9:0] data_out427;
  wire [9:0] data_out427;
  output [9:0] data_out428;
  wire [9:0] data_out428;
  output [9:0] data_out429;
  wire [9:0] data_out429;
  output [9:0] data_out430;
  wire [9:0] data_out430;
  output [9:0] data_out431;
  wire [9:0] data_out431;
  output [9:0] data_out432;
  wire [9:0] data_out432;
  output [9:0] data_out433;
  wire [9:0] data_out433;
  output [9:0] data_out434;
  wire [9:0] data_out434;
  output [9:0] data_out435;
  wire [9:0] data_out435;
  output [9:0] data_out436;
  wire [9:0] data_out436;
  output [9:0] data_out437;
  wire [9:0] data_out437;
  output [9:0] data_out438;
  wire [9:0] data_out438;
  output [9:0] data_out439;
  wire [9:0] data_out439;
  output [9:0] data_out440;
  wire [9:0] data_out440;
  output [9:0] data_out441;
  wire [9:0] data_out441;
  output [9:0] data_out442;
  wire [9:0] data_out442;
  output [9:0] data_out443;
  wire [9:0] data_out443;
  output [9:0] data_out444;
  wire [9:0] data_out444;
  output [9:0] data_out445;
  wire [9:0] data_out445;
  output [9:0] data_out446;
  wire [9:0] data_out446;
  output [9:0] data_out449;
  wire [9:0] data_out449;
  output [9:0] data_out450;
  wire [9:0] data_out450;
  output [9:0] data_out451;
  wire [9:0] data_out451;
  output [9:0] data_out452;
  wire [9:0] data_out452;
  output [9:0] data_out453;
  wire [9:0] data_out453;
  output [9:0] data_out454;
  wire [9:0] data_out454;
  output [9:0] data_out455;
  wire [9:0] data_out455;
  output [9:0] data_out456;
  wire [9:0] data_out456;
  output [9:0] data_out457;
  wire [9:0] data_out457;
  output [9:0] data_out458;
  wire [9:0] data_out458;
  output [9:0] data_out459;
  wire [9:0] data_out459;
  output [9:0] data_out460;
  wire [9:0] data_out460;
  output [9:0] data_out461;
  wire [9:0] data_out461;
  output [9:0] data_out462;
  wire [9:0] data_out462;
  output [9:0] data_out463;
  wire [9:0] data_out463;
  output [9:0] data_out464;
  wire [9:0] data_out464;
  output [9:0] data_out465;
  wire [9:0] data_out465;
  output [9:0] data_out466;
  wire [9:0] data_out466;
  output [9:0] data_out467;
  wire [9:0] data_out467;
  output [9:0] data_out468;
  wire [9:0] data_out468;
  output [9:0] data_out469;
  wire [9:0] data_out469;
  output [9:0] data_out470;
  wire [9:0] data_out470;
  output [9:0] data_out471;
  wire [9:0] data_out471;
  output [9:0] data_out472;
  wire [9:0] data_out472;
  output [9:0] data_out473;
  wire [9:0] data_out473;
  output [9:0] data_out474;
  wire [9:0] data_out474;
  output [9:0] data_out475;
  wire [9:0] data_out475;
  output [9:0] data_out476;
  wire [9:0] data_out476;
  output [9:0] data_out477;
  wire [9:0] data_out477;
  output [9:0] data_out478;
  wire [9:0] data_out478;
  output [9:0] startplot;
  wire [9:0] startplot;
  output [9:0] goalplot;
  wire [9:0] goalplot;
  input in_do;
  wire in_do;
  output out_do;
  wire out_do;
  output out_data;
  wire out_data;
  reg [9:0] startplot_reg;
  reg [9:0] goalplot_reg;
  wire [9:0] startplot_wire;
  wire [9:0] goalplot_wire;
  wire [9:0] _seach_blockx_map_block;
  wire [9:0] _seach_blockx_now;
  wire [9:0] _seach_blockx_start;
  wire [9:0] _seach_blockx_goal;
  wire [9:0] _seach_blockx_data_out;
  wire _seach_blockx_in_do;
  wire _seach_blockx_p_reset;
  wire _seach_blockx_m_clock;
  wire [9:0] _seach_blockx_419_map_block;
  wire [9:0] _seach_blockx_419_now;
  wire [9:0] _seach_blockx_419_start;
  wire [9:0] _seach_blockx_419_goal;
  wire [9:0] _seach_blockx_419_data_out;
  wire _seach_blockx_419_in_do;
  wire _seach_blockx_419_p_reset;
  wire _seach_blockx_419_m_clock;
  wire [9:0] _seach_blockx_418_map_block;
  wire [9:0] _seach_blockx_418_now;
  wire [9:0] _seach_blockx_418_start;
  wire [9:0] _seach_blockx_418_goal;
  wire [9:0] _seach_blockx_418_data_out;
  wire _seach_blockx_418_in_do;
  wire _seach_blockx_418_p_reset;
  wire _seach_blockx_418_m_clock;
  wire [9:0] _seach_blockx_417_map_block;
  wire [9:0] _seach_blockx_417_now;
  wire [9:0] _seach_blockx_417_start;
  wire [9:0] _seach_blockx_417_goal;
  wire [9:0] _seach_blockx_417_data_out;
  wire _seach_blockx_417_in_do;
  wire _seach_blockx_417_p_reset;
  wire _seach_blockx_417_m_clock;
  wire [9:0] _seach_blockx_416_map_block;
  wire [9:0] _seach_blockx_416_now;
  wire [9:0] _seach_blockx_416_start;
  wire [9:0] _seach_blockx_416_goal;
  wire [9:0] _seach_blockx_416_data_out;
  wire _seach_blockx_416_in_do;
  wire _seach_blockx_416_p_reset;
  wire _seach_blockx_416_m_clock;
  wire [9:0] _seach_blockx_415_map_block;
  wire [9:0] _seach_blockx_415_now;
  wire [9:0] _seach_blockx_415_start;
  wire [9:0] _seach_blockx_415_goal;
  wire [9:0] _seach_blockx_415_data_out;
  wire _seach_blockx_415_in_do;
  wire _seach_blockx_415_p_reset;
  wire _seach_blockx_415_m_clock;
  wire [9:0] _seach_blockx_414_map_block;
  wire [9:0] _seach_blockx_414_now;
  wire [9:0] _seach_blockx_414_start;
  wire [9:0] _seach_blockx_414_goal;
  wire [9:0] _seach_blockx_414_data_out;
  wire _seach_blockx_414_in_do;
  wire _seach_blockx_414_p_reset;
  wire _seach_blockx_414_m_clock;
  wire [9:0] _seach_blockx_413_map_block;
  wire [9:0] _seach_blockx_413_now;
  wire [9:0] _seach_blockx_413_start;
  wire [9:0] _seach_blockx_413_goal;
  wire [9:0] _seach_blockx_413_data_out;
  wire _seach_blockx_413_in_do;
  wire _seach_blockx_413_p_reset;
  wire _seach_blockx_413_m_clock;
  wire [9:0] _seach_blockx_412_map_block;
  wire [9:0] _seach_blockx_412_now;
  wire [9:0] _seach_blockx_412_start;
  wire [9:0] _seach_blockx_412_goal;
  wire [9:0] _seach_blockx_412_data_out;
  wire _seach_blockx_412_in_do;
  wire _seach_blockx_412_p_reset;
  wire _seach_blockx_412_m_clock;
  wire [9:0] _seach_blockx_411_map_block;
  wire [9:0] _seach_blockx_411_now;
  wire [9:0] _seach_blockx_411_start;
  wire [9:0] _seach_blockx_411_goal;
  wire [9:0] _seach_blockx_411_data_out;
  wire _seach_blockx_411_in_do;
  wire _seach_blockx_411_p_reset;
  wire _seach_blockx_411_m_clock;
  wire [9:0] _seach_blockx_410_map_block;
  wire [9:0] _seach_blockx_410_now;
  wire [9:0] _seach_blockx_410_start;
  wire [9:0] _seach_blockx_410_goal;
  wire [9:0] _seach_blockx_410_data_out;
  wire _seach_blockx_410_in_do;
  wire _seach_blockx_410_p_reset;
  wire _seach_blockx_410_m_clock;
  wire [9:0] _seach_blockx_409_map_block;
  wire [9:0] _seach_blockx_409_now;
  wire [9:0] _seach_blockx_409_start;
  wire [9:0] _seach_blockx_409_goal;
  wire [9:0] _seach_blockx_409_data_out;
  wire _seach_blockx_409_in_do;
  wire _seach_blockx_409_p_reset;
  wire _seach_blockx_409_m_clock;
  wire [9:0] _seach_blockx_408_map_block;
  wire [9:0] _seach_blockx_408_now;
  wire [9:0] _seach_blockx_408_start;
  wire [9:0] _seach_blockx_408_goal;
  wire [9:0] _seach_blockx_408_data_out;
  wire _seach_blockx_408_in_do;
  wire _seach_blockx_408_p_reset;
  wire _seach_blockx_408_m_clock;
  wire [9:0] _seach_blockx_407_map_block;
  wire [9:0] _seach_blockx_407_now;
  wire [9:0] _seach_blockx_407_start;
  wire [9:0] _seach_blockx_407_goal;
  wire [9:0] _seach_blockx_407_data_out;
  wire _seach_blockx_407_in_do;
  wire _seach_blockx_407_p_reset;
  wire _seach_blockx_407_m_clock;
  wire [9:0] _seach_blockx_406_map_block;
  wire [9:0] _seach_blockx_406_now;
  wire [9:0] _seach_blockx_406_start;
  wire [9:0] _seach_blockx_406_goal;
  wire [9:0] _seach_blockx_406_data_out;
  wire _seach_blockx_406_in_do;
  wire _seach_blockx_406_p_reset;
  wire _seach_blockx_406_m_clock;
  wire [9:0] _seach_blockx_405_map_block;
  wire [9:0] _seach_blockx_405_now;
  wire [9:0] _seach_blockx_405_start;
  wire [9:0] _seach_blockx_405_goal;
  wire [9:0] _seach_blockx_405_data_out;
  wire _seach_blockx_405_in_do;
  wire _seach_blockx_405_p_reset;
  wire _seach_blockx_405_m_clock;
  wire [9:0] _seach_blockx_404_map_block;
  wire [9:0] _seach_blockx_404_now;
  wire [9:0] _seach_blockx_404_start;
  wire [9:0] _seach_blockx_404_goal;
  wire [9:0] _seach_blockx_404_data_out;
  wire _seach_blockx_404_in_do;
  wire _seach_blockx_404_p_reset;
  wire _seach_blockx_404_m_clock;
  wire [9:0] _seach_blockx_403_map_block;
  wire [9:0] _seach_blockx_403_now;
  wire [9:0] _seach_blockx_403_start;
  wire [9:0] _seach_blockx_403_goal;
  wire [9:0] _seach_blockx_403_data_out;
  wire _seach_blockx_403_in_do;
  wire _seach_blockx_403_p_reset;
  wire _seach_blockx_403_m_clock;
  wire [9:0] _seach_blockx_402_map_block;
  wire [9:0] _seach_blockx_402_now;
  wire [9:0] _seach_blockx_402_start;
  wire [9:0] _seach_blockx_402_goal;
  wire [9:0] _seach_blockx_402_data_out;
  wire _seach_blockx_402_in_do;
  wire _seach_blockx_402_p_reset;
  wire _seach_blockx_402_m_clock;
  wire [9:0] _seach_blockx_401_map_block;
  wire [9:0] _seach_blockx_401_now;
  wire [9:0] _seach_blockx_401_start;
  wire [9:0] _seach_blockx_401_goal;
  wire [9:0] _seach_blockx_401_data_out;
  wire _seach_blockx_401_in_do;
  wire _seach_blockx_401_p_reset;
  wire _seach_blockx_401_m_clock;
  wire [9:0] _seach_blockx_400_map_block;
  wire [9:0] _seach_blockx_400_now;
  wire [9:0] _seach_blockx_400_start;
  wire [9:0] _seach_blockx_400_goal;
  wire [9:0] _seach_blockx_400_data_out;
  wire _seach_blockx_400_in_do;
  wire _seach_blockx_400_p_reset;
  wire _seach_blockx_400_m_clock;
  wire [9:0] _seach_blockx_399_map_block;
  wire [9:0] _seach_blockx_399_now;
  wire [9:0] _seach_blockx_399_start;
  wire [9:0] _seach_blockx_399_goal;
  wire [9:0] _seach_blockx_399_data_out;
  wire _seach_blockx_399_in_do;
  wire _seach_blockx_399_p_reset;
  wire _seach_blockx_399_m_clock;
  wire [9:0] _seach_blockx_398_map_block;
  wire [9:0] _seach_blockx_398_now;
  wire [9:0] _seach_blockx_398_start;
  wire [9:0] _seach_blockx_398_goal;
  wire [9:0] _seach_blockx_398_data_out;
  wire _seach_blockx_398_in_do;
  wire _seach_blockx_398_p_reset;
  wire _seach_blockx_398_m_clock;
  wire [9:0] _seach_blockx_397_map_block;
  wire [9:0] _seach_blockx_397_now;
  wire [9:0] _seach_blockx_397_start;
  wire [9:0] _seach_blockx_397_goal;
  wire [9:0] _seach_blockx_397_data_out;
  wire _seach_blockx_397_in_do;
  wire _seach_blockx_397_p_reset;
  wire _seach_blockx_397_m_clock;
  wire [9:0] _seach_blockx_396_map_block;
  wire [9:0] _seach_blockx_396_now;
  wire [9:0] _seach_blockx_396_start;
  wire [9:0] _seach_blockx_396_goal;
  wire [9:0] _seach_blockx_396_data_out;
  wire _seach_blockx_396_in_do;
  wire _seach_blockx_396_p_reset;
  wire _seach_blockx_396_m_clock;
  wire [9:0] _seach_blockx_395_map_block;
  wire [9:0] _seach_blockx_395_now;
  wire [9:0] _seach_blockx_395_start;
  wire [9:0] _seach_blockx_395_goal;
  wire [9:0] _seach_blockx_395_data_out;
  wire _seach_blockx_395_in_do;
  wire _seach_blockx_395_p_reset;
  wire _seach_blockx_395_m_clock;
  wire [9:0] _seach_blockx_394_map_block;
  wire [9:0] _seach_blockx_394_now;
  wire [9:0] _seach_blockx_394_start;
  wire [9:0] _seach_blockx_394_goal;
  wire [9:0] _seach_blockx_394_data_out;
  wire _seach_blockx_394_in_do;
  wire _seach_blockx_394_p_reset;
  wire _seach_blockx_394_m_clock;
  wire [9:0] _seach_blockx_393_map_block;
  wire [9:0] _seach_blockx_393_now;
  wire [9:0] _seach_blockx_393_start;
  wire [9:0] _seach_blockx_393_goal;
  wire [9:0] _seach_blockx_393_data_out;
  wire _seach_blockx_393_in_do;
  wire _seach_blockx_393_p_reset;
  wire _seach_blockx_393_m_clock;
  wire [9:0] _seach_blockx_392_map_block;
  wire [9:0] _seach_blockx_392_now;
  wire [9:0] _seach_blockx_392_start;
  wire [9:0] _seach_blockx_392_goal;
  wire [9:0] _seach_blockx_392_data_out;
  wire _seach_blockx_392_in_do;
  wire _seach_blockx_392_p_reset;
  wire _seach_blockx_392_m_clock;
  wire [9:0] _seach_blockx_391_map_block;
  wire [9:0] _seach_blockx_391_now;
  wire [9:0] _seach_blockx_391_start;
  wire [9:0] _seach_blockx_391_goal;
  wire [9:0] _seach_blockx_391_data_out;
  wire _seach_blockx_391_in_do;
  wire _seach_blockx_391_p_reset;
  wire _seach_blockx_391_m_clock;
  wire [9:0] _seach_blockx_390_map_block;
  wire [9:0] _seach_blockx_390_now;
  wire [9:0] _seach_blockx_390_start;
  wire [9:0] _seach_blockx_390_goal;
  wire [9:0] _seach_blockx_390_data_out;
  wire _seach_blockx_390_in_do;
  wire _seach_blockx_390_p_reset;
  wire _seach_blockx_390_m_clock;
  wire [9:0] _seach_blockx_389_map_block;
  wire [9:0] _seach_blockx_389_now;
  wire [9:0] _seach_blockx_389_start;
  wire [9:0] _seach_blockx_389_goal;
  wire [9:0] _seach_blockx_389_data_out;
  wire _seach_blockx_389_in_do;
  wire _seach_blockx_389_p_reset;
  wire _seach_blockx_389_m_clock;
  wire [9:0] _seach_blockx_388_map_block;
  wire [9:0] _seach_blockx_388_now;
  wire [9:0] _seach_blockx_388_start;
  wire [9:0] _seach_blockx_388_goal;
  wire [9:0] _seach_blockx_388_data_out;
  wire _seach_blockx_388_in_do;
  wire _seach_blockx_388_p_reset;
  wire _seach_blockx_388_m_clock;
  wire [9:0] _seach_blockx_387_map_block;
  wire [9:0] _seach_blockx_387_now;
  wire [9:0] _seach_blockx_387_start;
  wire [9:0] _seach_blockx_387_goal;
  wire [9:0] _seach_blockx_387_data_out;
  wire _seach_blockx_387_in_do;
  wire _seach_blockx_387_p_reset;
  wire _seach_blockx_387_m_clock;
  wire [9:0] _seach_blockx_386_map_block;
  wire [9:0] _seach_blockx_386_now;
  wire [9:0] _seach_blockx_386_start;
  wire [9:0] _seach_blockx_386_goal;
  wire [9:0] _seach_blockx_386_data_out;
  wire _seach_blockx_386_in_do;
  wire _seach_blockx_386_p_reset;
  wire _seach_blockx_386_m_clock;
  wire [9:0] _seach_blockx_385_map_block;
  wire [9:0] _seach_blockx_385_now;
  wire [9:0] _seach_blockx_385_start;
  wire [9:0] _seach_blockx_385_goal;
  wire [9:0] _seach_blockx_385_data_out;
  wire _seach_blockx_385_in_do;
  wire _seach_blockx_385_p_reset;
  wire _seach_blockx_385_m_clock;
  wire [9:0] _seach_blockx_384_map_block;
  wire [9:0] _seach_blockx_384_now;
  wire [9:0] _seach_blockx_384_start;
  wire [9:0] _seach_blockx_384_goal;
  wire [9:0] _seach_blockx_384_data_out;
  wire _seach_blockx_384_in_do;
  wire _seach_blockx_384_p_reset;
  wire _seach_blockx_384_m_clock;
  wire [9:0] _seach_blockx_383_map_block;
  wire [9:0] _seach_blockx_383_now;
  wire [9:0] _seach_blockx_383_start;
  wire [9:0] _seach_blockx_383_goal;
  wire [9:0] _seach_blockx_383_data_out;
  wire _seach_blockx_383_in_do;
  wire _seach_blockx_383_p_reset;
  wire _seach_blockx_383_m_clock;
  wire [9:0] _seach_blockx_382_map_block;
  wire [9:0] _seach_blockx_382_now;
  wire [9:0] _seach_blockx_382_start;
  wire [9:0] _seach_blockx_382_goal;
  wire [9:0] _seach_blockx_382_data_out;
  wire _seach_blockx_382_in_do;
  wire _seach_blockx_382_p_reset;
  wire _seach_blockx_382_m_clock;
  wire [9:0] _seach_blockx_381_map_block;
  wire [9:0] _seach_blockx_381_now;
  wire [9:0] _seach_blockx_381_start;
  wire [9:0] _seach_blockx_381_goal;
  wire [9:0] _seach_blockx_381_data_out;
  wire _seach_blockx_381_in_do;
  wire _seach_blockx_381_p_reset;
  wire _seach_blockx_381_m_clock;
  wire [9:0] _seach_blockx_380_map_block;
  wire [9:0] _seach_blockx_380_now;
  wire [9:0] _seach_blockx_380_start;
  wire [9:0] _seach_blockx_380_goal;
  wire [9:0] _seach_blockx_380_data_out;
  wire _seach_blockx_380_in_do;
  wire _seach_blockx_380_p_reset;
  wire _seach_blockx_380_m_clock;
  wire [9:0] _seach_blockx_379_map_block;
  wire [9:0] _seach_blockx_379_now;
  wire [9:0] _seach_blockx_379_start;
  wire [9:0] _seach_blockx_379_goal;
  wire [9:0] _seach_blockx_379_data_out;
  wire _seach_blockx_379_in_do;
  wire _seach_blockx_379_p_reset;
  wire _seach_blockx_379_m_clock;
  wire [9:0] _seach_blockx_378_map_block;
  wire [9:0] _seach_blockx_378_now;
  wire [9:0] _seach_blockx_378_start;
  wire [9:0] _seach_blockx_378_goal;
  wire [9:0] _seach_blockx_378_data_out;
  wire _seach_blockx_378_in_do;
  wire _seach_blockx_378_p_reset;
  wire _seach_blockx_378_m_clock;
  wire [9:0] _seach_blockx_377_map_block;
  wire [9:0] _seach_blockx_377_now;
  wire [9:0] _seach_blockx_377_start;
  wire [9:0] _seach_blockx_377_goal;
  wire [9:0] _seach_blockx_377_data_out;
  wire _seach_blockx_377_in_do;
  wire _seach_blockx_377_p_reset;
  wire _seach_blockx_377_m_clock;
  wire [9:0] _seach_blockx_376_map_block;
  wire [9:0] _seach_blockx_376_now;
  wire [9:0] _seach_blockx_376_start;
  wire [9:0] _seach_blockx_376_goal;
  wire [9:0] _seach_blockx_376_data_out;
  wire _seach_blockx_376_in_do;
  wire _seach_blockx_376_p_reset;
  wire _seach_blockx_376_m_clock;
  wire [9:0] _seach_blockx_375_map_block;
  wire [9:0] _seach_blockx_375_now;
  wire [9:0] _seach_blockx_375_start;
  wire [9:0] _seach_blockx_375_goal;
  wire [9:0] _seach_blockx_375_data_out;
  wire _seach_blockx_375_in_do;
  wire _seach_blockx_375_p_reset;
  wire _seach_blockx_375_m_clock;
  wire [9:0] _seach_blockx_374_map_block;
  wire [9:0] _seach_blockx_374_now;
  wire [9:0] _seach_blockx_374_start;
  wire [9:0] _seach_blockx_374_goal;
  wire [9:0] _seach_blockx_374_data_out;
  wire _seach_blockx_374_in_do;
  wire _seach_blockx_374_p_reset;
  wire _seach_blockx_374_m_clock;
  wire [9:0] _seach_blockx_373_map_block;
  wire [9:0] _seach_blockx_373_now;
  wire [9:0] _seach_blockx_373_start;
  wire [9:0] _seach_blockx_373_goal;
  wire [9:0] _seach_blockx_373_data_out;
  wire _seach_blockx_373_in_do;
  wire _seach_blockx_373_p_reset;
  wire _seach_blockx_373_m_clock;
  wire [9:0] _seach_blockx_372_map_block;
  wire [9:0] _seach_blockx_372_now;
  wire [9:0] _seach_blockx_372_start;
  wire [9:0] _seach_blockx_372_goal;
  wire [9:0] _seach_blockx_372_data_out;
  wire _seach_blockx_372_in_do;
  wire _seach_blockx_372_p_reset;
  wire _seach_blockx_372_m_clock;
  wire [9:0] _seach_blockx_371_map_block;
  wire [9:0] _seach_blockx_371_now;
  wire [9:0] _seach_blockx_371_start;
  wire [9:0] _seach_blockx_371_goal;
  wire [9:0] _seach_blockx_371_data_out;
  wire _seach_blockx_371_in_do;
  wire _seach_blockx_371_p_reset;
  wire _seach_blockx_371_m_clock;
  wire [9:0] _seach_blockx_370_map_block;
  wire [9:0] _seach_blockx_370_now;
  wire [9:0] _seach_blockx_370_start;
  wire [9:0] _seach_blockx_370_goal;
  wire [9:0] _seach_blockx_370_data_out;
  wire _seach_blockx_370_in_do;
  wire _seach_blockx_370_p_reset;
  wire _seach_blockx_370_m_clock;
  wire [9:0] _seach_blockx_369_map_block;
  wire [9:0] _seach_blockx_369_now;
  wire [9:0] _seach_blockx_369_start;
  wire [9:0] _seach_blockx_369_goal;
  wire [9:0] _seach_blockx_369_data_out;
  wire _seach_blockx_369_in_do;
  wire _seach_blockx_369_p_reset;
  wire _seach_blockx_369_m_clock;
  wire [9:0] _seach_blockx_368_map_block;
  wire [9:0] _seach_blockx_368_now;
  wire [9:0] _seach_blockx_368_start;
  wire [9:0] _seach_blockx_368_goal;
  wire [9:0] _seach_blockx_368_data_out;
  wire _seach_blockx_368_in_do;
  wire _seach_blockx_368_p_reset;
  wire _seach_blockx_368_m_clock;
  wire [9:0] _seach_blockx_367_map_block;
  wire [9:0] _seach_blockx_367_now;
  wire [9:0] _seach_blockx_367_start;
  wire [9:0] _seach_blockx_367_goal;
  wire [9:0] _seach_blockx_367_data_out;
  wire _seach_blockx_367_in_do;
  wire _seach_blockx_367_p_reset;
  wire _seach_blockx_367_m_clock;
  wire [9:0] _seach_blockx_366_map_block;
  wire [9:0] _seach_blockx_366_now;
  wire [9:0] _seach_blockx_366_start;
  wire [9:0] _seach_blockx_366_goal;
  wire [9:0] _seach_blockx_366_data_out;
  wire _seach_blockx_366_in_do;
  wire _seach_blockx_366_p_reset;
  wire _seach_blockx_366_m_clock;
  wire [9:0] _seach_blockx_365_map_block;
  wire [9:0] _seach_blockx_365_now;
  wire [9:0] _seach_blockx_365_start;
  wire [9:0] _seach_blockx_365_goal;
  wire [9:0] _seach_blockx_365_data_out;
  wire _seach_blockx_365_in_do;
  wire _seach_blockx_365_p_reset;
  wire _seach_blockx_365_m_clock;
  wire [9:0] _seach_blockx_364_map_block;
  wire [9:0] _seach_blockx_364_now;
  wire [9:0] _seach_blockx_364_start;
  wire [9:0] _seach_blockx_364_goal;
  wire [9:0] _seach_blockx_364_data_out;
  wire _seach_blockx_364_in_do;
  wire _seach_blockx_364_p_reset;
  wire _seach_blockx_364_m_clock;
  wire [9:0] _seach_blockx_363_map_block;
  wire [9:0] _seach_blockx_363_now;
  wire [9:0] _seach_blockx_363_start;
  wire [9:0] _seach_blockx_363_goal;
  wire [9:0] _seach_blockx_363_data_out;
  wire _seach_blockx_363_in_do;
  wire _seach_blockx_363_p_reset;
  wire _seach_blockx_363_m_clock;
  wire [9:0] _seach_blockx_362_map_block;
  wire [9:0] _seach_blockx_362_now;
  wire [9:0] _seach_blockx_362_start;
  wire [9:0] _seach_blockx_362_goal;
  wire [9:0] _seach_blockx_362_data_out;
  wire _seach_blockx_362_in_do;
  wire _seach_blockx_362_p_reset;
  wire _seach_blockx_362_m_clock;
  wire [9:0] _seach_blockx_361_map_block;
  wire [9:0] _seach_blockx_361_now;
  wire [9:0] _seach_blockx_361_start;
  wire [9:0] _seach_blockx_361_goal;
  wire [9:0] _seach_blockx_361_data_out;
  wire _seach_blockx_361_in_do;
  wire _seach_blockx_361_p_reset;
  wire _seach_blockx_361_m_clock;
  wire [9:0] _seach_blockx_360_map_block;
  wire [9:0] _seach_blockx_360_now;
  wire [9:0] _seach_blockx_360_start;
  wire [9:0] _seach_blockx_360_goal;
  wire [9:0] _seach_blockx_360_data_out;
  wire _seach_blockx_360_in_do;
  wire _seach_blockx_360_p_reset;
  wire _seach_blockx_360_m_clock;
  wire [9:0] _seach_blockx_359_map_block;
  wire [9:0] _seach_blockx_359_now;
  wire [9:0] _seach_blockx_359_start;
  wire [9:0] _seach_blockx_359_goal;
  wire [9:0] _seach_blockx_359_data_out;
  wire _seach_blockx_359_in_do;
  wire _seach_blockx_359_p_reset;
  wire _seach_blockx_359_m_clock;
  wire [9:0] _seach_blockx_358_map_block;
  wire [9:0] _seach_blockx_358_now;
  wire [9:0] _seach_blockx_358_start;
  wire [9:0] _seach_blockx_358_goal;
  wire [9:0] _seach_blockx_358_data_out;
  wire _seach_blockx_358_in_do;
  wire _seach_blockx_358_p_reset;
  wire _seach_blockx_358_m_clock;
  wire [9:0] _seach_blockx_357_map_block;
  wire [9:0] _seach_blockx_357_now;
  wire [9:0] _seach_blockx_357_start;
  wire [9:0] _seach_blockx_357_goal;
  wire [9:0] _seach_blockx_357_data_out;
  wire _seach_blockx_357_in_do;
  wire _seach_blockx_357_p_reset;
  wire _seach_blockx_357_m_clock;
  wire [9:0] _seach_blockx_356_map_block;
  wire [9:0] _seach_blockx_356_now;
  wire [9:0] _seach_blockx_356_start;
  wire [9:0] _seach_blockx_356_goal;
  wire [9:0] _seach_blockx_356_data_out;
  wire _seach_blockx_356_in_do;
  wire _seach_blockx_356_p_reset;
  wire _seach_blockx_356_m_clock;
  wire [9:0] _seach_blockx_355_map_block;
  wire [9:0] _seach_blockx_355_now;
  wire [9:0] _seach_blockx_355_start;
  wire [9:0] _seach_blockx_355_goal;
  wire [9:0] _seach_blockx_355_data_out;
  wire _seach_blockx_355_in_do;
  wire _seach_blockx_355_p_reset;
  wire _seach_blockx_355_m_clock;
  wire [9:0] _seach_blockx_354_map_block;
  wire [9:0] _seach_blockx_354_now;
  wire [9:0] _seach_blockx_354_start;
  wire [9:0] _seach_blockx_354_goal;
  wire [9:0] _seach_blockx_354_data_out;
  wire _seach_blockx_354_in_do;
  wire _seach_blockx_354_p_reset;
  wire _seach_blockx_354_m_clock;
  wire [9:0] _seach_blockx_353_map_block;
  wire [9:0] _seach_blockx_353_now;
  wire [9:0] _seach_blockx_353_start;
  wire [9:0] _seach_blockx_353_goal;
  wire [9:0] _seach_blockx_353_data_out;
  wire _seach_blockx_353_in_do;
  wire _seach_blockx_353_p_reset;
  wire _seach_blockx_353_m_clock;
  wire [9:0] _seach_blockx_352_map_block;
  wire [9:0] _seach_blockx_352_now;
  wire [9:0] _seach_blockx_352_start;
  wire [9:0] _seach_blockx_352_goal;
  wire [9:0] _seach_blockx_352_data_out;
  wire _seach_blockx_352_in_do;
  wire _seach_blockx_352_p_reset;
  wire _seach_blockx_352_m_clock;
  wire [9:0] _seach_blockx_351_map_block;
  wire [9:0] _seach_blockx_351_now;
  wire [9:0] _seach_blockx_351_start;
  wire [9:0] _seach_blockx_351_goal;
  wire [9:0] _seach_blockx_351_data_out;
  wire _seach_blockx_351_in_do;
  wire _seach_blockx_351_p_reset;
  wire _seach_blockx_351_m_clock;
  wire [9:0] _seach_blockx_350_map_block;
  wire [9:0] _seach_blockx_350_now;
  wire [9:0] _seach_blockx_350_start;
  wire [9:0] _seach_blockx_350_goal;
  wire [9:0] _seach_blockx_350_data_out;
  wire _seach_blockx_350_in_do;
  wire _seach_blockx_350_p_reset;
  wire _seach_blockx_350_m_clock;
  wire [9:0] _seach_blockx_349_map_block;
  wire [9:0] _seach_blockx_349_now;
  wire [9:0] _seach_blockx_349_start;
  wire [9:0] _seach_blockx_349_goal;
  wire [9:0] _seach_blockx_349_data_out;
  wire _seach_blockx_349_in_do;
  wire _seach_blockx_349_p_reset;
  wire _seach_blockx_349_m_clock;
  wire [9:0] _seach_blockx_348_map_block;
  wire [9:0] _seach_blockx_348_now;
  wire [9:0] _seach_blockx_348_start;
  wire [9:0] _seach_blockx_348_goal;
  wire [9:0] _seach_blockx_348_data_out;
  wire _seach_blockx_348_in_do;
  wire _seach_blockx_348_p_reset;
  wire _seach_blockx_348_m_clock;
  wire [9:0] _seach_blockx_347_map_block;
  wire [9:0] _seach_blockx_347_now;
  wire [9:0] _seach_blockx_347_start;
  wire [9:0] _seach_blockx_347_goal;
  wire [9:0] _seach_blockx_347_data_out;
  wire _seach_blockx_347_in_do;
  wire _seach_blockx_347_p_reset;
  wire _seach_blockx_347_m_clock;
  wire [9:0] _seach_blockx_346_map_block;
  wire [9:0] _seach_blockx_346_now;
  wire [9:0] _seach_blockx_346_start;
  wire [9:0] _seach_blockx_346_goal;
  wire [9:0] _seach_blockx_346_data_out;
  wire _seach_blockx_346_in_do;
  wire _seach_blockx_346_p_reset;
  wire _seach_blockx_346_m_clock;
  wire [9:0] _seach_blockx_345_map_block;
  wire [9:0] _seach_blockx_345_now;
  wire [9:0] _seach_blockx_345_start;
  wire [9:0] _seach_blockx_345_goal;
  wire [9:0] _seach_blockx_345_data_out;
  wire _seach_blockx_345_in_do;
  wire _seach_blockx_345_p_reset;
  wire _seach_blockx_345_m_clock;
  wire [9:0] _seach_blockx_344_map_block;
  wire [9:0] _seach_blockx_344_now;
  wire [9:0] _seach_blockx_344_start;
  wire [9:0] _seach_blockx_344_goal;
  wire [9:0] _seach_blockx_344_data_out;
  wire _seach_blockx_344_in_do;
  wire _seach_blockx_344_p_reset;
  wire _seach_blockx_344_m_clock;
  wire [9:0] _seach_blockx_343_map_block;
  wire [9:0] _seach_blockx_343_now;
  wire [9:0] _seach_blockx_343_start;
  wire [9:0] _seach_blockx_343_goal;
  wire [9:0] _seach_blockx_343_data_out;
  wire _seach_blockx_343_in_do;
  wire _seach_blockx_343_p_reset;
  wire _seach_blockx_343_m_clock;
  wire [9:0] _seach_blockx_342_map_block;
  wire [9:0] _seach_blockx_342_now;
  wire [9:0] _seach_blockx_342_start;
  wire [9:0] _seach_blockx_342_goal;
  wire [9:0] _seach_blockx_342_data_out;
  wire _seach_blockx_342_in_do;
  wire _seach_blockx_342_p_reset;
  wire _seach_blockx_342_m_clock;
  wire [9:0] _seach_blockx_341_map_block;
  wire [9:0] _seach_blockx_341_now;
  wire [9:0] _seach_blockx_341_start;
  wire [9:0] _seach_blockx_341_goal;
  wire [9:0] _seach_blockx_341_data_out;
  wire _seach_blockx_341_in_do;
  wire _seach_blockx_341_p_reset;
  wire _seach_blockx_341_m_clock;
  wire [9:0] _seach_blockx_340_map_block;
  wire [9:0] _seach_blockx_340_now;
  wire [9:0] _seach_blockx_340_start;
  wire [9:0] _seach_blockx_340_goal;
  wire [9:0] _seach_blockx_340_data_out;
  wire _seach_blockx_340_in_do;
  wire _seach_blockx_340_p_reset;
  wire _seach_blockx_340_m_clock;
  wire [9:0] _seach_blockx_339_map_block;
  wire [9:0] _seach_blockx_339_now;
  wire [9:0] _seach_blockx_339_start;
  wire [9:0] _seach_blockx_339_goal;
  wire [9:0] _seach_blockx_339_data_out;
  wire _seach_blockx_339_in_do;
  wire _seach_blockx_339_p_reset;
  wire _seach_blockx_339_m_clock;
  wire [9:0] _seach_blockx_338_map_block;
  wire [9:0] _seach_blockx_338_now;
  wire [9:0] _seach_blockx_338_start;
  wire [9:0] _seach_blockx_338_goal;
  wire [9:0] _seach_blockx_338_data_out;
  wire _seach_blockx_338_in_do;
  wire _seach_blockx_338_p_reset;
  wire _seach_blockx_338_m_clock;
  wire [9:0] _seach_blockx_337_map_block;
  wire [9:0] _seach_blockx_337_now;
  wire [9:0] _seach_blockx_337_start;
  wire [9:0] _seach_blockx_337_goal;
  wire [9:0] _seach_blockx_337_data_out;
  wire _seach_blockx_337_in_do;
  wire _seach_blockx_337_p_reset;
  wire _seach_blockx_337_m_clock;
  wire [9:0] _seach_blockx_336_map_block;
  wire [9:0] _seach_blockx_336_now;
  wire [9:0] _seach_blockx_336_start;
  wire [9:0] _seach_blockx_336_goal;
  wire [9:0] _seach_blockx_336_data_out;
  wire _seach_blockx_336_in_do;
  wire _seach_blockx_336_p_reset;
  wire _seach_blockx_336_m_clock;
  wire [9:0] _seach_blockx_335_map_block;
  wire [9:0] _seach_blockx_335_now;
  wire [9:0] _seach_blockx_335_start;
  wire [9:0] _seach_blockx_335_goal;
  wire [9:0] _seach_blockx_335_data_out;
  wire _seach_blockx_335_in_do;
  wire _seach_blockx_335_p_reset;
  wire _seach_blockx_335_m_clock;
  wire [9:0] _seach_blockx_334_map_block;
  wire [9:0] _seach_blockx_334_now;
  wire [9:0] _seach_blockx_334_start;
  wire [9:0] _seach_blockx_334_goal;
  wire [9:0] _seach_blockx_334_data_out;
  wire _seach_blockx_334_in_do;
  wire _seach_blockx_334_p_reset;
  wire _seach_blockx_334_m_clock;
  wire [9:0] _seach_blockx_333_map_block;
  wire [9:0] _seach_blockx_333_now;
  wire [9:0] _seach_blockx_333_start;
  wire [9:0] _seach_blockx_333_goal;
  wire [9:0] _seach_blockx_333_data_out;
  wire _seach_blockx_333_in_do;
  wire _seach_blockx_333_p_reset;
  wire _seach_blockx_333_m_clock;
  wire [9:0] _seach_blockx_332_map_block;
  wire [9:0] _seach_blockx_332_now;
  wire [9:0] _seach_blockx_332_start;
  wire [9:0] _seach_blockx_332_goal;
  wire [9:0] _seach_blockx_332_data_out;
  wire _seach_blockx_332_in_do;
  wire _seach_blockx_332_p_reset;
  wire _seach_blockx_332_m_clock;
  wire [9:0] _seach_blockx_331_map_block;
  wire [9:0] _seach_blockx_331_now;
  wire [9:0] _seach_blockx_331_start;
  wire [9:0] _seach_blockx_331_goal;
  wire [9:0] _seach_blockx_331_data_out;
  wire _seach_blockx_331_in_do;
  wire _seach_blockx_331_p_reset;
  wire _seach_blockx_331_m_clock;
  wire [9:0] _seach_blockx_330_map_block;
  wire [9:0] _seach_blockx_330_now;
  wire [9:0] _seach_blockx_330_start;
  wire [9:0] _seach_blockx_330_goal;
  wire [9:0] _seach_blockx_330_data_out;
  wire _seach_blockx_330_in_do;
  wire _seach_blockx_330_p_reset;
  wire _seach_blockx_330_m_clock;
  wire [9:0] _seach_blockx_329_map_block;
  wire [9:0] _seach_blockx_329_now;
  wire [9:0] _seach_blockx_329_start;
  wire [9:0] _seach_blockx_329_goal;
  wire [9:0] _seach_blockx_329_data_out;
  wire _seach_blockx_329_in_do;
  wire _seach_blockx_329_p_reset;
  wire _seach_blockx_329_m_clock;
  wire [9:0] _seach_blockx_328_map_block;
  wire [9:0] _seach_blockx_328_now;
  wire [9:0] _seach_blockx_328_start;
  wire [9:0] _seach_blockx_328_goal;
  wire [9:0] _seach_blockx_328_data_out;
  wire _seach_blockx_328_in_do;
  wire _seach_blockx_328_p_reset;
  wire _seach_blockx_328_m_clock;
  wire [9:0] _seach_blockx_327_map_block;
  wire [9:0] _seach_blockx_327_now;
  wire [9:0] _seach_blockx_327_start;
  wire [9:0] _seach_blockx_327_goal;
  wire [9:0] _seach_blockx_327_data_out;
  wire _seach_blockx_327_in_do;
  wire _seach_blockx_327_p_reset;
  wire _seach_blockx_327_m_clock;
  wire [9:0] _seach_blockx_326_map_block;
  wire [9:0] _seach_blockx_326_now;
  wire [9:0] _seach_blockx_326_start;
  wire [9:0] _seach_blockx_326_goal;
  wire [9:0] _seach_blockx_326_data_out;
  wire _seach_blockx_326_in_do;
  wire _seach_blockx_326_p_reset;
  wire _seach_blockx_326_m_clock;
  wire [9:0] _seach_blockx_325_map_block;
  wire [9:0] _seach_blockx_325_now;
  wire [9:0] _seach_blockx_325_start;
  wire [9:0] _seach_blockx_325_goal;
  wire [9:0] _seach_blockx_325_data_out;
  wire _seach_blockx_325_in_do;
  wire _seach_blockx_325_p_reset;
  wire _seach_blockx_325_m_clock;
  wire [9:0] _seach_blockx_324_map_block;
  wire [9:0] _seach_blockx_324_now;
  wire [9:0] _seach_blockx_324_start;
  wire [9:0] _seach_blockx_324_goal;
  wire [9:0] _seach_blockx_324_data_out;
  wire _seach_blockx_324_in_do;
  wire _seach_blockx_324_p_reset;
  wire _seach_blockx_324_m_clock;
  wire [9:0] _seach_blockx_323_map_block;
  wire [9:0] _seach_blockx_323_now;
  wire [9:0] _seach_blockx_323_start;
  wire [9:0] _seach_blockx_323_goal;
  wire [9:0] _seach_blockx_323_data_out;
  wire _seach_blockx_323_in_do;
  wire _seach_blockx_323_p_reset;
  wire _seach_blockx_323_m_clock;
  wire [9:0] _seach_blockx_322_map_block;
  wire [9:0] _seach_blockx_322_now;
  wire [9:0] _seach_blockx_322_start;
  wire [9:0] _seach_blockx_322_goal;
  wire [9:0] _seach_blockx_322_data_out;
  wire _seach_blockx_322_in_do;
  wire _seach_blockx_322_p_reset;
  wire _seach_blockx_322_m_clock;
  wire [9:0] _seach_blockx_321_map_block;
  wire [9:0] _seach_blockx_321_now;
  wire [9:0] _seach_blockx_321_start;
  wire [9:0] _seach_blockx_321_goal;
  wire [9:0] _seach_blockx_321_data_out;
  wire _seach_blockx_321_in_do;
  wire _seach_blockx_321_p_reset;
  wire _seach_blockx_321_m_clock;
  wire [9:0] _seach_blockx_320_map_block;
  wire [9:0] _seach_blockx_320_now;
  wire [9:0] _seach_blockx_320_start;
  wire [9:0] _seach_blockx_320_goal;
  wire [9:0] _seach_blockx_320_data_out;
  wire _seach_blockx_320_in_do;
  wire _seach_blockx_320_p_reset;
  wire _seach_blockx_320_m_clock;
  wire [9:0] _seach_blockx_319_map_block;
  wire [9:0] _seach_blockx_319_now;
  wire [9:0] _seach_blockx_319_start;
  wire [9:0] _seach_blockx_319_goal;
  wire [9:0] _seach_blockx_319_data_out;
  wire _seach_blockx_319_in_do;
  wire _seach_blockx_319_p_reset;
  wire _seach_blockx_319_m_clock;
  wire [9:0] _seach_blockx_318_map_block;
  wire [9:0] _seach_blockx_318_now;
  wire [9:0] _seach_blockx_318_start;
  wire [9:0] _seach_blockx_318_goal;
  wire [9:0] _seach_blockx_318_data_out;
  wire _seach_blockx_318_in_do;
  wire _seach_blockx_318_p_reset;
  wire _seach_blockx_318_m_clock;
  wire [9:0] _seach_blockx_317_map_block;
  wire [9:0] _seach_blockx_317_now;
  wire [9:0] _seach_blockx_317_start;
  wire [9:0] _seach_blockx_317_goal;
  wire [9:0] _seach_blockx_317_data_out;
  wire _seach_blockx_317_in_do;
  wire _seach_blockx_317_p_reset;
  wire _seach_blockx_317_m_clock;
  wire [9:0] _seach_blockx_316_map_block;
  wire [9:0] _seach_blockx_316_now;
  wire [9:0] _seach_blockx_316_start;
  wire [9:0] _seach_blockx_316_goal;
  wire [9:0] _seach_blockx_316_data_out;
  wire _seach_blockx_316_in_do;
  wire _seach_blockx_316_p_reset;
  wire _seach_blockx_316_m_clock;
  wire [9:0] _seach_blockx_315_map_block;
  wire [9:0] _seach_blockx_315_now;
  wire [9:0] _seach_blockx_315_start;
  wire [9:0] _seach_blockx_315_goal;
  wire [9:0] _seach_blockx_315_data_out;
  wire _seach_blockx_315_in_do;
  wire _seach_blockx_315_p_reset;
  wire _seach_blockx_315_m_clock;
  wire [9:0] _seach_blockx_314_map_block;
  wire [9:0] _seach_blockx_314_now;
  wire [9:0] _seach_blockx_314_start;
  wire [9:0] _seach_blockx_314_goal;
  wire [9:0] _seach_blockx_314_data_out;
  wire _seach_blockx_314_in_do;
  wire _seach_blockx_314_p_reset;
  wire _seach_blockx_314_m_clock;
  wire [9:0] _seach_blockx_313_map_block;
  wire [9:0] _seach_blockx_313_now;
  wire [9:0] _seach_blockx_313_start;
  wire [9:0] _seach_blockx_313_goal;
  wire [9:0] _seach_blockx_313_data_out;
  wire _seach_blockx_313_in_do;
  wire _seach_blockx_313_p_reset;
  wire _seach_blockx_313_m_clock;
  wire [9:0] _seach_blockx_312_map_block;
  wire [9:0] _seach_blockx_312_now;
  wire [9:0] _seach_blockx_312_start;
  wire [9:0] _seach_blockx_312_goal;
  wire [9:0] _seach_blockx_312_data_out;
  wire _seach_blockx_312_in_do;
  wire _seach_blockx_312_p_reset;
  wire _seach_blockx_312_m_clock;
  wire [9:0] _seach_blockx_311_map_block;
  wire [9:0] _seach_blockx_311_now;
  wire [9:0] _seach_blockx_311_start;
  wire [9:0] _seach_blockx_311_goal;
  wire [9:0] _seach_blockx_311_data_out;
  wire _seach_blockx_311_in_do;
  wire _seach_blockx_311_p_reset;
  wire _seach_blockx_311_m_clock;
  wire [9:0] _seach_blockx_310_map_block;
  wire [9:0] _seach_blockx_310_now;
  wire [9:0] _seach_blockx_310_start;
  wire [9:0] _seach_blockx_310_goal;
  wire [9:0] _seach_blockx_310_data_out;
  wire _seach_blockx_310_in_do;
  wire _seach_blockx_310_p_reset;
  wire _seach_blockx_310_m_clock;
  wire [9:0] _seach_blockx_309_map_block;
  wire [9:0] _seach_blockx_309_now;
  wire [9:0] _seach_blockx_309_start;
  wire [9:0] _seach_blockx_309_goal;
  wire [9:0] _seach_blockx_309_data_out;
  wire _seach_blockx_309_in_do;
  wire _seach_blockx_309_p_reset;
  wire _seach_blockx_309_m_clock;
  wire [9:0] _seach_blockx_308_map_block;
  wire [9:0] _seach_blockx_308_now;
  wire [9:0] _seach_blockx_308_start;
  wire [9:0] _seach_blockx_308_goal;
  wire [9:0] _seach_blockx_308_data_out;
  wire _seach_blockx_308_in_do;
  wire _seach_blockx_308_p_reset;
  wire _seach_blockx_308_m_clock;
  wire [9:0] _seach_blockx_307_map_block;
  wire [9:0] _seach_blockx_307_now;
  wire [9:0] _seach_blockx_307_start;
  wire [9:0] _seach_blockx_307_goal;
  wire [9:0] _seach_blockx_307_data_out;
  wire _seach_blockx_307_in_do;
  wire _seach_blockx_307_p_reset;
  wire _seach_blockx_307_m_clock;
  wire [9:0] _seach_blockx_306_map_block;
  wire [9:0] _seach_blockx_306_now;
  wire [9:0] _seach_blockx_306_start;
  wire [9:0] _seach_blockx_306_goal;
  wire [9:0] _seach_blockx_306_data_out;
  wire _seach_blockx_306_in_do;
  wire _seach_blockx_306_p_reset;
  wire _seach_blockx_306_m_clock;
  wire [9:0] _seach_blockx_305_map_block;
  wire [9:0] _seach_blockx_305_now;
  wire [9:0] _seach_blockx_305_start;
  wire [9:0] _seach_blockx_305_goal;
  wire [9:0] _seach_blockx_305_data_out;
  wire _seach_blockx_305_in_do;
  wire _seach_blockx_305_p_reset;
  wire _seach_blockx_305_m_clock;
  wire [9:0] _seach_blockx_304_map_block;
  wire [9:0] _seach_blockx_304_now;
  wire [9:0] _seach_blockx_304_start;
  wire [9:0] _seach_blockx_304_goal;
  wire [9:0] _seach_blockx_304_data_out;
  wire _seach_blockx_304_in_do;
  wire _seach_blockx_304_p_reset;
  wire _seach_blockx_304_m_clock;
  wire [9:0] _seach_blockx_303_map_block;
  wire [9:0] _seach_blockx_303_now;
  wire [9:0] _seach_blockx_303_start;
  wire [9:0] _seach_blockx_303_goal;
  wire [9:0] _seach_blockx_303_data_out;
  wire _seach_blockx_303_in_do;
  wire _seach_blockx_303_p_reset;
  wire _seach_blockx_303_m_clock;
  wire [9:0] _seach_blockx_302_map_block;
  wire [9:0] _seach_blockx_302_now;
  wire [9:0] _seach_blockx_302_start;
  wire [9:0] _seach_blockx_302_goal;
  wire [9:0] _seach_blockx_302_data_out;
  wire _seach_blockx_302_in_do;
  wire _seach_blockx_302_p_reset;
  wire _seach_blockx_302_m_clock;
  wire [9:0] _seach_blockx_301_map_block;
  wire [9:0] _seach_blockx_301_now;
  wire [9:0] _seach_blockx_301_start;
  wire [9:0] _seach_blockx_301_goal;
  wire [9:0] _seach_blockx_301_data_out;
  wire _seach_blockx_301_in_do;
  wire _seach_blockx_301_p_reset;
  wire _seach_blockx_301_m_clock;
  wire [9:0] _seach_blockx_300_map_block;
  wire [9:0] _seach_blockx_300_now;
  wire [9:0] _seach_blockx_300_start;
  wire [9:0] _seach_blockx_300_goal;
  wire [9:0] _seach_blockx_300_data_out;
  wire _seach_blockx_300_in_do;
  wire _seach_blockx_300_p_reset;
  wire _seach_blockx_300_m_clock;
  wire [9:0] _seach_blockx_299_map_block;
  wire [9:0] _seach_blockx_299_now;
  wire [9:0] _seach_blockx_299_start;
  wire [9:0] _seach_blockx_299_goal;
  wire [9:0] _seach_blockx_299_data_out;
  wire _seach_blockx_299_in_do;
  wire _seach_blockx_299_p_reset;
  wire _seach_blockx_299_m_clock;
  wire [9:0] _seach_blockx_298_map_block;
  wire [9:0] _seach_blockx_298_now;
  wire [9:0] _seach_blockx_298_start;
  wire [9:0] _seach_blockx_298_goal;
  wire [9:0] _seach_blockx_298_data_out;
  wire _seach_blockx_298_in_do;
  wire _seach_blockx_298_p_reset;
  wire _seach_blockx_298_m_clock;
  wire [9:0] _seach_blockx_297_map_block;
  wire [9:0] _seach_blockx_297_now;
  wire [9:0] _seach_blockx_297_start;
  wire [9:0] _seach_blockx_297_goal;
  wire [9:0] _seach_blockx_297_data_out;
  wire _seach_blockx_297_in_do;
  wire _seach_blockx_297_p_reset;
  wire _seach_blockx_297_m_clock;
  wire [9:0] _seach_blockx_296_map_block;
  wire [9:0] _seach_blockx_296_now;
  wire [9:0] _seach_blockx_296_start;
  wire [9:0] _seach_blockx_296_goal;
  wire [9:0] _seach_blockx_296_data_out;
  wire _seach_blockx_296_in_do;
  wire _seach_blockx_296_p_reset;
  wire _seach_blockx_296_m_clock;
  wire [9:0] _seach_blockx_295_map_block;
  wire [9:0] _seach_blockx_295_now;
  wire [9:0] _seach_blockx_295_start;
  wire [9:0] _seach_blockx_295_goal;
  wire [9:0] _seach_blockx_295_data_out;
  wire _seach_blockx_295_in_do;
  wire _seach_blockx_295_p_reset;
  wire _seach_blockx_295_m_clock;
  wire [9:0] _seach_blockx_294_map_block;
  wire [9:0] _seach_blockx_294_now;
  wire [9:0] _seach_blockx_294_start;
  wire [9:0] _seach_blockx_294_goal;
  wire [9:0] _seach_blockx_294_data_out;
  wire _seach_blockx_294_in_do;
  wire _seach_blockx_294_p_reset;
  wire _seach_blockx_294_m_clock;
  wire [9:0] _seach_blockx_293_map_block;
  wire [9:0] _seach_blockx_293_now;
  wire [9:0] _seach_blockx_293_start;
  wire [9:0] _seach_blockx_293_goal;
  wire [9:0] _seach_blockx_293_data_out;
  wire _seach_blockx_293_in_do;
  wire _seach_blockx_293_p_reset;
  wire _seach_blockx_293_m_clock;
  wire [9:0] _seach_blockx_292_map_block;
  wire [9:0] _seach_blockx_292_now;
  wire [9:0] _seach_blockx_292_start;
  wire [9:0] _seach_blockx_292_goal;
  wire [9:0] _seach_blockx_292_data_out;
  wire _seach_blockx_292_in_do;
  wire _seach_blockx_292_p_reset;
  wire _seach_blockx_292_m_clock;
  wire [9:0] _seach_blockx_291_map_block;
  wire [9:0] _seach_blockx_291_now;
  wire [9:0] _seach_blockx_291_start;
  wire [9:0] _seach_blockx_291_goal;
  wire [9:0] _seach_blockx_291_data_out;
  wire _seach_blockx_291_in_do;
  wire _seach_blockx_291_p_reset;
  wire _seach_blockx_291_m_clock;
  wire [9:0] _seach_blockx_290_map_block;
  wire [9:0] _seach_blockx_290_now;
  wire [9:0] _seach_blockx_290_start;
  wire [9:0] _seach_blockx_290_goal;
  wire [9:0] _seach_blockx_290_data_out;
  wire _seach_blockx_290_in_do;
  wire _seach_blockx_290_p_reset;
  wire _seach_blockx_290_m_clock;
  wire [9:0] _seach_blockx_289_map_block;
  wire [9:0] _seach_blockx_289_now;
  wire [9:0] _seach_blockx_289_start;
  wire [9:0] _seach_blockx_289_goal;
  wire [9:0] _seach_blockx_289_data_out;
  wire _seach_blockx_289_in_do;
  wire _seach_blockx_289_p_reset;
  wire _seach_blockx_289_m_clock;
  wire [9:0] _seach_blockx_288_map_block;
  wire [9:0] _seach_blockx_288_now;
  wire [9:0] _seach_blockx_288_start;
  wire [9:0] _seach_blockx_288_goal;
  wire [9:0] _seach_blockx_288_data_out;
  wire _seach_blockx_288_in_do;
  wire _seach_blockx_288_p_reset;
  wire _seach_blockx_288_m_clock;
  wire [9:0] _seach_blockx_287_map_block;
  wire [9:0] _seach_blockx_287_now;
  wire [9:0] _seach_blockx_287_start;
  wire [9:0] _seach_blockx_287_goal;
  wire [9:0] _seach_blockx_287_data_out;
  wire _seach_blockx_287_in_do;
  wire _seach_blockx_287_p_reset;
  wire _seach_blockx_287_m_clock;
  wire [9:0] _seach_blockx_286_map_block;
  wire [9:0] _seach_blockx_286_now;
  wire [9:0] _seach_blockx_286_start;
  wire [9:0] _seach_blockx_286_goal;
  wire [9:0] _seach_blockx_286_data_out;
  wire _seach_blockx_286_in_do;
  wire _seach_blockx_286_p_reset;
  wire _seach_blockx_286_m_clock;
  wire [9:0] _seach_blockx_285_map_block;
  wire [9:0] _seach_blockx_285_now;
  wire [9:0] _seach_blockx_285_start;
  wire [9:0] _seach_blockx_285_goal;
  wire [9:0] _seach_blockx_285_data_out;
  wire _seach_blockx_285_in_do;
  wire _seach_blockx_285_p_reset;
  wire _seach_blockx_285_m_clock;
  wire [9:0] _seach_blockx_284_map_block;
  wire [9:0] _seach_blockx_284_now;
  wire [9:0] _seach_blockx_284_start;
  wire [9:0] _seach_blockx_284_goal;
  wire [9:0] _seach_blockx_284_data_out;
  wire _seach_blockx_284_in_do;
  wire _seach_blockx_284_p_reset;
  wire _seach_blockx_284_m_clock;
  wire [9:0] _seach_blockx_283_map_block;
  wire [9:0] _seach_blockx_283_now;
  wire [9:0] _seach_blockx_283_start;
  wire [9:0] _seach_blockx_283_goal;
  wire [9:0] _seach_blockx_283_data_out;
  wire _seach_blockx_283_in_do;
  wire _seach_blockx_283_p_reset;
  wire _seach_blockx_283_m_clock;
  wire [9:0] _seach_blockx_282_map_block;
  wire [9:0] _seach_blockx_282_now;
  wire [9:0] _seach_blockx_282_start;
  wire [9:0] _seach_blockx_282_goal;
  wire [9:0] _seach_blockx_282_data_out;
  wire _seach_blockx_282_in_do;
  wire _seach_blockx_282_p_reset;
  wire _seach_blockx_282_m_clock;
  wire [9:0] _seach_blockx_281_map_block;
  wire [9:0] _seach_blockx_281_now;
  wire [9:0] _seach_blockx_281_start;
  wire [9:0] _seach_blockx_281_goal;
  wire [9:0] _seach_blockx_281_data_out;
  wire _seach_blockx_281_in_do;
  wire _seach_blockx_281_p_reset;
  wire _seach_blockx_281_m_clock;
  wire [9:0] _seach_blockx_280_map_block;
  wire [9:0] _seach_blockx_280_now;
  wire [9:0] _seach_blockx_280_start;
  wire [9:0] _seach_blockx_280_goal;
  wire [9:0] _seach_blockx_280_data_out;
  wire _seach_blockx_280_in_do;
  wire _seach_blockx_280_p_reset;
  wire _seach_blockx_280_m_clock;
  wire [9:0] _seach_blockx_279_map_block;
  wire [9:0] _seach_blockx_279_now;
  wire [9:0] _seach_blockx_279_start;
  wire [9:0] _seach_blockx_279_goal;
  wire [9:0] _seach_blockx_279_data_out;
  wire _seach_blockx_279_in_do;
  wire _seach_blockx_279_p_reset;
  wire _seach_blockx_279_m_clock;
  wire [9:0] _seach_blockx_278_map_block;
  wire [9:0] _seach_blockx_278_now;
  wire [9:0] _seach_blockx_278_start;
  wire [9:0] _seach_blockx_278_goal;
  wire [9:0] _seach_blockx_278_data_out;
  wire _seach_blockx_278_in_do;
  wire _seach_blockx_278_p_reset;
  wire _seach_blockx_278_m_clock;
  wire [9:0] _seach_blockx_277_map_block;
  wire [9:0] _seach_blockx_277_now;
  wire [9:0] _seach_blockx_277_start;
  wire [9:0] _seach_blockx_277_goal;
  wire [9:0] _seach_blockx_277_data_out;
  wire _seach_blockx_277_in_do;
  wire _seach_blockx_277_p_reset;
  wire _seach_blockx_277_m_clock;
  wire [9:0] _seach_blockx_276_map_block;
  wire [9:0] _seach_blockx_276_now;
  wire [9:0] _seach_blockx_276_start;
  wire [9:0] _seach_blockx_276_goal;
  wire [9:0] _seach_blockx_276_data_out;
  wire _seach_blockx_276_in_do;
  wire _seach_blockx_276_p_reset;
  wire _seach_blockx_276_m_clock;
  wire [9:0] _seach_blockx_275_map_block;
  wire [9:0] _seach_blockx_275_now;
  wire [9:0] _seach_blockx_275_start;
  wire [9:0] _seach_blockx_275_goal;
  wire [9:0] _seach_blockx_275_data_out;
  wire _seach_blockx_275_in_do;
  wire _seach_blockx_275_p_reset;
  wire _seach_blockx_275_m_clock;
  wire [9:0] _seach_blockx_274_map_block;
  wire [9:0] _seach_blockx_274_now;
  wire [9:0] _seach_blockx_274_start;
  wire [9:0] _seach_blockx_274_goal;
  wire [9:0] _seach_blockx_274_data_out;
  wire _seach_blockx_274_in_do;
  wire _seach_blockx_274_p_reset;
  wire _seach_blockx_274_m_clock;
  wire [9:0] _seach_blockx_273_map_block;
  wire [9:0] _seach_blockx_273_now;
  wire [9:0] _seach_blockx_273_start;
  wire [9:0] _seach_blockx_273_goal;
  wire [9:0] _seach_blockx_273_data_out;
  wire _seach_blockx_273_in_do;
  wire _seach_blockx_273_p_reset;
  wire _seach_blockx_273_m_clock;
  wire [9:0] _seach_blockx_272_map_block;
  wire [9:0] _seach_blockx_272_now;
  wire [9:0] _seach_blockx_272_start;
  wire [9:0] _seach_blockx_272_goal;
  wire [9:0] _seach_blockx_272_data_out;
  wire _seach_blockx_272_in_do;
  wire _seach_blockx_272_p_reset;
  wire _seach_blockx_272_m_clock;
  wire [9:0] _seach_blockx_271_map_block;
  wire [9:0] _seach_blockx_271_now;
  wire [9:0] _seach_blockx_271_start;
  wire [9:0] _seach_blockx_271_goal;
  wire [9:0] _seach_blockx_271_data_out;
  wire _seach_blockx_271_in_do;
  wire _seach_blockx_271_p_reset;
  wire _seach_blockx_271_m_clock;
  wire [9:0] _seach_blockx_270_map_block;
  wire [9:0] _seach_blockx_270_now;
  wire [9:0] _seach_blockx_270_start;
  wire [9:0] _seach_blockx_270_goal;
  wire [9:0] _seach_blockx_270_data_out;
  wire _seach_blockx_270_in_do;
  wire _seach_blockx_270_p_reset;
  wire _seach_blockx_270_m_clock;
  wire [9:0] _seach_blockx_269_map_block;
  wire [9:0] _seach_blockx_269_now;
  wire [9:0] _seach_blockx_269_start;
  wire [9:0] _seach_blockx_269_goal;
  wire [9:0] _seach_blockx_269_data_out;
  wire _seach_blockx_269_in_do;
  wire _seach_blockx_269_p_reset;
  wire _seach_blockx_269_m_clock;
  wire [9:0] _seach_blockx_268_map_block;
  wire [9:0] _seach_blockx_268_now;
  wire [9:0] _seach_blockx_268_start;
  wire [9:0] _seach_blockx_268_goal;
  wire [9:0] _seach_blockx_268_data_out;
  wire _seach_blockx_268_in_do;
  wire _seach_blockx_268_p_reset;
  wire _seach_blockx_268_m_clock;
  wire [9:0] _seach_blockx_267_map_block;
  wire [9:0] _seach_blockx_267_now;
  wire [9:0] _seach_blockx_267_start;
  wire [9:0] _seach_blockx_267_goal;
  wire [9:0] _seach_blockx_267_data_out;
  wire _seach_blockx_267_in_do;
  wire _seach_blockx_267_p_reset;
  wire _seach_blockx_267_m_clock;
  wire [9:0] _seach_blockx_266_map_block;
  wire [9:0] _seach_blockx_266_now;
  wire [9:0] _seach_blockx_266_start;
  wire [9:0] _seach_blockx_266_goal;
  wire [9:0] _seach_blockx_266_data_out;
  wire _seach_blockx_266_in_do;
  wire _seach_blockx_266_p_reset;
  wire _seach_blockx_266_m_clock;
  wire [9:0] _seach_blockx_265_map_block;
  wire [9:0] _seach_blockx_265_now;
  wire [9:0] _seach_blockx_265_start;
  wire [9:0] _seach_blockx_265_goal;
  wire [9:0] _seach_blockx_265_data_out;
  wire _seach_blockx_265_in_do;
  wire _seach_blockx_265_p_reset;
  wire _seach_blockx_265_m_clock;
  wire [9:0] _seach_blockx_264_map_block;
  wire [9:0] _seach_blockx_264_now;
  wire [9:0] _seach_blockx_264_start;
  wire [9:0] _seach_blockx_264_goal;
  wire [9:0] _seach_blockx_264_data_out;
  wire _seach_blockx_264_in_do;
  wire _seach_blockx_264_p_reset;
  wire _seach_blockx_264_m_clock;
  wire [9:0] _seach_blockx_263_map_block;
  wire [9:0] _seach_blockx_263_now;
  wire [9:0] _seach_blockx_263_start;
  wire [9:0] _seach_blockx_263_goal;
  wire [9:0] _seach_blockx_263_data_out;
  wire _seach_blockx_263_in_do;
  wire _seach_blockx_263_p_reset;
  wire _seach_blockx_263_m_clock;
  wire [9:0] _seach_blockx_262_map_block;
  wire [9:0] _seach_blockx_262_now;
  wire [9:0] _seach_blockx_262_start;
  wire [9:0] _seach_blockx_262_goal;
  wire [9:0] _seach_blockx_262_data_out;
  wire _seach_blockx_262_in_do;
  wire _seach_blockx_262_p_reset;
  wire _seach_blockx_262_m_clock;
  wire [9:0] _seach_blockx_261_map_block;
  wire [9:0] _seach_blockx_261_now;
  wire [9:0] _seach_blockx_261_start;
  wire [9:0] _seach_blockx_261_goal;
  wire [9:0] _seach_blockx_261_data_out;
  wire _seach_blockx_261_in_do;
  wire _seach_blockx_261_p_reset;
  wire _seach_blockx_261_m_clock;
  wire [9:0] _seach_blockx_260_map_block;
  wire [9:0] _seach_blockx_260_now;
  wire [9:0] _seach_blockx_260_start;
  wire [9:0] _seach_blockx_260_goal;
  wire [9:0] _seach_blockx_260_data_out;
  wire _seach_blockx_260_in_do;
  wire _seach_blockx_260_p_reset;
  wire _seach_blockx_260_m_clock;
  wire [9:0] _seach_blockx_259_map_block;
  wire [9:0] _seach_blockx_259_now;
  wire [9:0] _seach_blockx_259_start;
  wire [9:0] _seach_blockx_259_goal;
  wire [9:0] _seach_blockx_259_data_out;
  wire _seach_blockx_259_in_do;
  wire _seach_blockx_259_p_reset;
  wire _seach_blockx_259_m_clock;
  wire [9:0] _seach_blockx_258_map_block;
  wire [9:0] _seach_blockx_258_now;
  wire [9:0] _seach_blockx_258_start;
  wire [9:0] _seach_blockx_258_goal;
  wire [9:0] _seach_blockx_258_data_out;
  wire _seach_blockx_258_in_do;
  wire _seach_blockx_258_p_reset;
  wire _seach_blockx_258_m_clock;
  wire [9:0] _seach_blockx_257_map_block;
  wire [9:0] _seach_blockx_257_now;
  wire [9:0] _seach_blockx_257_start;
  wire [9:0] _seach_blockx_257_goal;
  wire [9:0] _seach_blockx_257_data_out;
  wire _seach_blockx_257_in_do;
  wire _seach_blockx_257_p_reset;
  wire _seach_blockx_257_m_clock;
  wire [9:0] _seach_blockx_256_map_block;
  wire [9:0] _seach_blockx_256_now;
  wire [9:0] _seach_blockx_256_start;
  wire [9:0] _seach_blockx_256_goal;
  wire [9:0] _seach_blockx_256_data_out;
  wire _seach_blockx_256_in_do;
  wire _seach_blockx_256_p_reset;
  wire _seach_blockx_256_m_clock;
  wire [9:0] _seach_blockx_255_map_block;
  wire [9:0] _seach_blockx_255_now;
  wire [9:0] _seach_blockx_255_start;
  wire [9:0] _seach_blockx_255_goal;
  wire [9:0] _seach_blockx_255_data_out;
  wire _seach_blockx_255_in_do;
  wire _seach_blockx_255_p_reset;
  wire _seach_blockx_255_m_clock;
  wire [9:0] _seach_blockx_254_map_block;
  wire [9:0] _seach_blockx_254_now;
  wire [9:0] _seach_blockx_254_start;
  wire [9:0] _seach_blockx_254_goal;
  wire [9:0] _seach_blockx_254_data_out;
  wire _seach_blockx_254_in_do;
  wire _seach_blockx_254_p_reset;
  wire _seach_blockx_254_m_clock;
  wire [9:0] _seach_blockx_253_map_block;
  wire [9:0] _seach_blockx_253_now;
  wire [9:0] _seach_blockx_253_start;
  wire [9:0] _seach_blockx_253_goal;
  wire [9:0] _seach_blockx_253_data_out;
  wire _seach_blockx_253_in_do;
  wire _seach_blockx_253_p_reset;
  wire _seach_blockx_253_m_clock;
  wire [9:0] _seach_blockx_252_map_block;
  wire [9:0] _seach_blockx_252_now;
  wire [9:0] _seach_blockx_252_start;
  wire [9:0] _seach_blockx_252_goal;
  wire [9:0] _seach_blockx_252_data_out;
  wire _seach_blockx_252_in_do;
  wire _seach_blockx_252_p_reset;
  wire _seach_blockx_252_m_clock;
  wire [9:0] _seach_blockx_251_map_block;
  wire [9:0] _seach_blockx_251_now;
  wire [9:0] _seach_blockx_251_start;
  wire [9:0] _seach_blockx_251_goal;
  wire [9:0] _seach_blockx_251_data_out;
  wire _seach_blockx_251_in_do;
  wire _seach_blockx_251_p_reset;
  wire _seach_blockx_251_m_clock;
  wire [9:0] _seach_blockx_250_map_block;
  wire [9:0] _seach_blockx_250_now;
  wire [9:0] _seach_blockx_250_start;
  wire [9:0] _seach_blockx_250_goal;
  wire [9:0] _seach_blockx_250_data_out;
  wire _seach_blockx_250_in_do;
  wire _seach_blockx_250_p_reset;
  wire _seach_blockx_250_m_clock;
  wire [9:0] _seach_blockx_249_map_block;
  wire [9:0] _seach_blockx_249_now;
  wire [9:0] _seach_blockx_249_start;
  wire [9:0] _seach_blockx_249_goal;
  wire [9:0] _seach_blockx_249_data_out;
  wire _seach_blockx_249_in_do;
  wire _seach_blockx_249_p_reset;
  wire _seach_blockx_249_m_clock;
  wire [9:0] _seach_blockx_248_map_block;
  wire [9:0] _seach_blockx_248_now;
  wire [9:0] _seach_blockx_248_start;
  wire [9:0] _seach_blockx_248_goal;
  wire [9:0] _seach_blockx_248_data_out;
  wire _seach_blockx_248_in_do;
  wire _seach_blockx_248_p_reset;
  wire _seach_blockx_248_m_clock;
  wire [9:0] _seach_blockx_247_map_block;
  wire [9:0] _seach_blockx_247_now;
  wire [9:0] _seach_blockx_247_start;
  wire [9:0] _seach_blockx_247_goal;
  wire [9:0] _seach_blockx_247_data_out;
  wire _seach_blockx_247_in_do;
  wire _seach_blockx_247_p_reset;
  wire _seach_blockx_247_m_clock;
  wire [9:0] _seach_blockx_246_map_block;
  wire [9:0] _seach_blockx_246_now;
  wire [9:0] _seach_blockx_246_start;
  wire [9:0] _seach_blockx_246_goal;
  wire [9:0] _seach_blockx_246_data_out;
  wire _seach_blockx_246_in_do;
  wire _seach_blockx_246_p_reset;
  wire _seach_blockx_246_m_clock;
  wire [9:0] _seach_blockx_245_map_block;
  wire [9:0] _seach_blockx_245_now;
  wire [9:0] _seach_blockx_245_start;
  wire [9:0] _seach_blockx_245_goal;
  wire [9:0] _seach_blockx_245_data_out;
  wire _seach_blockx_245_in_do;
  wire _seach_blockx_245_p_reset;
  wire _seach_blockx_245_m_clock;
  wire [9:0] _seach_blockx_244_map_block;
  wire [9:0] _seach_blockx_244_now;
  wire [9:0] _seach_blockx_244_start;
  wire [9:0] _seach_blockx_244_goal;
  wire [9:0] _seach_blockx_244_data_out;
  wire _seach_blockx_244_in_do;
  wire _seach_blockx_244_p_reset;
  wire _seach_blockx_244_m_clock;
  wire [9:0] _seach_blockx_243_map_block;
  wire [9:0] _seach_blockx_243_now;
  wire [9:0] _seach_blockx_243_start;
  wire [9:0] _seach_blockx_243_goal;
  wire [9:0] _seach_blockx_243_data_out;
  wire _seach_blockx_243_in_do;
  wire _seach_blockx_243_p_reset;
  wire _seach_blockx_243_m_clock;
  wire [9:0] _seach_blockx_242_map_block;
  wire [9:0] _seach_blockx_242_now;
  wire [9:0] _seach_blockx_242_start;
  wire [9:0] _seach_blockx_242_goal;
  wire [9:0] _seach_blockx_242_data_out;
  wire _seach_blockx_242_in_do;
  wire _seach_blockx_242_p_reset;
  wire _seach_blockx_242_m_clock;
  wire [9:0] _seach_blockx_241_map_block;
  wire [9:0] _seach_blockx_241_now;
  wire [9:0] _seach_blockx_241_start;
  wire [9:0] _seach_blockx_241_goal;
  wire [9:0] _seach_blockx_241_data_out;
  wire _seach_blockx_241_in_do;
  wire _seach_blockx_241_p_reset;
  wire _seach_blockx_241_m_clock;
  wire [9:0] _seach_blockx_240_map_block;
  wire [9:0] _seach_blockx_240_now;
  wire [9:0] _seach_blockx_240_start;
  wire [9:0] _seach_blockx_240_goal;
  wire [9:0] _seach_blockx_240_data_out;
  wire _seach_blockx_240_in_do;
  wire _seach_blockx_240_p_reset;
  wire _seach_blockx_240_m_clock;
  wire [9:0] _seach_blockx_239_map_block;
  wire [9:0] _seach_blockx_239_now;
  wire [9:0] _seach_blockx_239_start;
  wire [9:0] _seach_blockx_239_goal;
  wire [9:0] _seach_blockx_239_data_out;
  wire _seach_blockx_239_in_do;
  wire _seach_blockx_239_p_reset;
  wire _seach_blockx_239_m_clock;
  wire [9:0] _seach_blockx_238_map_block;
  wire [9:0] _seach_blockx_238_now;
  wire [9:0] _seach_blockx_238_start;
  wire [9:0] _seach_blockx_238_goal;
  wire [9:0] _seach_blockx_238_data_out;
  wire _seach_blockx_238_in_do;
  wire _seach_blockx_238_p_reset;
  wire _seach_blockx_238_m_clock;
  wire [9:0] _seach_blockx_237_map_block;
  wire [9:0] _seach_blockx_237_now;
  wire [9:0] _seach_blockx_237_start;
  wire [9:0] _seach_blockx_237_goal;
  wire [9:0] _seach_blockx_237_data_out;
  wire _seach_blockx_237_in_do;
  wire _seach_blockx_237_p_reset;
  wire _seach_blockx_237_m_clock;
  wire [9:0] _seach_blockx_236_map_block;
  wire [9:0] _seach_blockx_236_now;
  wire [9:0] _seach_blockx_236_start;
  wire [9:0] _seach_blockx_236_goal;
  wire [9:0] _seach_blockx_236_data_out;
  wire _seach_blockx_236_in_do;
  wire _seach_blockx_236_p_reset;
  wire _seach_blockx_236_m_clock;
  wire [9:0] _seach_blockx_235_map_block;
  wire [9:0] _seach_blockx_235_now;
  wire [9:0] _seach_blockx_235_start;
  wire [9:0] _seach_blockx_235_goal;
  wire [9:0] _seach_blockx_235_data_out;
  wire _seach_blockx_235_in_do;
  wire _seach_blockx_235_p_reset;
  wire _seach_blockx_235_m_clock;
  wire [9:0] _seach_blockx_234_map_block;
  wire [9:0] _seach_blockx_234_now;
  wire [9:0] _seach_blockx_234_start;
  wire [9:0] _seach_blockx_234_goal;
  wire [9:0] _seach_blockx_234_data_out;
  wire _seach_blockx_234_in_do;
  wire _seach_blockx_234_p_reset;
  wire _seach_blockx_234_m_clock;
  wire [9:0] _seach_blockx_233_map_block;
  wire [9:0] _seach_blockx_233_now;
  wire [9:0] _seach_blockx_233_start;
  wire [9:0] _seach_blockx_233_goal;
  wire [9:0] _seach_blockx_233_data_out;
  wire _seach_blockx_233_in_do;
  wire _seach_blockx_233_p_reset;
  wire _seach_blockx_233_m_clock;
  wire [9:0] _seach_blockx_232_map_block;
  wire [9:0] _seach_blockx_232_now;
  wire [9:0] _seach_blockx_232_start;
  wire [9:0] _seach_blockx_232_goal;
  wire [9:0] _seach_blockx_232_data_out;
  wire _seach_blockx_232_in_do;
  wire _seach_blockx_232_p_reset;
  wire _seach_blockx_232_m_clock;
  wire [9:0] _seach_blockx_231_map_block;
  wire [9:0] _seach_blockx_231_now;
  wire [9:0] _seach_blockx_231_start;
  wire [9:0] _seach_blockx_231_goal;
  wire [9:0] _seach_blockx_231_data_out;
  wire _seach_blockx_231_in_do;
  wire _seach_blockx_231_p_reset;
  wire _seach_blockx_231_m_clock;
  wire [9:0] _seach_blockx_230_map_block;
  wire [9:0] _seach_blockx_230_now;
  wire [9:0] _seach_blockx_230_start;
  wire [9:0] _seach_blockx_230_goal;
  wire [9:0] _seach_blockx_230_data_out;
  wire _seach_blockx_230_in_do;
  wire _seach_blockx_230_p_reset;
  wire _seach_blockx_230_m_clock;
  wire [9:0] _seach_blockx_229_map_block;
  wire [9:0] _seach_blockx_229_now;
  wire [9:0] _seach_blockx_229_start;
  wire [9:0] _seach_blockx_229_goal;
  wire [9:0] _seach_blockx_229_data_out;
  wire _seach_blockx_229_in_do;
  wire _seach_blockx_229_p_reset;
  wire _seach_blockx_229_m_clock;
  wire [9:0] _seach_blockx_228_map_block;
  wire [9:0] _seach_blockx_228_now;
  wire [9:0] _seach_blockx_228_start;
  wire [9:0] _seach_blockx_228_goal;
  wire [9:0] _seach_blockx_228_data_out;
  wire _seach_blockx_228_in_do;
  wire _seach_blockx_228_p_reset;
  wire _seach_blockx_228_m_clock;
  wire [9:0] _seach_blockx_227_map_block;
  wire [9:0] _seach_blockx_227_now;
  wire [9:0] _seach_blockx_227_start;
  wire [9:0] _seach_blockx_227_goal;
  wire [9:0] _seach_blockx_227_data_out;
  wire _seach_blockx_227_in_do;
  wire _seach_blockx_227_p_reset;
  wire _seach_blockx_227_m_clock;
  wire [9:0] _seach_blockx_226_map_block;
  wire [9:0] _seach_blockx_226_now;
  wire [9:0] _seach_blockx_226_start;
  wire [9:0] _seach_blockx_226_goal;
  wire [9:0] _seach_blockx_226_data_out;
  wire _seach_blockx_226_in_do;
  wire _seach_blockx_226_p_reset;
  wire _seach_blockx_226_m_clock;
  wire [9:0] _seach_blockx_225_map_block;
  wire [9:0] _seach_blockx_225_now;
  wire [9:0] _seach_blockx_225_start;
  wire [9:0] _seach_blockx_225_goal;
  wire [9:0] _seach_blockx_225_data_out;
  wire _seach_blockx_225_in_do;
  wire _seach_blockx_225_p_reset;
  wire _seach_blockx_225_m_clock;
  wire [9:0] _seach_blockx_224_map_block;
  wire [9:0] _seach_blockx_224_now;
  wire [9:0] _seach_blockx_224_start;
  wire [9:0] _seach_blockx_224_goal;
  wire [9:0] _seach_blockx_224_data_out;
  wire _seach_blockx_224_in_do;
  wire _seach_blockx_224_p_reset;
  wire _seach_blockx_224_m_clock;
  wire [9:0] _seach_blockx_223_map_block;
  wire [9:0] _seach_blockx_223_now;
  wire [9:0] _seach_blockx_223_start;
  wire [9:0] _seach_blockx_223_goal;
  wire [9:0] _seach_blockx_223_data_out;
  wire _seach_blockx_223_in_do;
  wire _seach_blockx_223_p_reset;
  wire _seach_blockx_223_m_clock;
  wire [9:0] _seach_blockx_222_map_block;
  wire [9:0] _seach_blockx_222_now;
  wire [9:0] _seach_blockx_222_start;
  wire [9:0] _seach_blockx_222_goal;
  wire [9:0] _seach_blockx_222_data_out;
  wire _seach_blockx_222_in_do;
  wire _seach_blockx_222_p_reset;
  wire _seach_blockx_222_m_clock;
  wire [9:0] _seach_blockx_221_map_block;
  wire [9:0] _seach_blockx_221_now;
  wire [9:0] _seach_blockx_221_start;
  wire [9:0] _seach_blockx_221_goal;
  wire [9:0] _seach_blockx_221_data_out;
  wire _seach_blockx_221_in_do;
  wire _seach_blockx_221_p_reset;
  wire _seach_blockx_221_m_clock;
  wire [9:0] _seach_blockx_220_map_block;
  wire [9:0] _seach_blockx_220_now;
  wire [9:0] _seach_blockx_220_start;
  wire [9:0] _seach_blockx_220_goal;
  wire [9:0] _seach_blockx_220_data_out;
  wire _seach_blockx_220_in_do;
  wire _seach_blockx_220_p_reset;
  wire _seach_blockx_220_m_clock;
  wire [9:0] _seach_blockx_219_map_block;
  wire [9:0] _seach_blockx_219_now;
  wire [9:0] _seach_blockx_219_start;
  wire [9:0] _seach_blockx_219_goal;
  wire [9:0] _seach_blockx_219_data_out;
  wire _seach_blockx_219_in_do;
  wire _seach_blockx_219_p_reset;
  wire _seach_blockx_219_m_clock;
  wire [9:0] _seach_blockx_218_map_block;
  wire [9:0] _seach_blockx_218_now;
  wire [9:0] _seach_blockx_218_start;
  wire [9:0] _seach_blockx_218_goal;
  wire [9:0] _seach_blockx_218_data_out;
  wire _seach_blockx_218_in_do;
  wire _seach_blockx_218_p_reset;
  wire _seach_blockx_218_m_clock;
  wire [9:0] _seach_blockx_217_map_block;
  wire [9:0] _seach_blockx_217_now;
  wire [9:0] _seach_blockx_217_start;
  wire [9:0] _seach_blockx_217_goal;
  wire [9:0] _seach_blockx_217_data_out;
  wire _seach_blockx_217_in_do;
  wire _seach_blockx_217_p_reset;
  wire _seach_blockx_217_m_clock;
  wire [9:0] _seach_blockx_216_map_block;
  wire [9:0] _seach_blockx_216_now;
  wire [9:0] _seach_blockx_216_start;
  wire [9:0] _seach_blockx_216_goal;
  wire [9:0] _seach_blockx_216_data_out;
  wire _seach_blockx_216_in_do;
  wire _seach_blockx_216_p_reset;
  wire _seach_blockx_216_m_clock;
  wire [9:0] _seach_blockx_215_map_block;
  wire [9:0] _seach_blockx_215_now;
  wire [9:0] _seach_blockx_215_start;
  wire [9:0] _seach_blockx_215_goal;
  wire [9:0] _seach_blockx_215_data_out;
  wire _seach_blockx_215_in_do;
  wire _seach_blockx_215_p_reset;
  wire _seach_blockx_215_m_clock;
  wire [9:0] _seach_blockx_214_map_block;
  wire [9:0] _seach_blockx_214_now;
  wire [9:0] _seach_blockx_214_start;
  wire [9:0] _seach_blockx_214_goal;
  wire [9:0] _seach_blockx_214_data_out;
  wire _seach_blockx_214_in_do;
  wire _seach_blockx_214_p_reset;
  wire _seach_blockx_214_m_clock;
  wire [9:0] _seach_blockx_213_map_block;
  wire [9:0] _seach_blockx_213_now;
  wire [9:0] _seach_blockx_213_start;
  wire [9:0] _seach_blockx_213_goal;
  wire [9:0] _seach_blockx_213_data_out;
  wire _seach_blockx_213_in_do;
  wire _seach_blockx_213_p_reset;
  wire _seach_blockx_213_m_clock;
  wire [9:0] _seach_blockx_212_map_block;
  wire [9:0] _seach_blockx_212_now;
  wire [9:0] _seach_blockx_212_start;
  wire [9:0] _seach_blockx_212_goal;
  wire [9:0] _seach_blockx_212_data_out;
  wire _seach_blockx_212_in_do;
  wire _seach_blockx_212_p_reset;
  wire _seach_blockx_212_m_clock;
  wire [9:0] _seach_blockx_211_map_block;
  wire [9:0] _seach_blockx_211_now;
  wire [9:0] _seach_blockx_211_start;
  wire [9:0] _seach_blockx_211_goal;
  wire [9:0] _seach_blockx_211_data_out;
  wire _seach_blockx_211_in_do;
  wire _seach_blockx_211_p_reset;
  wire _seach_blockx_211_m_clock;
  wire [9:0] _seach_blockx_210_map_block;
  wire [9:0] _seach_blockx_210_now;
  wire [9:0] _seach_blockx_210_start;
  wire [9:0] _seach_blockx_210_goal;
  wire [9:0] _seach_blockx_210_data_out;
  wire _seach_blockx_210_in_do;
  wire _seach_blockx_210_p_reset;
  wire _seach_blockx_210_m_clock;
  wire [9:0] _seach_blockx_209_map_block;
  wire [9:0] _seach_blockx_209_now;
  wire [9:0] _seach_blockx_209_start;
  wire [9:0] _seach_blockx_209_goal;
  wire [9:0] _seach_blockx_209_data_out;
  wire _seach_blockx_209_in_do;
  wire _seach_blockx_209_p_reset;
  wire _seach_blockx_209_m_clock;
  wire [9:0] _seach_blockx_208_map_block;
  wire [9:0] _seach_blockx_208_now;
  wire [9:0] _seach_blockx_208_start;
  wire [9:0] _seach_blockx_208_goal;
  wire [9:0] _seach_blockx_208_data_out;
  wire _seach_blockx_208_in_do;
  wire _seach_blockx_208_p_reset;
  wire _seach_blockx_208_m_clock;
  wire [9:0] _seach_blockx_207_map_block;
  wire [9:0] _seach_blockx_207_now;
  wire [9:0] _seach_blockx_207_start;
  wire [9:0] _seach_blockx_207_goal;
  wire [9:0] _seach_blockx_207_data_out;
  wire _seach_blockx_207_in_do;
  wire _seach_blockx_207_p_reset;
  wire _seach_blockx_207_m_clock;
  wire [9:0] _seach_blockx_206_map_block;
  wire [9:0] _seach_blockx_206_now;
  wire [9:0] _seach_blockx_206_start;
  wire [9:0] _seach_blockx_206_goal;
  wire [9:0] _seach_blockx_206_data_out;
  wire _seach_blockx_206_in_do;
  wire _seach_blockx_206_p_reset;
  wire _seach_blockx_206_m_clock;
  wire [9:0] _seach_blockx_205_map_block;
  wire [9:0] _seach_blockx_205_now;
  wire [9:0] _seach_blockx_205_start;
  wire [9:0] _seach_blockx_205_goal;
  wire [9:0] _seach_blockx_205_data_out;
  wire _seach_blockx_205_in_do;
  wire _seach_blockx_205_p_reset;
  wire _seach_blockx_205_m_clock;
  wire [9:0] _seach_blockx_204_map_block;
  wire [9:0] _seach_blockx_204_now;
  wire [9:0] _seach_blockx_204_start;
  wire [9:0] _seach_blockx_204_goal;
  wire [9:0] _seach_blockx_204_data_out;
  wire _seach_blockx_204_in_do;
  wire _seach_blockx_204_p_reset;
  wire _seach_blockx_204_m_clock;
  wire [9:0] _seach_blockx_203_map_block;
  wire [9:0] _seach_blockx_203_now;
  wire [9:0] _seach_blockx_203_start;
  wire [9:0] _seach_blockx_203_goal;
  wire [9:0] _seach_blockx_203_data_out;
  wire _seach_blockx_203_in_do;
  wire _seach_blockx_203_p_reset;
  wire _seach_blockx_203_m_clock;
  wire [9:0] _seach_blockx_202_map_block;
  wire [9:0] _seach_blockx_202_now;
  wire [9:0] _seach_blockx_202_start;
  wire [9:0] _seach_blockx_202_goal;
  wire [9:0] _seach_blockx_202_data_out;
  wire _seach_blockx_202_in_do;
  wire _seach_blockx_202_p_reset;
  wire _seach_blockx_202_m_clock;
  wire [9:0] _seach_blockx_201_map_block;
  wire [9:0] _seach_blockx_201_now;
  wire [9:0] _seach_blockx_201_start;
  wire [9:0] _seach_blockx_201_goal;
  wire [9:0] _seach_blockx_201_data_out;
  wire _seach_blockx_201_in_do;
  wire _seach_blockx_201_p_reset;
  wire _seach_blockx_201_m_clock;
  wire [9:0] _seach_blockx_200_map_block;
  wire [9:0] _seach_blockx_200_now;
  wire [9:0] _seach_blockx_200_start;
  wire [9:0] _seach_blockx_200_goal;
  wire [9:0] _seach_blockx_200_data_out;
  wire _seach_blockx_200_in_do;
  wire _seach_blockx_200_p_reset;
  wire _seach_blockx_200_m_clock;
  wire [9:0] _seach_blockx_199_map_block;
  wire [9:0] _seach_blockx_199_now;
  wire [9:0] _seach_blockx_199_start;
  wire [9:0] _seach_blockx_199_goal;
  wire [9:0] _seach_blockx_199_data_out;
  wire _seach_blockx_199_in_do;
  wire _seach_blockx_199_p_reset;
  wire _seach_blockx_199_m_clock;
  wire [9:0] _seach_blockx_198_map_block;
  wire [9:0] _seach_blockx_198_now;
  wire [9:0] _seach_blockx_198_start;
  wire [9:0] _seach_blockx_198_goal;
  wire [9:0] _seach_blockx_198_data_out;
  wire _seach_blockx_198_in_do;
  wire _seach_blockx_198_p_reset;
  wire _seach_blockx_198_m_clock;
  wire [9:0] _seach_blockx_197_map_block;
  wire [9:0] _seach_blockx_197_now;
  wire [9:0] _seach_blockx_197_start;
  wire [9:0] _seach_blockx_197_goal;
  wire [9:0] _seach_blockx_197_data_out;
  wire _seach_blockx_197_in_do;
  wire _seach_blockx_197_p_reset;
  wire _seach_blockx_197_m_clock;
  wire [9:0] _seach_blockx_196_map_block;
  wire [9:0] _seach_blockx_196_now;
  wire [9:0] _seach_blockx_196_start;
  wire [9:0] _seach_blockx_196_goal;
  wire [9:0] _seach_blockx_196_data_out;
  wire _seach_blockx_196_in_do;
  wire _seach_blockx_196_p_reset;
  wire _seach_blockx_196_m_clock;
  wire [9:0] _seach_blockx_195_map_block;
  wire [9:0] _seach_blockx_195_now;
  wire [9:0] _seach_blockx_195_start;
  wire [9:0] _seach_blockx_195_goal;
  wire [9:0] _seach_blockx_195_data_out;
  wire _seach_blockx_195_in_do;
  wire _seach_blockx_195_p_reset;
  wire _seach_blockx_195_m_clock;
  wire [9:0] _seach_blockx_194_map_block;
  wire [9:0] _seach_blockx_194_now;
  wire [9:0] _seach_blockx_194_start;
  wire [9:0] _seach_blockx_194_goal;
  wire [9:0] _seach_blockx_194_data_out;
  wire _seach_blockx_194_in_do;
  wire _seach_blockx_194_p_reset;
  wire _seach_blockx_194_m_clock;
  wire [9:0] _seach_blockx_193_map_block;
  wire [9:0] _seach_blockx_193_now;
  wire [9:0] _seach_blockx_193_start;
  wire [9:0] _seach_blockx_193_goal;
  wire [9:0] _seach_blockx_193_data_out;
  wire _seach_blockx_193_in_do;
  wire _seach_blockx_193_p_reset;
  wire _seach_blockx_193_m_clock;
  wire [9:0] _seach_blockx_192_map_block;
  wire [9:0] _seach_blockx_192_now;
  wire [9:0] _seach_blockx_192_start;
  wire [9:0] _seach_blockx_192_goal;
  wire [9:0] _seach_blockx_192_data_out;
  wire _seach_blockx_192_in_do;
  wire _seach_blockx_192_p_reset;
  wire _seach_blockx_192_m_clock;
  wire [9:0] _seach_blockx_191_map_block;
  wire [9:0] _seach_blockx_191_now;
  wire [9:0] _seach_blockx_191_start;
  wire [9:0] _seach_blockx_191_goal;
  wire [9:0] _seach_blockx_191_data_out;
  wire _seach_blockx_191_in_do;
  wire _seach_blockx_191_p_reset;
  wire _seach_blockx_191_m_clock;
  wire [9:0] _seach_blockx_190_map_block;
  wire [9:0] _seach_blockx_190_now;
  wire [9:0] _seach_blockx_190_start;
  wire [9:0] _seach_blockx_190_goal;
  wire [9:0] _seach_blockx_190_data_out;
  wire _seach_blockx_190_in_do;
  wire _seach_blockx_190_p_reset;
  wire _seach_blockx_190_m_clock;
  wire [9:0] _seach_blockx_189_map_block;
  wire [9:0] _seach_blockx_189_now;
  wire [9:0] _seach_blockx_189_start;
  wire [9:0] _seach_blockx_189_goal;
  wire [9:0] _seach_blockx_189_data_out;
  wire _seach_blockx_189_in_do;
  wire _seach_blockx_189_p_reset;
  wire _seach_blockx_189_m_clock;
  wire [9:0] _seach_blockx_188_map_block;
  wire [9:0] _seach_blockx_188_now;
  wire [9:0] _seach_blockx_188_start;
  wire [9:0] _seach_blockx_188_goal;
  wire [9:0] _seach_blockx_188_data_out;
  wire _seach_blockx_188_in_do;
  wire _seach_blockx_188_p_reset;
  wire _seach_blockx_188_m_clock;
  wire [9:0] _seach_blockx_187_map_block;
  wire [9:0] _seach_blockx_187_now;
  wire [9:0] _seach_blockx_187_start;
  wire [9:0] _seach_blockx_187_goal;
  wire [9:0] _seach_blockx_187_data_out;
  wire _seach_blockx_187_in_do;
  wire _seach_blockx_187_p_reset;
  wire _seach_blockx_187_m_clock;
  wire [9:0] _seach_blockx_186_map_block;
  wire [9:0] _seach_blockx_186_now;
  wire [9:0] _seach_blockx_186_start;
  wire [9:0] _seach_blockx_186_goal;
  wire [9:0] _seach_blockx_186_data_out;
  wire _seach_blockx_186_in_do;
  wire _seach_blockx_186_p_reset;
  wire _seach_blockx_186_m_clock;
  wire [9:0] _seach_blockx_185_map_block;
  wire [9:0] _seach_blockx_185_now;
  wire [9:0] _seach_blockx_185_start;
  wire [9:0] _seach_blockx_185_goal;
  wire [9:0] _seach_blockx_185_data_out;
  wire _seach_blockx_185_in_do;
  wire _seach_blockx_185_p_reset;
  wire _seach_blockx_185_m_clock;
  wire [9:0] _seach_blockx_184_map_block;
  wire [9:0] _seach_blockx_184_now;
  wire [9:0] _seach_blockx_184_start;
  wire [9:0] _seach_blockx_184_goal;
  wire [9:0] _seach_blockx_184_data_out;
  wire _seach_blockx_184_in_do;
  wire _seach_blockx_184_p_reset;
  wire _seach_blockx_184_m_clock;
  wire [9:0] _seach_blockx_183_map_block;
  wire [9:0] _seach_blockx_183_now;
  wire [9:0] _seach_blockx_183_start;
  wire [9:0] _seach_blockx_183_goal;
  wire [9:0] _seach_blockx_183_data_out;
  wire _seach_blockx_183_in_do;
  wire _seach_blockx_183_p_reset;
  wire _seach_blockx_183_m_clock;
  wire [9:0] _seach_blockx_182_map_block;
  wire [9:0] _seach_blockx_182_now;
  wire [9:0] _seach_blockx_182_start;
  wire [9:0] _seach_blockx_182_goal;
  wire [9:0] _seach_blockx_182_data_out;
  wire _seach_blockx_182_in_do;
  wire _seach_blockx_182_p_reset;
  wire _seach_blockx_182_m_clock;
  wire [9:0] _seach_blockx_181_map_block;
  wire [9:0] _seach_blockx_181_now;
  wire [9:0] _seach_blockx_181_start;
  wire [9:0] _seach_blockx_181_goal;
  wire [9:0] _seach_blockx_181_data_out;
  wire _seach_blockx_181_in_do;
  wire _seach_blockx_181_p_reset;
  wire _seach_blockx_181_m_clock;
  wire [9:0] _seach_blockx_180_map_block;
  wire [9:0] _seach_blockx_180_now;
  wire [9:0] _seach_blockx_180_start;
  wire [9:0] _seach_blockx_180_goal;
  wire [9:0] _seach_blockx_180_data_out;
  wire _seach_blockx_180_in_do;
  wire _seach_blockx_180_p_reset;
  wire _seach_blockx_180_m_clock;
  wire [9:0] _seach_blockx_179_map_block;
  wire [9:0] _seach_blockx_179_now;
  wire [9:0] _seach_blockx_179_start;
  wire [9:0] _seach_blockx_179_goal;
  wire [9:0] _seach_blockx_179_data_out;
  wire _seach_blockx_179_in_do;
  wire _seach_blockx_179_p_reset;
  wire _seach_blockx_179_m_clock;
  wire [9:0] _seach_blockx_178_map_block;
  wire [9:0] _seach_blockx_178_now;
  wire [9:0] _seach_blockx_178_start;
  wire [9:0] _seach_blockx_178_goal;
  wire [9:0] _seach_blockx_178_data_out;
  wire _seach_blockx_178_in_do;
  wire _seach_blockx_178_p_reset;
  wire _seach_blockx_178_m_clock;
  wire [9:0] _seach_blockx_177_map_block;
  wire [9:0] _seach_blockx_177_now;
  wire [9:0] _seach_blockx_177_start;
  wire [9:0] _seach_blockx_177_goal;
  wire [9:0] _seach_blockx_177_data_out;
  wire _seach_blockx_177_in_do;
  wire _seach_blockx_177_p_reset;
  wire _seach_blockx_177_m_clock;
  wire [9:0] _seach_blockx_176_map_block;
  wire [9:0] _seach_blockx_176_now;
  wire [9:0] _seach_blockx_176_start;
  wire [9:0] _seach_blockx_176_goal;
  wire [9:0] _seach_blockx_176_data_out;
  wire _seach_blockx_176_in_do;
  wire _seach_blockx_176_p_reset;
  wire _seach_blockx_176_m_clock;
  wire [9:0] _seach_blockx_175_map_block;
  wire [9:0] _seach_blockx_175_now;
  wire [9:0] _seach_blockx_175_start;
  wire [9:0] _seach_blockx_175_goal;
  wire [9:0] _seach_blockx_175_data_out;
  wire _seach_blockx_175_in_do;
  wire _seach_blockx_175_p_reset;
  wire _seach_blockx_175_m_clock;
  wire [9:0] _seach_blockx_174_map_block;
  wire [9:0] _seach_blockx_174_now;
  wire [9:0] _seach_blockx_174_start;
  wire [9:0] _seach_blockx_174_goal;
  wire [9:0] _seach_blockx_174_data_out;
  wire _seach_blockx_174_in_do;
  wire _seach_blockx_174_p_reset;
  wire _seach_blockx_174_m_clock;
  wire [9:0] _seach_blockx_173_map_block;
  wire [9:0] _seach_blockx_173_now;
  wire [9:0] _seach_blockx_173_start;
  wire [9:0] _seach_blockx_173_goal;
  wire [9:0] _seach_blockx_173_data_out;
  wire _seach_blockx_173_in_do;
  wire _seach_blockx_173_p_reset;
  wire _seach_blockx_173_m_clock;
  wire [9:0] _seach_blockx_172_map_block;
  wire [9:0] _seach_blockx_172_now;
  wire [9:0] _seach_blockx_172_start;
  wire [9:0] _seach_blockx_172_goal;
  wire [9:0] _seach_blockx_172_data_out;
  wire _seach_blockx_172_in_do;
  wire _seach_blockx_172_p_reset;
  wire _seach_blockx_172_m_clock;
  wire [9:0] _seach_blockx_171_map_block;
  wire [9:0] _seach_blockx_171_now;
  wire [9:0] _seach_blockx_171_start;
  wire [9:0] _seach_blockx_171_goal;
  wire [9:0] _seach_blockx_171_data_out;
  wire _seach_blockx_171_in_do;
  wire _seach_blockx_171_p_reset;
  wire _seach_blockx_171_m_clock;
  wire [9:0] _seach_blockx_170_map_block;
  wire [9:0] _seach_blockx_170_now;
  wire [9:0] _seach_blockx_170_start;
  wire [9:0] _seach_blockx_170_goal;
  wire [9:0] _seach_blockx_170_data_out;
  wire _seach_blockx_170_in_do;
  wire _seach_blockx_170_p_reset;
  wire _seach_blockx_170_m_clock;
  wire [9:0] _seach_blockx_169_map_block;
  wire [9:0] _seach_blockx_169_now;
  wire [9:0] _seach_blockx_169_start;
  wire [9:0] _seach_blockx_169_goal;
  wire [9:0] _seach_blockx_169_data_out;
  wire _seach_blockx_169_in_do;
  wire _seach_blockx_169_p_reset;
  wire _seach_blockx_169_m_clock;
  wire [9:0] _seach_blockx_168_map_block;
  wire [9:0] _seach_blockx_168_now;
  wire [9:0] _seach_blockx_168_start;
  wire [9:0] _seach_blockx_168_goal;
  wire [9:0] _seach_blockx_168_data_out;
  wire _seach_blockx_168_in_do;
  wire _seach_blockx_168_p_reset;
  wire _seach_blockx_168_m_clock;
  wire [9:0] _seach_blockx_167_map_block;
  wire [9:0] _seach_blockx_167_now;
  wire [9:0] _seach_blockx_167_start;
  wire [9:0] _seach_blockx_167_goal;
  wire [9:0] _seach_blockx_167_data_out;
  wire _seach_blockx_167_in_do;
  wire _seach_blockx_167_p_reset;
  wire _seach_blockx_167_m_clock;
  wire [9:0] _seach_blockx_166_map_block;
  wire [9:0] _seach_blockx_166_now;
  wire [9:0] _seach_blockx_166_start;
  wire [9:0] _seach_blockx_166_goal;
  wire [9:0] _seach_blockx_166_data_out;
  wire _seach_blockx_166_in_do;
  wire _seach_blockx_166_p_reset;
  wire _seach_blockx_166_m_clock;
  wire [9:0] _seach_blockx_165_map_block;
  wire [9:0] _seach_blockx_165_now;
  wire [9:0] _seach_blockx_165_start;
  wire [9:0] _seach_blockx_165_goal;
  wire [9:0] _seach_blockx_165_data_out;
  wire _seach_blockx_165_in_do;
  wire _seach_blockx_165_p_reset;
  wire _seach_blockx_165_m_clock;
  wire [9:0] _seach_blockx_164_map_block;
  wire [9:0] _seach_blockx_164_now;
  wire [9:0] _seach_blockx_164_start;
  wire [9:0] _seach_blockx_164_goal;
  wire [9:0] _seach_blockx_164_data_out;
  wire _seach_blockx_164_in_do;
  wire _seach_blockx_164_p_reset;
  wire _seach_blockx_164_m_clock;
  wire [9:0] _seach_blockx_163_map_block;
  wire [9:0] _seach_blockx_163_now;
  wire [9:0] _seach_blockx_163_start;
  wire [9:0] _seach_blockx_163_goal;
  wire [9:0] _seach_blockx_163_data_out;
  wire _seach_blockx_163_in_do;
  wire _seach_blockx_163_p_reset;
  wire _seach_blockx_163_m_clock;
  wire [9:0] _seach_blockx_162_map_block;
  wire [9:0] _seach_blockx_162_now;
  wire [9:0] _seach_blockx_162_start;
  wire [9:0] _seach_blockx_162_goal;
  wire [9:0] _seach_blockx_162_data_out;
  wire _seach_blockx_162_in_do;
  wire _seach_blockx_162_p_reset;
  wire _seach_blockx_162_m_clock;
  wire [9:0] _seach_blockx_161_map_block;
  wire [9:0] _seach_blockx_161_now;
  wire [9:0] _seach_blockx_161_start;
  wire [9:0] _seach_blockx_161_goal;
  wire [9:0] _seach_blockx_161_data_out;
  wire _seach_blockx_161_in_do;
  wire _seach_blockx_161_p_reset;
  wire _seach_blockx_161_m_clock;
  wire [9:0] _seach_blockx_160_map_block;
  wire [9:0] _seach_blockx_160_now;
  wire [9:0] _seach_blockx_160_start;
  wire [9:0] _seach_blockx_160_goal;
  wire [9:0] _seach_blockx_160_data_out;
  wire _seach_blockx_160_in_do;
  wire _seach_blockx_160_p_reset;
  wire _seach_blockx_160_m_clock;
  wire [9:0] _seach_blockx_159_map_block;
  wire [9:0] _seach_blockx_159_now;
  wire [9:0] _seach_blockx_159_start;
  wire [9:0] _seach_blockx_159_goal;
  wire [9:0] _seach_blockx_159_data_out;
  wire _seach_blockx_159_in_do;
  wire _seach_blockx_159_p_reset;
  wire _seach_blockx_159_m_clock;
  wire [9:0] _seach_blockx_158_map_block;
  wire [9:0] _seach_blockx_158_now;
  wire [9:0] _seach_blockx_158_start;
  wire [9:0] _seach_blockx_158_goal;
  wire [9:0] _seach_blockx_158_data_out;
  wire _seach_blockx_158_in_do;
  wire _seach_blockx_158_p_reset;
  wire _seach_blockx_158_m_clock;
  wire [9:0] _seach_blockx_157_map_block;
  wire [9:0] _seach_blockx_157_now;
  wire [9:0] _seach_blockx_157_start;
  wire [9:0] _seach_blockx_157_goal;
  wire [9:0] _seach_blockx_157_data_out;
  wire _seach_blockx_157_in_do;
  wire _seach_blockx_157_p_reset;
  wire _seach_blockx_157_m_clock;
  wire [9:0] _seach_blockx_156_map_block;
  wire [9:0] _seach_blockx_156_now;
  wire [9:0] _seach_blockx_156_start;
  wire [9:0] _seach_blockx_156_goal;
  wire [9:0] _seach_blockx_156_data_out;
  wire _seach_blockx_156_in_do;
  wire _seach_blockx_156_p_reset;
  wire _seach_blockx_156_m_clock;
  wire [9:0] _seach_blockx_155_map_block;
  wire [9:0] _seach_blockx_155_now;
  wire [9:0] _seach_blockx_155_start;
  wire [9:0] _seach_blockx_155_goal;
  wire [9:0] _seach_blockx_155_data_out;
  wire _seach_blockx_155_in_do;
  wire _seach_blockx_155_p_reset;
  wire _seach_blockx_155_m_clock;
  wire [9:0] _seach_blockx_154_map_block;
  wire [9:0] _seach_blockx_154_now;
  wire [9:0] _seach_blockx_154_start;
  wire [9:0] _seach_blockx_154_goal;
  wire [9:0] _seach_blockx_154_data_out;
  wire _seach_blockx_154_in_do;
  wire _seach_blockx_154_p_reset;
  wire _seach_blockx_154_m_clock;
  wire [9:0] _seach_blockx_153_map_block;
  wire [9:0] _seach_blockx_153_now;
  wire [9:0] _seach_blockx_153_start;
  wire [9:0] _seach_blockx_153_goal;
  wire [9:0] _seach_blockx_153_data_out;
  wire _seach_blockx_153_in_do;
  wire _seach_blockx_153_p_reset;
  wire _seach_blockx_153_m_clock;
  wire [9:0] _seach_blockx_152_map_block;
  wire [9:0] _seach_blockx_152_now;
  wire [9:0] _seach_blockx_152_start;
  wire [9:0] _seach_blockx_152_goal;
  wire [9:0] _seach_blockx_152_data_out;
  wire _seach_blockx_152_in_do;
  wire _seach_blockx_152_p_reset;
  wire _seach_blockx_152_m_clock;
  wire [9:0] _seach_blockx_151_map_block;
  wire [9:0] _seach_blockx_151_now;
  wire [9:0] _seach_blockx_151_start;
  wire [9:0] _seach_blockx_151_goal;
  wire [9:0] _seach_blockx_151_data_out;
  wire _seach_blockx_151_in_do;
  wire _seach_blockx_151_p_reset;
  wire _seach_blockx_151_m_clock;
  wire [9:0] _seach_blockx_150_map_block;
  wire [9:0] _seach_blockx_150_now;
  wire [9:0] _seach_blockx_150_start;
  wire [9:0] _seach_blockx_150_goal;
  wire [9:0] _seach_blockx_150_data_out;
  wire _seach_blockx_150_in_do;
  wire _seach_blockx_150_p_reset;
  wire _seach_blockx_150_m_clock;
  wire [9:0] _seach_blockx_149_map_block;
  wire [9:0] _seach_blockx_149_now;
  wire [9:0] _seach_blockx_149_start;
  wire [9:0] _seach_blockx_149_goal;
  wire [9:0] _seach_blockx_149_data_out;
  wire _seach_blockx_149_in_do;
  wire _seach_blockx_149_p_reset;
  wire _seach_blockx_149_m_clock;
  wire [9:0] _seach_blockx_148_map_block;
  wire [9:0] _seach_blockx_148_now;
  wire [9:0] _seach_blockx_148_start;
  wire [9:0] _seach_blockx_148_goal;
  wire [9:0] _seach_blockx_148_data_out;
  wire _seach_blockx_148_in_do;
  wire _seach_blockx_148_p_reset;
  wire _seach_blockx_148_m_clock;
  wire [9:0] _seach_blockx_147_map_block;
  wire [9:0] _seach_blockx_147_now;
  wire [9:0] _seach_blockx_147_start;
  wire [9:0] _seach_blockx_147_goal;
  wire [9:0] _seach_blockx_147_data_out;
  wire _seach_blockx_147_in_do;
  wire _seach_blockx_147_p_reset;
  wire _seach_blockx_147_m_clock;
  wire [9:0] _seach_blockx_146_map_block;
  wire [9:0] _seach_blockx_146_now;
  wire [9:0] _seach_blockx_146_start;
  wire [9:0] _seach_blockx_146_goal;
  wire [9:0] _seach_blockx_146_data_out;
  wire _seach_blockx_146_in_do;
  wire _seach_blockx_146_p_reset;
  wire _seach_blockx_146_m_clock;
  wire [9:0] _seach_blockx_145_map_block;
  wire [9:0] _seach_blockx_145_now;
  wire [9:0] _seach_blockx_145_start;
  wire [9:0] _seach_blockx_145_goal;
  wire [9:0] _seach_blockx_145_data_out;
  wire _seach_blockx_145_in_do;
  wire _seach_blockx_145_p_reset;
  wire _seach_blockx_145_m_clock;
  wire [9:0] _seach_blockx_144_map_block;
  wire [9:0] _seach_blockx_144_now;
  wire [9:0] _seach_blockx_144_start;
  wire [9:0] _seach_blockx_144_goal;
  wire [9:0] _seach_blockx_144_data_out;
  wire _seach_blockx_144_in_do;
  wire _seach_blockx_144_p_reset;
  wire _seach_blockx_144_m_clock;
  wire [9:0] _seach_blockx_143_map_block;
  wire [9:0] _seach_blockx_143_now;
  wire [9:0] _seach_blockx_143_start;
  wire [9:0] _seach_blockx_143_goal;
  wire [9:0] _seach_blockx_143_data_out;
  wire _seach_blockx_143_in_do;
  wire _seach_blockx_143_p_reset;
  wire _seach_blockx_143_m_clock;
  wire [9:0] _seach_blockx_142_map_block;
  wire [9:0] _seach_blockx_142_now;
  wire [9:0] _seach_blockx_142_start;
  wire [9:0] _seach_blockx_142_goal;
  wire [9:0] _seach_blockx_142_data_out;
  wire _seach_blockx_142_in_do;
  wire _seach_blockx_142_p_reset;
  wire _seach_blockx_142_m_clock;
  wire [9:0] _seach_blockx_141_map_block;
  wire [9:0] _seach_blockx_141_now;
  wire [9:0] _seach_blockx_141_start;
  wire [9:0] _seach_blockx_141_goal;
  wire [9:0] _seach_blockx_141_data_out;
  wire _seach_blockx_141_in_do;
  wire _seach_blockx_141_p_reset;
  wire _seach_blockx_141_m_clock;
  wire [9:0] _seach_blockx_140_map_block;
  wire [9:0] _seach_blockx_140_now;
  wire [9:0] _seach_blockx_140_start;
  wire [9:0] _seach_blockx_140_goal;
  wire [9:0] _seach_blockx_140_data_out;
  wire _seach_blockx_140_in_do;
  wire _seach_blockx_140_p_reset;
  wire _seach_blockx_140_m_clock;
  wire [9:0] _seach_blockx_139_map_block;
  wire [9:0] _seach_blockx_139_now;
  wire [9:0] _seach_blockx_139_start;
  wire [9:0] _seach_blockx_139_goal;
  wire [9:0] _seach_blockx_139_data_out;
  wire _seach_blockx_139_in_do;
  wire _seach_blockx_139_p_reset;
  wire _seach_blockx_139_m_clock;
  wire [9:0] _seach_blockx_138_map_block;
  wire [9:0] _seach_blockx_138_now;
  wire [9:0] _seach_blockx_138_start;
  wire [9:0] _seach_blockx_138_goal;
  wire [9:0] _seach_blockx_138_data_out;
  wire _seach_blockx_138_in_do;
  wire _seach_blockx_138_p_reset;
  wire _seach_blockx_138_m_clock;
  wire [9:0] _seach_blockx_137_map_block;
  wire [9:0] _seach_blockx_137_now;
  wire [9:0] _seach_blockx_137_start;
  wire [9:0] _seach_blockx_137_goal;
  wire [9:0] _seach_blockx_137_data_out;
  wire _seach_blockx_137_in_do;
  wire _seach_blockx_137_p_reset;
  wire _seach_blockx_137_m_clock;
  wire [9:0] _seach_blockx_136_map_block;
  wire [9:0] _seach_blockx_136_now;
  wire [9:0] _seach_blockx_136_start;
  wire [9:0] _seach_blockx_136_goal;
  wire [9:0] _seach_blockx_136_data_out;
  wire _seach_blockx_136_in_do;
  wire _seach_blockx_136_p_reset;
  wire _seach_blockx_136_m_clock;
  wire [9:0] _seach_blockx_135_map_block;
  wire [9:0] _seach_blockx_135_now;
  wire [9:0] _seach_blockx_135_start;
  wire [9:0] _seach_blockx_135_goal;
  wire [9:0] _seach_blockx_135_data_out;
  wire _seach_blockx_135_in_do;
  wire _seach_blockx_135_p_reset;
  wire _seach_blockx_135_m_clock;
  wire [9:0] _seach_blockx_134_map_block;
  wire [9:0] _seach_blockx_134_now;
  wire [9:0] _seach_blockx_134_start;
  wire [9:0] _seach_blockx_134_goal;
  wire [9:0] _seach_blockx_134_data_out;
  wire _seach_blockx_134_in_do;
  wire _seach_blockx_134_p_reset;
  wire _seach_blockx_134_m_clock;
  wire [9:0] _seach_blockx_133_map_block;
  wire [9:0] _seach_blockx_133_now;
  wire [9:0] _seach_blockx_133_start;
  wire [9:0] _seach_blockx_133_goal;
  wire [9:0] _seach_blockx_133_data_out;
  wire _seach_blockx_133_in_do;
  wire _seach_blockx_133_p_reset;
  wire _seach_blockx_133_m_clock;
  wire [9:0] _seach_blockx_132_map_block;
  wire [9:0] _seach_blockx_132_now;
  wire [9:0] _seach_blockx_132_start;
  wire [9:0] _seach_blockx_132_goal;
  wire [9:0] _seach_blockx_132_data_out;
  wire _seach_blockx_132_in_do;
  wire _seach_blockx_132_p_reset;
  wire _seach_blockx_132_m_clock;
  wire [9:0] _seach_blockx_131_map_block;
  wire [9:0] _seach_blockx_131_now;
  wire [9:0] _seach_blockx_131_start;
  wire [9:0] _seach_blockx_131_goal;
  wire [9:0] _seach_blockx_131_data_out;
  wire _seach_blockx_131_in_do;
  wire _seach_blockx_131_p_reset;
  wire _seach_blockx_131_m_clock;
  wire [9:0] _seach_blockx_130_map_block;
  wire [9:0] _seach_blockx_130_now;
  wire [9:0] _seach_blockx_130_start;
  wire [9:0] _seach_blockx_130_goal;
  wire [9:0] _seach_blockx_130_data_out;
  wire _seach_blockx_130_in_do;
  wire _seach_blockx_130_p_reset;
  wire _seach_blockx_130_m_clock;
  wire [9:0] _seach_blockx_129_map_block;
  wire [9:0] _seach_blockx_129_now;
  wire [9:0] _seach_blockx_129_start;
  wire [9:0] _seach_blockx_129_goal;
  wire [9:0] _seach_blockx_129_data_out;
  wire _seach_blockx_129_in_do;
  wire _seach_blockx_129_p_reset;
  wire _seach_blockx_129_m_clock;
  wire [9:0] _seach_blockx_128_map_block;
  wire [9:0] _seach_blockx_128_now;
  wire [9:0] _seach_blockx_128_start;
  wire [9:0] _seach_blockx_128_goal;
  wire [9:0] _seach_blockx_128_data_out;
  wire _seach_blockx_128_in_do;
  wire _seach_blockx_128_p_reset;
  wire _seach_blockx_128_m_clock;
  wire [9:0] _seach_blockx_127_map_block;
  wire [9:0] _seach_blockx_127_now;
  wire [9:0] _seach_blockx_127_start;
  wire [9:0] _seach_blockx_127_goal;
  wire [9:0] _seach_blockx_127_data_out;
  wire _seach_blockx_127_in_do;
  wire _seach_blockx_127_p_reset;
  wire _seach_blockx_127_m_clock;
  wire [9:0] _seach_blockx_126_map_block;
  wire [9:0] _seach_blockx_126_now;
  wire [9:0] _seach_blockx_126_start;
  wire [9:0] _seach_blockx_126_goal;
  wire [9:0] _seach_blockx_126_data_out;
  wire _seach_blockx_126_in_do;
  wire _seach_blockx_126_p_reset;
  wire _seach_blockx_126_m_clock;
  wire [9:0] _seach_blockx_125_map_block;
  wire [9:0] _seach_blockx_125_now;
  wire [9:0] _seach_blockx_125_start;
  wire [9:0] _seach_blockx_125_goal;
  wire [9:0] _seach_blockx_125_data_out;
  wire _seach_blockx_125_in_do;
  wire _seach_blockx_125_p_reset;
  wire _seach_blockx_125_m_clock;
  wire [9:0] _seach_blockx_124_map_block;
  wire [9:0] _seach_blockx_124_now;
  wire [9:0] _seach_blockx_124_start;
  wire [9:0] _seach_blockx_124_goal;
  wire [9:0] _seach_blockx_124_data_out;
  wire _seach_blockx_124_in_do;
  wire _seach_blockx_124_p_reset;
  wire _seach_blockx_124_m_clock;
  wire [9:0] _seach_blockx_123_map_block;
  wire [9:0] _seach_blockx_123_now;
  wire [9:0] _seach_blockx_123_start;
  wire [9:0] _seach_blockx_123_goal;
  wire [9:0] _seach_blockx_123_data_out;
  wire _seach_blockx_123_in_do;
  wire _seach_blockx_123_p_reset;
  wire _seach_blockx_123_m_clock;
  wire [9:0] _seach_blockx_122_map_block;
  wire [9:0] _seach_blockx_122_now;
  wire [9:0] _seach_blockx_122_start;
  wire [9:0] _seach_blockx_122_goal;
  wire [9:0] _seach_blockx_122_data_out;
  wire _seach_blockx_122_in_do;
  wire _seach_blockx_122_p_reset;
  wire _seach_blockx_122_m_clock;
  wire [9:0] _seach_blockx_121_map_block;
  wire [9:0] _seach_blockx_121_now;
  wire [9:0] _seach_blockx_121_start;
  wire [9:0] _seach_blockx_121_goal;
  wire [9:0] _seach_blockx_121_data_out;
  wire _seach_blockx_121_in_do;
  wire _seach_blockx_121_p_reset;
  wire _seach_blockx_121_m_clock;
  wire [9:0] _seach_blockx_120_map_block;
  wire [9:0] _seach_blockx_120_now;
  wire [9:0] _seach_blockx_120_start;
  wire [9:0] _seach_blockx_120_goal;
  wire [9:0] _seach_blockx_120_data_out;
  wire _seach_blockx_120_in_do;
  wire _seach_blockx_120_p_reset;
  wire _seach_blockx_120_m_clock;
  wire [9:0] _seach_blockx_119_map_block;
  wire [9:0] _seach_blockx_119_now;
  wire [9:0] _seach_blockx_119_start;
  wire [9:0] _seach_blockx_119_goal;
  wire [9:0] _seach_blockx_119_data_out;
  wire _seach_blockx_119_in_do;
  wire _seach_blockx_119_p_reset;
  wire _seach_blockx_119_m_clock;
  wire [9:0] _seach_blockx_118_map_block;
  wire [9:0] _seach_blockx_118_now;
  wire [9:0] _seach_blockx_118_start;
  wire [9:0] _seach_blockx_118_goal;
  wire [9:0] _seach_blockx_118_data_out;
  wire _seach_blockx_118_in_do;
  wire _seach_blockx_118_p_reset;
  wire _seach_blockx_118_m_clock;
  wire [9:0] _seach_blockx_117_map_block;
  wire [9:0] _seach_blockx_117_now;
  wire [9:0] _seach_blockx_117_start;
  wire [9:0] _seach_blockx_117_goal;
  wire [9:0] _seach_blockx_117_data_out;
  wire _seach_blockx_117_in_do;
  wire _seach_blockx_117_p_reset;
  wire _seach_blockx_117_m_clock;
  wire [9:0] _seach_blockx_116_map_block;
  wire [9:0] _seach_blockx_116_now;
  wire [9:0] _seach_blockx_116_start;
  wire [9:0] _seach_blockx_116_goal;
  wire [9:0] _seach_blockx_116_data_out;
  wire _seach_blockx_116_in_do;
  wire _seach_blockx_116_p_reset;
  wire _seach_blockx_116_m_clock;
  wire [9:0] _seach_blockx_115_map_block;
  wire [9:0] _seach_blockx_115_now;
  wire [9:0] _seach_blockx_115_start;
  wire [9:0] _seach_blockx_115_goal;
  wire [9:0] _seach_blockx_115_data_out;
  wire _seach_blockx_115_in_do;
  wire _seach_blockx_115_p_reset;
  wire _seach_blockx_115_m_clock;
  wire [9:0] _seach_blockx_114_map_block;
  wire [9:0] _seach_blockx_114_now;
  wire [9:0] _seach_blockx_114_start;
  wire [9:0] _seach_blockx_114_goal;
  wire [9:0] _seach_blockx_114_data_out;
  wire _seach_blockx_114_in_do;
  wire _seach_blockx_114_p_reset;
  wire _seach_blockx_114_m_clock;
  wire [9:0] _seach_blockx_113_map_block;
  wire [9:0] _seach_blockx_113_now;
  wire [9:0] _seach_blockx_113_start;
  wire [9:0] _seach_blockx_113_goal;
  wire [9:0] _seach_blockx_113_data_out;
  wire _seach_blockx_113_in_do;
  wire _seach_blockx_113_p_reset;
  wire _seach_blockx_113_m_clock;
  wire [9:0] _seach_blockx_112_map_block;
  wire [9:0] _seach_blockx_112_now;
  wire [9:0] _seach_blockx_112_start;
  wire [9:0] _seach_blockx_112_goal;
  wire [9:0] _seach_blockx_112_data_out;
  wire _seach_blockx_112_in_do;
  wire _seach_blockx_112_p_reset;
  wire _seach_blockx_112_m_clock;
  wire [9:0] _seach_blockx_111_map_block;
  wire [9:0] _seach_blockx_111_now;
  wire [9:0] _seach_blockx_111_start;
  wire [9:0] _seach_blockx_111_goal;
  wire [9:0] _seach_blockx_111_data_out;
  wire _seach_blockx_111_in_do;
  wire _seach_blockx_111_p_reset;
  wire _seach_blockx_111_m_clock;
  wire [9:0] _seach_blockx_110_map_block;
  wire [9:0] _seach_blockx_110_now;
  wire [9:0] _seach_blockx_110_start;
  wire [9:0] _seach_blockx_110_goal;
  wire [9:0] _seach_blockx_110_data_out;
  wire _seach_blockx_110_in_do;
  wire _seach_blockx_110_p_reset;
  wire _seach_blockx_110_m_clock;
  wire [9:0] _seach_blockx_109_map_block;
  wire [9:0] _seach_blockx_109_now;
  wire [9:0] _seach_blockx_109_start;
  wire [9:0] _seach_blockx_109_goal;
  wire [9:0] _seach_blockx_109_data_out;
  wire _seach_blockx_109_in_do;
  wire _seach_blockx_109_p_reset;
  wire _seach_blockx_109_m_clock;
  wire [9:0] _seach_blockx_108_map_block;
  wire [9:0] _seach_blockx_108_now;
  wire [9:0] _seach_blockx_108_start;
  wire [9:0] _seach_blockx_108_goal;
  wire [9:0] _seach_blockx_108_data_out;
  wire _seach_blockx_108_in_do;
  wire _seach_blockx_108_p_reset;
  wire _seach_blockx_108_m_clock;
  wire [9:0] _seach_blockx_107_map_block;
  wire [9:0] _seach_blockx_107_now;
  wire [9:0] _seach_blockx_107_start;
  wire [9:0] _seach_blockx_107_goal;
  wire [9:0] _seach_blockx_107_data_out;
  wire _seach_blockx_107_in_do;
  wire _seach_blockx_107_p_reset;
  wire _seach_blockx_107_m_clock;
  wire [9:0] _seach_blockx_106_map_block;
  wire [9:0] _seach_blockx_106_now;
  wire [9:0] _seach_blockx_106_start;
  wire [9:0] _seach_blockx_106_goal;
  wire [9:0] _seach_blockx_106_data_out;
  wire _seach_blockx_106_in_do;
  wire _seach_blockx_106_p_reset;
  wire _seach_blockx_106_m_clock;
  wire [9:0] _seach_blockx_105_map_block;
  wire [9:0] _seach_blockx_105_now;
  wire [9:0] _seach_blockx_105_start;
  wire [9:0] _seach_blockx_105_goal;
  wire [9:0] _seach_blockx_105_data_out;
  wire _seach_blockx_105_in_do;
  wire _seach_blockx_105_p_reset;
  wire _seach_blockx_105_m_clock;
  wire [9:0] _seach_blockx_104_map_block;
  wire [9:0] _seach_blockx_104_now;
  wire [9:0] _seach_blockx_104_start;
  wire [9:0] _seach_blockx_104_goal;
  wire [9:0] _seach_blockx_104_data_out;
  wire _seach_blockx_104_in_do;
  wire _seach_blockx_104_p_reset;
  wire _seach_blockx_104_m_clock;
  wire [9:0] _seach_blockx_103_map_block;
  wire [9:0] _seach_blockx_103_now;
  wire [9:0] _seach_blockx_103_start;
  wire [9:0] _seach_blockx_103_goal;
  wire [9:0] _seach_blockx_103_data_out;
  wire _seach_blockx_103_in_do;
  wire _seach_blockx_103_p_reset;
  wire _seach_blockx_103_m_clock;
  wire [9:0] _seach_blockx_102_map_block;
  wire [9:0] _seach_blockx_102_now;
  wire [9:0] _seach_blockx_102_start;
  wire [9:0] _seach_blockx_102_goal;
  wire [9:0] _seach_blockx_102_data_out;
  wire _seach_blockx_102_in_do;
  wire _seach_blockx_102_p_reset;
  wire _seach_blockx_102_m_clock;
  wire [9:0] _seach_blockx_101_map_block;
  wire [9:0] _seach_blockx_101_now;
  wire [9:0] _seach_blockx_101_start;
  wire [9:0] _seach_blockx_101_goal;
  wire [9:0] _seach_blockx_101_data_out;
  wire _seach_blockx_101_in_do;
  wire _seach_blockx_101_p_reset;
  wire _seach_blockx_101_m_clock;
  wire [9:0] _seach_blockx_100_map_block;
  wire [9:0] _seach_blockx_100_now;
  wire [9:0] _seach_blockx_100_start;
  wire [9:0] _seach_blockx_100_goal;
  wire [9:0] _seach_blockx_100_data_out;
  wire _seach_blockx_100_in_do;
  wire _seach_blockx_100_p_reset;
  wire _seach_blockx_100_m_clock;
  wire [9:0] _seach_blockx_99_map_block;
  wire [9:0] _seach_blockx_99_now;
  wire [9:0] _seach_blockx_99_start;
  wire [9:0] _seach_blockx_99_goal;
  wire [9:0] _seach_blockx_99_data_out;
  wire _seach_blockx_99_in_do;
  wire _seach_blockx_99_p_reset;
  wire _seach_blockx_99_m_clock;
  wire [9:0] _seach_blockx_98_map_block;
  wire [9:0] _seach_blockx_98_now;
  wire [9:0] _seach_blockx_98_start;
  wire [9:0] _seach_blockx_98_goal;
  wire [9:0] _seach_blockx_98_data_out;
  wire _seach_blockx_98_in_do;
  wire _seach_blockx_98_p_reset;
  wire _seach_blockx_98_m_clock;
  wire [9:0] _seach_blockx_97_map_block;
  wire [9:0] _seach_blockx_97_now;
  wire [9:0] _seach_blockx_97_start;
  wire [9:0] _seach_blockx_97_goal;
  wire [9:0] _seach_blockx_97_data_out;
  wire _seach_blockx_97_in_do;
  wire _seach_blockx_97_p_reset;
  wire _seach_blockx_97_m_clock;
  wire [9:0] _seach_blockx_96_map_block;
  wire [9:0] _seach_blockx_96_now;
  wire [9:0] _seach_blockx_96_start;
  wire [9:0] _seach_blockx_96_goal;
  wire [9:0] _seach_blockx_96_data_out;
  wire _seach_blockx_96_in_do;
  wire _seach_blockx_96_p_reset;
  wire _seach_blockx_96_m_clock;
  wire [9:0] _seach_blockx_95_map_block;
  wire [9:0] _seach_blockx_95_now;
  wire [9:0] _seach_blockx_95_start;
  wire [9:0] _seach_blockx_95_goal;
  wire [9:0] _seach_blockx_95_data_out;
  wire _seach_blockx_95_in_do;
  wire _seach_blockx_95_p_reset;
  wire _seach_blockx_95_m_clock;
  wire [9:0] _seach_blockx_94_map_block;
  wire [9:0] _seach_blockx_94_now;
  wire [9:0] _seach_blockx_94_start;
  wire [9:0] _seach_blockx_94_goal;
  wire [9:0] _seach_blockx_94_data_out;
  wire _seach_blockx_94_in_do;
  wire _seach_blockx_94_p_reset;
  wire _seach_blockx_94_m_clock;
  wire [9:0] _seach_blockx_93_map_block;
  wire [9:0] _seach_blockx_93_now;
  wire [9:0] _seach_blockx_93_start;
  wire [9:0] _seach_blockx_93_goal;
  wire [9:0] _seach_blockx_93_data_out;
  wire _seach_blockx_93_in_do;
  wire _seach_blockx_93_p_reset;
  wire _seach_blockx_93_m_clock;
  wire [9:0] _seach_blockx_92_map_block;
  wire [9:0] _seach_blockx_92_now;
  wire [9:0] _seach_blockx_92_start;
  wire [9:0] _seach_blockx_92_goal;
  wire [9:0] _seach_blockx_92_data_out;
  wire _seach_blockx_92_in_do;
  wire _seach_blockx_92_p_reset;
  wire _seach_blockx_92_m_clock;
  wire [9:0] _seach_blockx_91_map_block;
  wire [9:0] _seach_blockx_91_now;
  wire [9:0] _seach_blockx_91_start;
  wire [9:0] _seach_blockx_91_goal;
  wire [9:0] _seach_blockx_91_data_out;
  wire _seach_blockx_91_in_do;
  wire _seach_blockx_91_p_reset;
  wire _seach_blockx_91_m_clock;
  wire [9:0] _seach_blockx_90_map_block;
  wire [9:0] _seach_blockx_90_now;
  wire [9:0] _seach_blockx_90_start;
  wire [9:0] _seach_blockx_90_goal;
  wire [9:0] _seach_blockx_90_data_out;
  wire _seach_blockx_90_in_do;
  wire _seach_blockx_90_p_reset;
  wire _seach_blockx_90_m_clock;
  wire [9:0] _seach_blockx_89_map_block;
  wire [9:0] _seach_blockx_89_now;
  wire [9:0] _seach_blockx_89_start;
  wire [9:0] _seach_blockx_89_goal;
  wire [9:0] _seach_blockx_89_data_out;
  wire _seach_blockx_89_in_do;
  wire _seach_blockx_89_p_reset;
  wire _seach_blockx_89_m_clock;
  wire [9:0] _seach_blockx_88_map_block;
  wire [9:0] _seach_blockx_88_now;
  wire [9:0] _seach_blockx_88_start;
  wire [9:0] _seach_blockx_88_goal;
  wire [9:0] _seach_blockx_88_data_out;
  wire _seach_blockx_88_in_do;
  wire _seach_blockx_88_p_reset;
  wire _seach_blockx_88_m_clock;
  wire [9:0] _seach_blockx_87_map_block;
  wire [9:0] _seach_blockx_87_now;
  wire [9:0] _seach_blockx_87_start;
  wire [9:0] _seach_blockx_87_goal;
  wire [9:0] _seach_blockx_87_data_out;
  wire _seach_blockx_87_in_do;
  wire _seach_blockx_87_p_reset;
  wire _seach_blockx_87_m_clock;
  wire [9:0] _seach_blockx_86_map_block;
  wire [9:0] _seach_blockx_86_now;
  wire [9:0] _seach_blockx_86_start;
  wire [9:0] _seach_blockx_86_goal;
  wire [9:0] _seach_blockx_86_data_out;
  wire _seach_blockx_86_in_do;
  wire _seach_blockx_86_p_reset;
  wire _seach_blockx_86_m_clock;
  wire [9:0] _seach_blockx_85_map_block;
  wire [9:0] _seach_blockx_85_now;
  wire [9:0] _seach_blockx_85_start;
  wire [9:0] _seach_blockx_85_goal;
  wire [9:0] _seach_blockx_85_data_out;
  wire _seach_blockx_85_in_do;
  wire _seach_blockx_85_p_reset;
  wire _seach_blockx_85_m_clock;
  wire [9:0] _seach_blockx_84_map_block;
  wire [9:0] _seach_blockx_84_now;
  wire [9:0] _seach_blockx_84_start;
  wire [9:0] _seach_blockx_84_goal;
  wire [9:0] _seach_blockx_84_data_out;
  wire _seach_blockx_84_in_do;
  wire _seach_blockx_84_p_reset;
  wire _seach_blockx_84_m_clock;
  wire [9:0] _seach_blockx_83_map_block;
  wire [9:0] _seach_blockx_83_now;
  wire [9:0] _seach_blockx_83_start;
  wire [9:0] _seach_blockx_83_goal;
  wire [9:0] _seach_blockx_83_data_out;
  wire _seach_blockx_83_in_do;
  wire _seach_blockx_83_p_reset;
  wire _seach_blockx_83_m_clock;
  wire [9:0] _seach_blockx_82_map_block;
  wire [9:0] _seach_blockx_82_now;
  wire [9:0] _seach_blockx_82_start;
  wire [9:0] _seach_blockx_82_goal;
  wire [9:0] _seach_blockx_82_data_out;
  wire _seach_blockx_82_in_do;
  wire _seach_blockx_82_p_reset;
  wire _seach_blockx_82_m_clock;
  wire [9:0] _seach_blockx_81_map_block;
  wire [9:0] _seach_blockx_81_now;
  wire [9:0] _seach_blockx_81_start;
  wire [9:0] _seach_blockx_81_goal;
  wire [9:0] _seach_blockx_81_data_out;
  wire _seach_blockx_81_in_do;
  wire _seach_blockx_81_p_reset;
  wire _seach_blockx_81_m_clock;
  wire [9:0] _seach_blockx_80_map_block;
  wire [9:0] _seach_blockx_80_now;
  wire [9:0] _seach_blockx_80_start;
  wire [9:0] _seach_blockx_80_goal;
  wire [9:0] _seach_blockx_80_data_out;
  wire _seach_blockx_80_in_do;
  wire _seach_blockx_80_p_reset;
  wire _seach_blockx_80_m_clock;
  wire [9:0] _seach_blockx_79_map_block;
  wire [9:0] _seach_blockx_79_now;
  wire [9:0] _seach_blockx_79_start;
  wire [9:0] _seach_blockx_79_goal;
  wire [9:0] _seach_blockx_79_data_out;
  wire _seach_blockx_79_in_do;
  wire _seach_blockx_79_p_reset;
  wire _seach_blockx_79_m_clock;
  wire [9:0] _seach_blockx_78_map_block;
  wire [9:0] _seach_blockx_78_now;
  wire [9:0] _seach_blockx_78_start;
  wire [9:0] _seach_blockx_78_goal;
  wire [9:0] _seach_blockx_78_data_out;
  wire _seach_blockx_78_in_do;
  wire _seach_blockx_78_p_reset;
  wire _seach_blockx_78_m_clock;
  wire [9:0] _seach_blockx_77_map_block;
  wire [9:0] _seach_blockx_77_now;
  wire [9:0] _seach_blockx_77_start;
  wire [9:0] _seach_blockx_77_goal;
  wire [9:0] _seach_blockx_77_data_out;
  wire _seach_blockx_77_in_do;
  wire _seach_blockx_77_p_reset;
  wire _seach_blockx_77_m_clock;
  wire [9:0] _seach_blockx_76_map_block;
  wire [9:0] _seach_blockx_76_now;
  wire [9:0] _seach_blockx_76_start;
  wire [9:0] _seach_blockx_76_goal;
  wire [9:0] _seach_blockx_76_data_out;
  wire _seach_blockx_76_in_do;
  wire _seach_blockx_76_p_reset;
  wire _seach_blockx_76_m_clock;
  wire [9:0] _seach_blockx_75_map_block;
  wire [9:0] _seach_blockx_75_now;
  wire [9:0] _seach_blockx_75_start;
  wire [9:0] _seach_blockx_75_goal;
  wire [9:0] _seach_blockx_75_data_out;
  wire _seach_blockx_75_in_do;
  wire _seach_blockx_75_p_reset;
  wire _seach_blockx_75_m_clock;
  wire [9:0] _seach_blockx_74_map_block;
  wire [9:0] _seach_blockx_74_now;
  wire [9:0] _seach_blockx_74_start;
  wire [9:0] _seach_blockx_74_goal;
  wire [9:0] _seach_blockx_74_data_out;
  wire _seach_blockx_74_in_do;
  wire _seach_blockx_74_p_reset;
  wire _seach_blockx_74_m_clock;
  wire [9:0] _seach_blockx_73_map_block;
  wire [9:0] _seach_blockx_73_now;
  wire [9:0] _seach_blockx_73_start;
  wire [9:0] _seach_blockx_73_goal;
  wire [9:0] _seach_blockx_73_data_out;
  wire _seach_blockx_73_in_do;
  wire _seach_blockx_73_p_reset;
  wire _seach_blockx_73_m_clock;
  wire [9:0] _seach_blockx_72_map_block;
  wire [9:0] _seach_blockx_72_now;
  wire [9:0] _seach_blockx_72_start;
  wire [9:0] _seach_blockx_72_goal;
  wire [9:0] _seach_blockx_72_data_out;
  wire _seach_blockx_72_in_do;
  wire _seach_blockx_72_p_reset;
  wire _seach_blockx_72_m_clock;
  wire [9:0] _seach_blockx_71_map_block;
  wire [9:0] _seach_blockx_71_now;
  wire [9:0] _seach_blockx_71_start;
  wire [9:0] _seach_blockx_71_goal;
  wire [9:0] _seach_blockx_71_data_out;
  wire _seach_blockx_71_in_do;
  wire _seach_blockx_71_p_reset;
  wire _seach_blockx_71_m_clock;
  wire [9:0] _seach_blockx_70_map_block;
  wire [9:0] _seach_blockx_70_now;
  wire [9:0] _seach_blockx_70_start;
  wire [9:0] _seach_blockx_70_goal;
  wire [9:0] _seach_blockx_70_data_out;
  wire _seach_blockx_70_in_do;
  wire _seach_blockx_70_p_reset;
  wire _seach_blockx_70_m_clock;
  wire [9:0] _seach_blockx_69_map_block;
  wire [9:0] _seach_blockx_69_now;
  wire [9:0] _seach_blockx_69_start;
  wire [9:0] _seach_blockx_69_goal;
  wire [9:0] _seach_blockx_69_data_out;
  wire _seach_blockx_69_in_do;
  wire _seach_blockx_69_p_reset;
  wire _seach_blockx_69_m_clock;
  wire [9:0] _seach_blockx_68_map_block;
  wire [9:0] _seach_blockx_68_now;
  wire [9:0] _seach_blockx_68_start;
  wire [9:0] _seach_blockx_68_goal;
  wire [9:0] _seach_blockx_68_data_out;
  wire _seach_blockx_68_in_do;
  wire _seach_blockx_68_p_reset;
  wire _seach_blockx_68_m_clock;
  wire [9:0] _seach_blockx_67_map_block;
  wire [9:0] _seach_blockx_67_now;
  wire [9:0] _seach_blockx_67_start;
  wire [9:0] _seach_blockx_67_goal;
  wire [9:0] _seach_blockx_67_data_out;
  wire _seach_blockx_67_in_do;
  wire _seach_blockx_67_p_reset;
  wire _seach_blockx_67_m_clock;
  wire [9:0] _seach_blockx_66_map_block;
  wire [9:0] _seach_blockx_66_now;
  wire [9:0] _seach_blockx_66_start;
  wire [9:0] _seach_blockx_66_goal;
  wire [9:0] _seach_blockx_66_data_out;
  wire _seach_blockx_66_in_do;
  wire _seach_blockx_66_p_reset;
  wire _seach_blockx_66_m_clock;
  wire [9:0] _seach_blockx_65_map_block;
  wire [9:0] _seach_blockx_65_now;
  wire [9:0] _seach_blockx_65_start;
  wire [9:0] _seach_blockx_65_goal;
  wire [9:0] _seach_blockx_65_data_out;
  wire _seach_blockx_65_in_do;
  wire _seach_blockx_65_p_reset;
  wire _seach_blockx_65_m_clock;
  wire [9:0] _seach_blockx_64_map_block;
  wire [9:0] _seach_blockx_64_now;
  wire [9:0] _seach_blockx_64_start;
  wire [9:0] _seach_blockx_64_goal;
  wire [9:0] _seach_blockx_64_data_out;
  wire _seach_blockx_64_in_do;
  wire _seach_blockx_64_p_reset;
  wire _seach_blockx_64_m_clock;
  wire [9:0] _seach_blockx_63_map_block;
  wire [9:0] _seach_blockx_63_now;
  wire [9:0] _seach_blockx_63_start;
  wire [9:0] _seach_blockx_63_goal;
  wire [9:0] _seach_blockx_63_data_out;
  wire _seach_blockx_63_in_do;
  wire _seach_blockx_63_p_reset;
  wire _seach_blockx_63_m_clock;
  wire [9:0] _seach_blockx_62_map_block;
  wire [9:0] _seach_blockx_62_now;
  wire [9:0] _seach_blockx_62_start;
  wire [9:0] _seach_blockx_62_goal;
  wire [9:0] _seach_blockx_62_data_out;
  wire _seach_blockx_62_in_do;
  wire _seach_blockx_62_p_reset;
  wire _seach_blockx_62_m_clock;
  wire [9:0] _seach_blockx_61_map_block;
  wire [9:0] _seach_blockx_61_now;
  wire [9:0] _seach_blockx_61_start;
  wire [9:0] _seach_blockx_61_goal;
  wire [9:0] _seach_blockx_61_data_out;
  wire _seach_blockx_61_in_do;
  wire _seach_blockx_61_p_reset;
  wire _seach_blockx_61_m_clock;
  wire [9:0] _seach_blockx_60_map_block;
  wire [9:0] _seach_blockx_60_now;
  wire [9:0] _seach_blockx_60_start;
  wire [9:0] _seach_blockx_60_goal;
  wire [9:0] _seach_blockx_60_data_out;
  wire _seach_blockx_60_in_do;
  wire _seach_blockx_60_p_reset;
  wire _seach_blockx_60_m_clock;
  wire [9:0] _seach_blockx_59_map_block;
  wire [9:0] _seach_blockx_59_now;
  wire [9:0] _seach_blockx_59_start;
  wire [9:0] _seach_blockx_59_goal;
  wire [9:0] _seach_blockx_59_data_out;
  wire _seach_blockx_59_in_do;
  wire _seach_blockx_59_p_reset;
  wire _seach_blockx_59_m_clock;
  wire [9:0] _seach_blockx_58_map_block;
  wire [9:0] _seach_blockx_58_now;
  wire [9:0] _seach_blockx_58_start;
  wire [9:0] _seach_blockx_58_goal;
  wire [9:0] _seach_blockx_58_data_out;
  wire _seach_blockx_58_in_do;
  wire _seach_blockx_58_p_reset;
  wire _seach_blockx_58_m_clock;
  wire [9:0] _seach_blockx_57_map_block;
  wire [9:0] _seach_blockx_57_now;
  wire [9:0] _seach_blockx_57_start;
  wire [9:0] _seach_blockx_57_goal;
  wire [9:0] _seach_blockx_57_data_out;
  wire _seach_blockx_57_in_do;
  wire _seach_blockx_57_p_reset;
  wire _seach_blockx_57_m_clock;
  wire [9:0] _seach_blockx_56_map_block;
  wire [9:0] _seach_blockx_56_now;
  wire [9:0] _seach_blockx_56_start;
  wire [9:0] _seach_blockx_56_goal;
  wire [9:0] _seach_blockx_56_data_out;
  wire _seach_blockx_56_in_do;
  wire _seach_blockx_56_p_reset;
  wire _seach_blockx_56_m_clock;
  wire [9:0] _seach_blockx_55_map_block;
  wire [9:0] _seach_blockx_55_now;
  wire [9:0] _seach_blockx_55_start;
  wire [9:0] _seach_blockx_55_goal;
  wire [9:0] _seach_blockx_55_data_out;
  wire _seach_blockx_55_in_do;
  wire _seach_blockx_55_p_reset;
  wire _seach_blockx_55_m_clock;
  wire [9:0] _seach_blockx_54_map_block;
  wire [9:0] _seach_blockx_54_now;
  wire [9:0] _seach_blockx_54_start;
  wire [9:0] _seach_blockx_54_goal;
  wire [9:0] _seach_blockx_54_data_out;
  wire _seach_blockx_54_in_do;
  wire _seach_blockx_54_p_reset;
  wire _seach_blockx_54_m_clock;
  wire [9:0] _seach_blockx_53_map_block;
  wire [9:0] _seach_blockx_53_now;
  wire [9:0] _seach_blockx_53_start;
  wire [9:0] _seach_blockx_53_goal;
  wire [9:0] _seach_blockx_53_data_out;
  wire _seach_blockx_53_in_do;
  wire _seach_blockx_53_p_reset;
  wire _seach_blockx_53_m_clock;
  wire [9:0] _seach_blockx_52_map_block;
  wire [9:0] _seach_blockx_52_now;
  wire [9:0] _seach_blockx_52_start;
  wire [9:0] _seach_blockx_52_goal;
  wire [9:0] _seach_blockx_52_data_out;
  wire _seach_blockx_52_in_do;
  wire _seach_blockx_52_p_reset;
  wire _seach_blockx_52_m_clock;
  wire [9:0] _seach_blockx_51_map_block;
  wire [9:0] _seach_blockx_51_now;
  wire [9:0] _seach_blockx_51_start;
  wire [9:0] _seach_blockx_51_goal;
  wire [9:0] _seach_blockx_51_data_out;
  wire _seach_blockx_51_in_do;
  wire _seach_blockx_51_p_reset;
  wire _seach_blockx_51_m_clock;
  wire [9:0] _seach_blockx_50_map_block;
  wire [9:0] _seach_blockx_50_now;
  wire [9:0] _seach_blockx_50_start;
  wire [9:0] _seach_blockx_50_goal;
  wire [9:0] _seach_blockx_50_data_out;
  wire _seach_blockx_50_in_do;
  wire _seach_blockx_50_p_reset;
  wire _seach_blockx_50_m_clock;
  wire [9:0] _seach_blockx_49_map_block;
  wire [9:0] _seach_blockx_49_now;
  wire [9:0] _seach_blockx_49_start;
  wire [9:0] _seach_blockx_49_goal;
  wire [9:0] _seach_blockx_49_data_out;
  wire _seach_blockx_49_in_do;
  wire _seach_blockx_49_p_reset;
  wire _seach_blockx_49_m_clock;
  wire [9:0] _seach_blockx_48_map_block;
  wire [9:0] _seach_blockx_48_now;
  wire [9:0] _seach_blockx_48_start;
  wire [9:0] _seach_blockx_48_goal;
  wire [9:0] _seach_blockx_48_data_out;
  wire _seach_blockx_48_in_do;
  wire _seach_blockx_48_p_reset;
  wire _seach_blockx_48_m_clock;
  wire [9:0] _seach_blockx_47_map_block;
  wire [9:0] _seach_blockx_47_now;
  wire [9:0] _seach_blockx_47_start;
  wire [9:0] _seach_blockx_47_goal;
  wire [9:0] _seach_blockx_47_data_out;
  wire _seach_blockx_47_in_do;
  wire _seach_blockx_47_p_reset;
  wire _seach_blockx_47_m_clock;
  wire [9:0] _seach_blockx_46_map_block;
  wire [9:0] _seach_blockx_46_now;
  wire [9:0] _seach_blockx_46_start;
  wire [9:0] _seach_blockx_46_goal;
  wire [9:0] _seach_blockx_46_data_out;
  wire _seach_blockx_46_in_do;
  wire _seach_blockx_46_p_reset;
  wire _seach_blockx_46_m_clock;
  wire [9:0] _seach_blockx_45_map_block;
  wire [9:0] _seach_blockx_45_now;
  wire [9:0] _seach_blockx_45_start;
  wire [9:0] _seach_blockx_45_goal;
  wire [9:0] _seach_blockx_45_data_out;
  wire _seach_blockx_45_in_do;
  wire _seach_blockx_45_p_reset;
  wire _seach_blockx_45_m_clock;
  wire [9:0] _seach_blockx_44_map_block;
  wire [9:0] _seach_blockx_44_now;
  wire [9:0] _seach_blockx_44_start;
  wire [9:0] _seach_blockx_44_goal;
  wire [9:0] _seach_blockx_44_data_out;
  wire _seach_blockx_44_in_do;
  wire _seach_blockx_44_p_reset;
  wire _seach_blockx_44_m_clock;
  wire [9:0] _seach_blockx_43_map_block;
  wire [9:0] _seach_blockx_43_now;
  wire [9:0] _seach_blockx_43_start;
  wire [9:0] _seach_blockx_43_goal;
  wire [9:0] _seach_blockx_43_data_out;
  wire _seach_blockx_43_in_do;
  wire _seach_blockx_43_p_reset;
  wire _seach_blockx_43_m_clock;
  wire [9:0] _seach_blockx_42_map_block;
  wire [9:0] _seach_blockx_42_now;
  wire [9:0] _seach_blockx_42_start;
  wire [9:0] _seach_blockx_42_goal;
  wire [9:0] _seach_blockx_42_data_out;
  wire _seach_blockx_42_in_do;
  wire _seach_blockx_42_p_reset;
  wire _seach_blockx_42_m_clock;
  wire [9:0] _seach_blockx_41_map_block;
  wire [9:0] _seach_blockx_41_now;
  wire [9:0] _seach_blockx_41_start;
  wire [9:0] _seach_blockx_41_goal;
  wire [9:0] _seach_blockx_41_data_out;
  wire _seach_blockx_41_in_do;
  wire _seach_blockx_41_p_reset;
  wire _seach_blockx_41_m_clock;
  wire [9:0] _seach_blockx_40_map_block;
  wire [9:0] _seach_blockx_40_now;
  wire [9:0] _seach_blockx_40_start;
  wire [9:0] _seach_blockx_40_goal;
  wire [9:0] _seach_blockx_40_data_out;
  wire _seach_blockx_40_in_do;
  wire _seach_blockx_40_p_reset;
  wire _seach_blockx_40_m_clock;
  wire [9:0] _seach_blockx_39_map_block;
  wire [9:0] _seach_blockx_39_now;
  wire [9:0] _seach_blockx_39_start;
  wire [9:0] _seach_blockx_39_goal;
  wire [9:0] _seach_blockx_39_data_out;
  wire _seach_blockx_39_in_do;
  wire _seach_blockx_39_p_reset;
  wire _seach_blockx_39_m_clock;
  wire [9:0] _seach_blockx_38_map_block;
  wire [9:0] _seach_blockx_38_now;
  wire [9:0] _seach_blockx_38_start;
  wire [9:0] _seach_blockx_38_goal;
  wire [9:0] _seach_blockx_38_data_out;
  wire _seach_blockx_38_in_do;
  wire _seach_blockx_38_p_reset;
  wire _seach_blockx_38_m_clock;
  wire [9:0] _seach_blockx_37_map_block;
  wire [9:0] _seach_blockx_37_now;
  wire [9:0] _seach_blockx_37_start;
  wire [9:0] _seach_blockx_37_goal;
  wire [9:0] _seach_blockx_37_data_out;
  wire _seach_blockx_37_in_do;
  wire _seach_blockx_37_p_reset;
  wire _seach_blockx_37_m_clock;
  wire [9:0] _seach_blockx_36_map_block;
  wire [9:0] _seach_blockx_36_now;
  wire [9:0] _seach_blockx_36_start;
  wire [9:0] _seach_blockx_36_goal;
  wire [9:0] _seach_blockx_36_data_out;
  wire _seach_blockx_36_in_do;
  wire _seach_blockx_36_p_reset;
  wire _seach_blockx_36_m_clock;
  wire [9:0] _seach_blockx_35_map_block;
  wire [9:0] _seach_blockx_35_now;
  wire [9:0] _seach_blockx_35_start;
  wire [9:0] _seach_blockx_35_goal;
  wire [9:0] _seach_blockx_35_data_out;
  wire _seach_blockx_35_in_do;
  wire _seach_blockx_35_p_reset;
  wire _seach_blockx_35_m_clock;
  wire [9:0] _seach_blockx_34_map_block;
  wire [9:0] _seach_blockx_34_now;
  wire [9:0] _seach_blockx_34_start;
  wire [9:0] _seach_blockx_34_goal;
  wire [9:0] _seach_blockx_34_data_out;
  wire _seach_blockx_34_in_do;
  wire _seach_blockx_34_p_reset;
  wire _seach_blockx_34_m_clock;
  wire [9:0] _seach_blockx_33_map_block;
  wire [9:0] _seach_blockx_33_now;
  wire [9:0] _seach_blockx_33_start;
  wire [9:0] _seach_blockx_33_goal;
  wire [9:0] _seach_blockx_33_data_out;
  wire _seach_blockx_33_in_do;
  wire _seach_blockx_33_p_reset;
  wire _seach_blockx_33_m_clock;
  wire [9:0] _seach_blockx_32_map_block;
  wire [9:0] _seach_blockx_32_now;
  wire [9:0] _seach_blockx_32_start;
  wire [9:0] _seach_blockx_32_goal;
  wire [9:0] _seach_blockx_32_data_out;
  wire _seach_blockx_32_in_do;
  wire _seach_blockx_32_p_reset;
  wire _seach_blockx_32_m_clock;
  wire [9:0] _seach_blockx_31_map_block;
  wire [9:0] _seach_blockx_31_now;
  wire [9:0] _seach_blockx_31_start;
  wire [9:0] _seach_blockx_31_goal;
  wire [9:0] _seach_blockx_31_data_out;
  wire _seach_blockx_31_in_do;
  wire _seach_blockx_31_p_reset;
  wire _seach_blockx_31_m_clock;
  wire [9:0] _seach_blockx_30_map_block;
  wire [9:0] _seach_blockx_30_now;
  wire [9:0] _seach_blockx_30_start;
  wire [9:0] _seach_blockx_30_goal;
  wire [9:0] _seach_blockx_30_data_out;
  wire _seach_blockx_30_in_do;
  wire _seach_blockx_30_p_reset;
  wire _seach_blockx_30_m_clock;
  wire [9:0] _seach_blockx_29_map_block;
  wire [9:0] _seach_blockx_29_now;
  wire [9:0] _seach_blockx_29_start;
  wire [9:0] _seach_blockx_29_goal;
  wire [9:0] _seach_blockx_29_data_out;
  wire _seach_blockx_29_in_do;
  wire _seach_blockx_29_p_reset;
  wire _seach_blockx_29_m_clock;
  wire [9:0] _seach_blockx_28_map_block;
  wire [9:0] _seach_blockx_28_now;
  wire [9:0] _seach_blockx_28_start;
  wire [9:0] _seach_blockx_28_goal;
  wire [9:0] _seach_blockx_28_data_out;
  wire _seach_blockx_28_in_do;
  wire _seach_blockx_28_p_reset;
  wire _seach_blockx_28_m_clock;
  wire [9:0] _seach_blockx_27_map_block;
  wire [9:0] _seach_blockx_27_now;
  wire [9:0] _seach_blockx_27_start;
  wire [9:0] _seach_blockx_27_goal;
  wire [9:0] _seach_blockx_27_data_out;
  wire _seach_blockx_27_in_do;
  wire _seach_blockx_27_p_reset;
  wire _seach_blockx_27_m_clock;
  wire [9:0] _seach_blockx_26_map_block;
  wire [9:0] _seach_blockx_26_now;
  wire [9:0] _seach_blockx_26_start;
  wire [9:0] _seach_blockx_26_goal;
  wire [9:0] _seach_blockx_26_data_out;
  wire _seach_blockx_26_in_do;
  wire _seach_blockx_26_p_reset;
  wire _seach_blockx_26_m_clock;
  wire [9:0] _seach_blockx_25_map_block;
  wire [9:0] _seach_blockx_25_now;
  wire [9:0] _seach_blockx_25_start;
  wire [9:0] _seach_blockx_25_goal;
  wire [9:0] _seach_blockx_25_data_out;
  wire _seach_blockx_25_in_do;
  wire _seach_blockx_25_p_reset;
  wire _seach_blockx_25_m_clock;
  wire [9:0] _seach_blockx_24_map_block;
  wire [9:0] _seach_blockx_24_now;
  wire [9:0] _seach_blockx_24_start;
  wire [9:0] _seach_blockx_24_goal;
  wire [9:0] _seach_blockx_24_data_out;
  wire _seach_blockx_24_in_do;
  wire _seach_blockx_24_p_reset;
  wire _seach_blockx_24_m_clock;
  wire [9:0] _seach_blockx_23_map_block;
  wire [9:0] _seach_blockx_23_now;
  wire [9:0] _seach_blockx_23_start;
  wire [9:0] _seach_blockx_23_goal;
  wire [9:0] _seach_blockx_23_data_out;
  wire _seach_blockx_23_in_do;
  wire _seach_blockx_23_p_reset;
  wire _seach_blockx_23_m_clock;
  wire [9:0] _seach_blockx_22_map_block;
  wire [9:0] _seach_blockx_22_now;
  wire [9:0] _seach_blockx_22_start;
  wire [9:0] _seach_blockx_22_goal;
  wire [9:0] _seach_blockx_22_data_out;
  wire _seach_blockx_22_in_do;
  wire _seach_blockx_22_p_reset;
  wire _seach_blockx_22_m_clock;
  wire [9:0] _seach_blockx_21_map_block;
  wire [9:0] _seach_blockx_21_now;
  wire [9:0] _seach_blockx_21_start;
  wire [9:0] _seach_blockx_21_goal;
  wire [9:0] _seach_blockx_21_data_out;
  wire _seach_blockx_21_in_do;
  wire _seach_blockx_21_p_reset;
  wire _seach_blockx_21_m_clock;
  wire [9:0] _seach_blockx_20_map_block;
  wire [9:0] _seach_blockx_20_now;
  wire [9:0] _seach_blockx_20_start;
  wire [9:0] _seach_blockx_20_goal;
  wire [9:0] _seach_blockx_20_data_out;
  wire _seach_blockx_20_in_do;
  wire _seach_blockx_20_p_reset;
  wire _seach_blockx_20_m_clock;
  wire [9:0] _seach_blockx_19_map_block;
  wire [9:0] _seach_blockx_19_now;
  wire [9:0] _seach_blockx_19_start;
  wire [9:0] _seach_blockx_19_goal;
  wire [9:0] _seach_blockx_19_data_out;
  wire _seach_blockx_19_in_do;
  wire _seach_blockx_19_p_reset;
  wire _seach_blockx_19_m_clock;
  wire [9:0] _seach_blockx_18_map_block;
  wire [9:0] _seach_blockx_18_now;
  wire [9:0] _seach_blockx_18_start;
  wire [9:0] _seach_blockx_18_goal;
  wire [9:0] _seach_blockx_18_data_out;
  wire _seach_blockx_18_in_do;
  wire _seach_blockx_18_p_reset;
  wire _seach_blockx_18_m_clock;
  wire [9:0] _seach_blockx_17_map_block;
  wire [9:0] _seach_blockx_17_now;
  wire [9:0] _seach_blockx_17_start;
  wire [9:0] _seach_blockx_17_goal;
  wire [9:0] _seach_blockx_17_data_out;
  wire _seach_blockx_17_in_do;
  wire _seach_blockx_17_p_reset;
  wire _seach_blockx_17_m_clock;
  wire [9:0] _seach_blockx_16_map_block;
  wire [9:0] _seach_blockx_16_now;
  wire [9:0] _seach_blockx_16_start;
  wire [9:0] _seach_blockx_16_goal;
  wire [9:0] _seach_blockx_16_data_out;
  wire _seach_blockx_16_in_do;
  wire _seach_blockx_16_p_reset;
  wire _seach_blockx_16_m_clock;
  wire [9:0] _seach_blockx_15_map_block;
  wire [9:0] _seach_blockx_15_now;
  wire [9:0] _seach_blockx_15_start;
  wire [9:0] _seach_blockx_15_goal;
  wire [9:0] _seach_blockx_15_data_out;
  wire _seach_blockx_15_in_do;
  wire _seach_blockx_15_p_reset;
  wire _seach_blockx_15_m_clock;
  wire [9:0] _seach_blockx_14_map_block;
  wire [9:0] _seach_blockx_14_now;
  wire [9:0] _seach_blockx_14_start;
  wire [9:0] _seach_blockx_14_goal;
  wire [9:0] _seach_blockx_14_data_out;
  wire _seach_blockx_14_in_do;
  wire _seach_blockx_14_p_reset;
  wire _seach_blockx_14_m_clock;
  wire [9:0] _seach_blockx_13_map_block;
  wire [9:0] _seach_blockx_13_now;
  wire [9:0] _seach_blockx_13_start;
  wire [9:0] _seach_blockx_13_goal;
  wire [9:0] _seach_blockx_13_data_out;
  wire _seach_blockx_13_in_do;
  wire _seach_blockx_13_p_reset;
  wire _seach_blockx_13_m_clock;
  wire [9:0] _seach_blockx_12_map_block;
  wire [9:0] _seach_blockx_12_now;
  wire [9:0] _seach_blockx_12_start;
  wire [9:0] _seach_blockx_12_goal;
  wire [9:0] _seach_blockx_12_data_out;
  wire _seach_blockx_12_in_do;
  wire _seach_blockx_12_p_reset;
  wire _seach_blockx_12_m_clock;
  wire [9:0] _seach_blockx_11_map_block;
  wire [9:0] _seach_blockx_11_now;
  wire [9:0] _seach_blockx_11_start;
  wire [9:0] _seach_blockx_11_goal;
  wire [9:0] _seach_blockx_11_data_out;
  wire _seach_blockx_11_in_do;
  wire _seach_blockx_11_p_reset;
  wire _seach_blockx_11_m_clock;
  wire [9:0] _seach_blockx_10_map_block;
  wire [9:0] _seach_blockx_10_now;
  wire [9:0] _seach_blockx_10_start;
  wire [9:0] _seach_blockx_10_goal;
  wire [9:0] _seach_blockx_10_data_out;
  wire _seach_blockx_10_in_do;
  wire _seach_blockx_10_p_reset;
  wire _seach_blockx_10_m_clock;
  wire [9:0] _seach_blockx_9_map_block;
  wire [9:0] _seach_blockx_9_now;
  wire [9:0] _seach_blockx_9_start;
  wire [9:0] _seach_blockx_9_goal;
  wire [9:0] _seach_blockx_9_data_out;
  wire _seach_blockx_9_in_do;
  wire _seach_blockx_9_p_reset;
  wire _seach_blockx_9_m_clock;
  wire [9:0] _seach_blockx_8_map_block;
  wire [9:0] _seach_blockx_8_now;
  wire [9:0] _seach_blockx_8_start;
  wire [9:0] _seach_blockx_8_goal;
  wire [9:0] _seach_blockx_8_data_out;
  wire _seach_blockx_8_in_do;
  wire _seach_blockx_8_p_reset;
  wire _seach_blockx_8_m_clock;
  wire [9:0] _seach_blockx_7_map_block;
  wire [9:0] _seach_blockx_7_now;
  wire [9:0] _seach_blockx_7_start;
  wire [9:0] _seach_blockx_7_goal;
  wire [9:0] _seach_blockx_7_data_out;
  wire _seach_blockx_7_in_do;
  wire _seach_blockx_7_p_reset;
  wire _seach_blockx_7_m_clock;
  wire [9:0] _seach_blockx_6_map_block;
  wire [9:0] _seach_blockx_6_now;
  wire [9:0] _seach_blockx_6_start;
  wire [9:0] _seach_blockx_6_goal;
  wire [9:0] _seach_blockx_6_data_out;
  wire _seach_blockx_6_in_do;
  wire _seach_blockx_6_p_reset;
  wire _seach_blockx_6_m_clock;
  wire [9:0] _seach_blockx_5_map_block;
  wire [9:0] _seach_blockx_5_now;
  wire [9:0] _seach_blockx_5_start;
  wire [9:0] _seach_blockx_5_goal;
  wire [9:0] _seach_blockx_5_data_out;
  wire _seach_blockx_5_in_do;
  wire _seach_blockx_5_p_reset;
  wire _seach_blockx_5_m_clock;
  wire [9:0] _seach_blockx_4_map_block;
  wire [9:0] _seach_blockx_4_now;
  wire [9:0] _seach_blockx_4_start;
  wire [9:0] _seach_blockx_4_goal;
  wire [9:0] _seach_blockx_4_data_out;
  wire _seach_blockx_4_in_do;
  wire _seach_blockx_4_p_reset;
  wire _seach_blockx_4_m_clock;
  wire [9:0] _seach_blockx_3_map_block;
  wire [9:0] _seach_blockx_3_now;
  wire [9:0] _seach_blockx_3_start;
  wire [9:0] _seach_blockx_3_goal;
  wire [9:0] _seach_blockx_3_data_out;
  wire _seach_blockx_3_in_do;
  wire _seach_blockx_3_p_reset;
  wire _seach_blockx_3_m_clock;
  wire [9:0] _seach_blockx_2_map_block;
  wire [9:0] _seach_blockx_2_now;
  wire [9:0] _seach_blockx_2_start;
  wire [9:0] _seach_blockx_2_goal;
  wire [9:0] _seach_blockx_2_data_out;
  wire _seach_blockx_2_in_do;
  wire _seach_blockx_2_p_reset;
  wire _seach_blockx_2_m_clock;
  wire [9:0] _seach_blockx_1_map_block;
  wire [9:0] _seach_blockx_1_now;
  wire [9:0] _seach_blockx_1_start;
  wire [9:0] _seach_blockx_1_goal;
  wire [9:0] _seach_blockx_1_data_out;
  wire _seach_blockx_1_in_do;
  wire _seach_blockx_1_p_reset;
  wire _seach_blockx_1_m_clock;
  reg _reg_0;
  reg _reg_1;
  wire _net_2;
  wire _net_3;
  wire _net_4;
  wire _net_5;
  wire _net_6;
  wire _net_7;
  wire _net_8;
  wire _net_9;
  wire _net_10;
  wire _net_11;
  wire _net_12;
  wire _net_13;
  wire _net_14;
  wire _net_15;
  wire _net_16;
  wire _net_17;
  wire _net_18;
  wire _net_19;
  wire _net_20;
  wire _net_21;
  wire _net_22;
  wire _net_23;
  wire _net_24;
  wire _net_25;
  wire _net_26;
  wire _net_27;
  wire _net_28;
  wire _net_29;
  wire _net_30;
  wire _net_31;
  wire _net_32;
  wire _net_33;
  wire _net_34;
  wire _net_35;
  wire _net_36;
  wire _net_37;
  wire _net_38;
  wire _net_39;
  wire _net_40;
  wire _net_41;
  wire _net_42;
  wire _net_43;
  wire _net_44;
  wire _net_45;
  wire _net_46;
  wire _net_47;
  wire _net_48;
  wire _net_49;
  wire _net_50;
  wire _net_51;
  wire _net_52;
  wire _net_53;
  wire _net_54;
  wire _net_55;
  wire _net_56;
  wire _net_57;
  wire _net_58;
  wire _net_59;
  wire _net_60;
  wire _net_61;
  wire _net_62;
  wire _net_63;
  wire _net_64;
  wire _net_65;
  wire _net_66;
  wire _net_67;
  wire _net_68;
  wire _net_69;
  wire _net_70;
  wire _net_71;
  wire _net_72;
  wire _net_73;
  wire _net_74;
  wire _net_75;
  wire _net_76;
  wire _net_77;
  wire _net_78;
  wire _net_79;
  wire _net_80;
  wire _net_81;
  wire _net_82;
  wire _net_83;
  wire _net_84;
  wire _net_85;
  wire _net_86;
  wire _net_87;
  wire _net_88;
  wire _net_89;
  wire _net_90;
  wire _net_91;
  wire _net_92;
  wire _net_93;
  wire _net_94;
  wire _net_95;
  wire _net_96;
  wire _net_97;
  wire _net_98;
  wire _net_99;
  wire _net_100;
  wire _net_101;
  wire _net_102;
  wire _net_103;
  wire _net_104;
  wire _net_105;
  wire _net_106;
  wire _net_107;
  wire _net_108;
  wire _net_109;
  wire _net_110;
  wire _net_111;
  wire _net_112;
  wire _net_113;
  wire _net_114;
  wire _net_115;
  wire _net_116;
  wire _net_117;
  wire _net_118;
  wire _net_119;
  wire _net_120;
  wire _net_121;
  wire _net_122;
  wire _net_123;
  wire _net_124;
  wire _net_125;
  wire _net_126;
  wire _net_127;
  wire _net_128;
  wire _net_129;
  wire _net_130;
  wire _net_131;
  wire _net_132;
  wire _net_133;
  wire _net_134;
  wire _net_135;
  wire _net_136;
  wire _net_137;
  wire _net_138;
  wire _net_139;
  wire _net_140;
  wire _net_141;
  wire _net_142;
  wire _net_143;
  wire _net_144;
  wire _net_145;
  wire _net_146;
  wire _net_147;
  wire _net_148;
  wire _net_149;
  wire _net_150;
  wire _net_151;
  wire _net_152;
  wire _net_153;
  wire _net_154;
  wire _net_155;
  wire _net_156;
  wire _net_157;
  wire _net_158;
  wire _net_159;
  wire _net_160;
  wire _net_161;
  wire _net_162;
  wire _net_163;
  wire _net_164;
  wire _net_165;
  wire _net_166;
  wire _net_167;
  wire _net_168;
  wire _net_169;
  wire _net_170;
  wire _net_171;
  wire _net_172;
  wire _net_173;
  wire _net_174;
  wire _net_175;
  wire _net_176;
  wire _net_177;
  wire _net_178;
  wire _net_179;
  wire _net_180;
  wire _net_181;
  wire _net_182;
  wire _net_183;
  wire _net_184;
  wire _net_185;
  wire _net_186;
  wire _net_187;
  wire _net_188;
  wire _net_189;
  wire _net_190;
  wire _net_191;
  wire _net_192;
  wire _net_193;
  wire _net_194;
  wire _net_195;
  wire _net_196;
  wire _net_197;
  wire _net_198;
  wire _net_199;
  wire _net_200;
  wire _net_201;
  wire _net_202;
  wire _net_203;
  wire _net_204;
  wire _net_205;
  wire _net_206;
  wire _net_207;
  wire _net_208;
  wire _net_209;
  wire _net_210;
  wire _net_211;
  wire _net_212;
  wire _net_213;
  wire _net_214;
  wire _net_215;
  wire _net_216;
  wire _net_217;
  wire _net_218;
  wire _net_219;
  wire _net_220;
  wire _net_221;
  wire _net_222;
  wire _net_223;
  wire _net_224;
  wire _net_225;
  wire _net_226;
  wire _net_227;
  wire _net_228;
  wire _net_229;
  wire _net_230;
  wire _net_231;
  wire _net_232;
  wire _net_233;
  wire _net_234;
  wire _net_235;
  wire _net_236;
  wire _net_237;
  wire _net_238;
  wire _net_239;
  wire _net_240;
  wire _net_241;
  wire _net_242;
  wire _net_243;
  wire _net_244;
  wire _net_245;
  wire _net_246;
  wire _net_247;
  wire _net_248;
  wire _net_249;
  wire _net_250;
  wire _net_251;
  wire _net_252;
  wire _net_253;
  wire _net_254;
  wire _net_255;
  wire _net_256;
  wire _net_257;
  wire _net_258;
  wire _net_259;
  wire _net_260;
  wire _net_261;
  wire _net_262;
  wire _net_263;
  wire _net_264;
  wire _net_265;
  wire _net_266;
  wire _net_267;
  wire _net_268;
  wire _net_269;
  wire _net_270;
  wire _net_271;
  wire _net_272;
  wire _net_273;
  wire _net_274;
  wire _net_275;
  wire _net_276;
  wire _net_277;
  wire _net_278;
  wire _net_279;
  wire _net_280;
  wire _net_281;
  wire _net_282;
  wire _net_283;
  wire _net_284;
  wire _net_285;
  wire _net_286;
  wire _net_287;
  wire _net_288;
  wire _net_289;
  wire _net_290;
  wire _net_291;
  wire _net_292;
  wire _net_293;
  wire _net_294;
  wire _net_295;
  wire _net_296;
  wire _net_297;
  wire _net_298;
  wire _net_299;
  wire _net_300;
  wire _net_301;
  wire _net_302;
  wire _net_303;
  wire _net_304;
  wire _net_305;
  wire _net_306;
  wire _net_307;
  wire _net_308;
  wire _net_309;
  wire _net_310;
  wire _net_311;
  wire _net_312;
  wire _net_313;
  wire _net_314;
  wire _net_315;
  wire _net_316;
  wire _net_317;
  wire _net_318;
  wire _net_319;
  wire _net_320;
  wire _net_321;
  wire _net_322;
  wire _net_323;
  wire _net_324;
  wire _net_325;
  wire _net_326;
  wire _net_327;
  wire _net_328;
  wire _net_329;
  wire _net_330;
  wire _net_331;
  wire _net_332;
  wire _net_333;
  wire _net_334;
  wire _net_335;
  wire _net_336;
  wire _net_337;
  wire _net_338;
  wire _net_339;
  wire _net_340;
  wire _net_341;
  wire _net_342;
  wire _net_343;
  wire _net_344;
  wire _net_345;
  wire _net_346;
  wire _net_347;
  wire _net_348;
  wire _net_349;
  wire _net_350;
  wire _net_351;
  wire _net_352;
  wire _net_353;
  wire _net_354;
  wire _net_355;
  wire _net_356;
  wire _net_357;
  wire _net_358;
  wire _net_359;
  wire _net_360;
  wire _net_361;
  wire _net_362;
  wire _net_363;
  wire _net_364;
  wire _net_365;
  wire _net_366;
  wire _net_367;
  wire _net_368;
  wire _net_369;
  wire _net_370;
  wire _net_371;
  wire _net_372;
  wire _net_373;
  wire _net_374;
  wire _net_375;
  wire _net_376;
  wire _net_377;
  wire _net_378;
  wire _net_379;
  wire _net_380;
  wire _net_381;
  wire _net_382;
  wire _net_383;
  wire _net_384;
  wire _net_385;
  wire _net_386;
  wire _net_387;
  wire _net_388;
  wire _net_389;
  wire _net_390;
  wire _net_391;
  wire _net_392;
  wire _net_393;
  wire _net_394;
  wire _net_395;
  wire _net_396;
  wire _net_397;
  wire _net_398;
  wire _net_399;
  wire _net_400;
  wire _net_401;
  wire _net_402;
  wire _net_403;
  wire _net_404;
  wire _net_405;
  wire _net_406;
  wire _net_407;
  wire _net_408;
  wire _net_409;
  wire _net_410;
  wire _net_411;
  wire _net_412;
  wire _net_413;
  wire _net_414;
  wire _net_415;
  wire _net_416;
  wire _net_417;
  wire _net_418;
  wire _net_419;
  wire _net_420;
  wire _net_421;
  wire _net_422;
  wire _net_423;
  wire _net_424;
  wire _net_425;
  wire _net_426;
  wire _net_427;
  wire _net_428;
  wire _net_429;
  wire _net_430;
  wire _net_431;
  wire _net_432;
  wire _net_433;
  wire _net_434;
  wire _net_435;
  wire _net_436;
  wire _net_437;
  wire _net_438;
  wire _net_439;
  wire _net_440;
  wire _net_441;
  wire _net_442;
  wire _net_443;
  wire _net_444;
  wire _net_445;
  wire _net_446;
  wire _net_447;
  wire _net_448;
  wire _net_449;
  wire _net_450;
  wire _net_451;
  wire _net_452;
  wire _net_453;
  wire _net_454;
  wire _net_455;
  wire _net_456;
  wire _net_457;
  wire _net_458;
  wire _net_459;
  wire _net_460;
  wire _net_461;
  wire _net_462;
  wire _net_463;
  wire _net_464;
  wire _net_465;
  wire _net_466;
  wire _net_467;
  wire _net_468;
  wire _net_469;
  wire _net_470;
  wire _net_471;
  wire _net_472;
  wire _net_473;
  wire _net_474;
  wire _net_475;
  wire _net_476;
  wire _net_477;
  wire _net_478;
  wire _net_479;
  wire _net_480;
  wire _net_481;
  wire _net_482;
  wire _net_483;
  wire _net_484;
  wire _net_485;
  wire _net_486;
  wire _net_487;
  wire _net_488;
  wire _net_489;
  wire _net_490;
  wire _net_491;
  wire _net_492;
  wire _net_493;
  wire _net_494;
  wire _net_495;
  wire _net_496;
  wire _net_497;
  wire _net_498;
  wire _net_499;
  wire _net_500;
  wire _net_501;
  wire _net_502;
  wire _net_503;
  wire _net_504;
  wire _net_505;
  wire _net_506;
  wire _net_507;
  wire _net_508;
  wire _net_509;
  wire _net_510;
  wire _net_511;
  wire _net_512;
  wire _net_513;
  wire _net_514;
  wire _net_515;
  wire _net_516;
  wire _net_517;
  wire _net_518;
  wire _net_519;
  wire _net_520;
  wire _net_521;
  wire _net_522;
  wire _net_523;
  wire _net_524;
  wire _net_525;
  wire _net_526;
  wire _net_527;
  wire _net_528;
  wire _net_529;
  wire _net_530;
  wire _net_531;
  wire _net_532;
  wire _net_533;
  wire _net_534;
  wire _net_535;
  wire _net_536;
  wire _net_537;
  wire _net_538;
  wire _net_539;
  wire _net_540;
  wire _net_541;
  wire _net_542;
  wire _net_543;
  wire _net_544;
  wire _net_545;
  wire _net_546;
  wire _net_547;
  wire _net_548;
  wire _net_549;
  wire _net_550;
  wire _net_551;
  wire _net_552;
  wire _net_553;
  wire _net_554;
  wire _net_555;
  wire _net_556;
  wire _net_557;
  wire _net_558;
  wire _net_559;
  wire _net_560;
  wire _net_561;
  wire _net_562;
  wire _net_563;
  wire _net_564;
  wire _net_565;
  wire _net_566;
  wire _net_567;
  wire _net_568;
  wire _net_569;
  wire _net_570;
  wire _net_571;
  wire _net_572;
  wire _net_573;
  wire _net_574;
  wire _net_575;
  wire _net_576;
  wire _net_577;
  wire _net_578;
  wire _net_579;
  wire _net_580;
  wire _net_581;
  wire _net_582;
  wire _net_583;
  wire _net_584;
  wire _net_585;
  wire _net_586;
  wire _net_587;
  wire _net_588;
  wire _net_589;
  wire _net_590;
  wire _net_591;
  wire _net_592;
  wire _net_593;
  wire _net_594;
  wire _net_595;
  wire _net_596;
  wire _net_597;
  wire _net_598;
  wire _net_599;
  wire _net_600;
  wire _net_601;
  wire _net_602;
  wire _net_603;
  wire _net_604;
  wire _net_605;
  wire _net_606;
  wire _net_607;
  wire _net_608;
  wire _net_609;
  wire _net_610;
  wire _net_611;
  wire _net_612;
  wire _net_613;
  wire _net_614;
  wire _net_615;
  wire _net_616;
  wire _net_617;
  wire _net_618;
  wire _net_619;
  wire _net_620;
  wire _net_621;
  wire _net_622;
  wire _net_623;
  wire _net_624;
  wire _net_625;
  wire _net_626;
  wire _net_627;
  wire _net_628;
  wire _net_629;
  wire _net_630;
  wire _net_631;
  wire _net_632;
  wire _net_633;
  wire _net_634;
  wire _net_635;
  wire _net_636;
  wire _net_637;
  wire _net_638;
  wire _net_639;
  wire _net_640;
  wire _net_641;
  wire _net_642;
  wire _net_643;
  wire _net_644;
  wire _net_645;
  wire _net_646;
  wire _net_647;
  wire _net_648;
  wire _net_649;
  wire _net_650;
  wire _net_651;
  wire _net_652;
  wire _net_653;
  wire _net_654;
  wire _net_655;
  wire _net_656;
  wire _net_657;
  wire _net_658;
  wire _net_659;
  wire _net_660;
  wire _net_661;
  wire _net_662;
  wire _net_663;
  wire _net_664;
  wire _net_665;
  wire _net_666;
  wire _net_667;
  wire _net_668;
  wire _net_669;
  wire _net_670;
  wire _net_671;
  wire _net_672;
  wire _net_673;
  wire _net_674;
  wire _net_675;
  wire _net_676;
  wire _net_677;
  wire _net_678;
  wire _net_679;
  wire _net_680;
  wire _net_681;
  wire _net_682;
  wire _net_683;
  wire _net_684;
  wire _net_685;
  wire _net_686;
  wire _net_687;
  wire _net_688;
  wire _net_689;
  wire _net_690;
  wire _net_691;
  wire _net_692;
  wire _net_693;
  wire _net_694;
  wire _net_695;
  wire _net_696;
  wire _net_697;
  wire _net_698;
  wire _net_699;
  wire _net_700;
  wire _net_701;
  wire _net_702;
  wire _net_703;
  wire _net_704;
  wire _net_705;
  wire _net_706;
  wire _net_707;
  wire _net_708;
  wire _net_709;
  wire _net_710;
  wire _net_711;
  wire _net_712;
  wire _net_713;
  wire _net_714;
  wire _net_715;
  wire _net_716;
  wire _net_717;
  wire _net_718;
  wire _net_719;
  wire _net_720;
  wire _net_721;
  wire _net_722;
  wire _net_723;
  wire _net_724;
  wire _net_725;
  wire _net_726;
  wire _net_727;
  wire _net_728;
  wire _net_729;
  wire _net_730;
  wire _net_731;
  wire _net_732;
  wire _net_733;
  wire _net_734;
  wire _net_735;
  wire _net_736;
  wire _net_737;
  wire _net_738;
  wire _net_739;
  wire _net_740;
  wire _net_741;
  wire _net_742;
  wire _net_743;
  wire _net_744;
  wire _net_745;
  wire _net_746;
  wire _net_747;
  wire _net_748;
  wire _net_749;
  wire _net_750;
  wire _net_751;
  wire _net_752;
  wire _net_753;
  wire _net_754;
  wire _net_755;
  wire _net_756;
  wire _net_757;
  wire _net_758;
  wire _net_759;
  wire _net_760;
  wire _net_761;
  wire _net_762;
  wire _net_763;
  wire _net_764;
  wire _net_765;
  wire _net_766;
  wire _net_767;
  wire _net_768;
  wire _net_769;
  wire _net_770;
  wire _net_771;
  wire _net_772;
  wire _net_773;
  wire _net_774;
  wire _net_775;
  wire _net_776;
  wire _net_777;
  wire _net_778;
  wire _net_779;
  wire _net_780;
  wire _net_781;
  wire _net_782;
  wire _net_783;
  wire _net_784;
  wire _net_785;
  wire _net_786;
  wire _net_787;
  wire _net_788;
  wire _net_789;
  wire _net_790;
  wire _net_791;
  wire _net_792;
  wire _net_793;
  wire _net_794;
  wire _net_795;
  wire _net_796;
  wire _net_797;
  wire _net_798;
  wire _net_799;
  wire _net_800;
  wire _net_801;
  wire _net_802;
  wire _net_803;
  wire _net_804;
  wire _net_805;
  wire _net_806;
  wire _net_807;
  wire _net_808;
  wire _net_809;
  wire _net_810;
  wire _net_811;
  wire _net_812;
  wire _net_813;
  wire _net_814;
  wire _net_815;
  wire _net_816;
  wire _net_817;
  wire _net_818;
  wire _net_819;
  wire _net_820;
  wire _net_821;
  wire _net_822;
  wire _net_823;
  wire _net_824;
  wire _net_825;
  wire _net_826;
  wire _net_827;
  wire _net_828;
  wire _net_829;
  wire _net_830;
  wire _net_831;
  wire _net_832;
  wire _net_833;
  wire _net_834;
  wire _net_835;
  wire _net_836;
  wire _net_837;
  wire _net_838;
  wire _net_839;
  wire _net_840;
  wire _net_841;
  wire _net_842;
  wire _net_843;
  wire _net_844;
  wire _net_845;
  wire _net_846;
  wire _net_847;
  wire _net_848;
  wire _net_849;
  wire _net_850;
  wire _net_851;
  wire _net_852;
  wire _net_853;
  wire _net_854;
  wire _net_855;
  wire _net_856;
  wire _net_857;
  wire _net_858;
  wire _net_859;
  wire _net_860;
  wire _net_861;
  wire _net_862;
  wire _net_863;
  wire _net_864;
  wire _net_865;
  wire _net_866;
  wire _net_867;
  wire _net_868;
  wire _net_869;
  wire _net_870;
  wire _net_871;
  wire _net_872;
  wire _net_873;
  wire _net_874;
  wire _net_875;
  wire _net_876;
  wire _net_877;
  wire _net_878;
  wire _net_879;
  wire _net_880;
  wire _net_881;
  wire _net_882;
  wire _net_883;
  wire _net_884;
  wire _net_885;
  wire _net_886;
  wire _net_887;
  wire _net_888;
  wire _net_889;
  wire _net_890;
  wire _net_891;
  wire _net_892;
  wire _net_893;
  wire _net_894;
  wire _net_895;
  wire _net_896;
  wire _net_897;
  wire _net_898;
  wire _net_899;
  wire _net_900;
  wire _net_901;
  wire _net_902;
  wire _net_903;
  wire _net_904;
  wire _net_905;
  wire _net_906;
  wire _net_907;
  wire _net_908;
  wire _net_909;
  wire _net_910;
  wire _net_911;
  wire _net_912;
  wire _net_913;
  wire _net_914;
  wire _net_915;
  wire _net_916;
  wire _net_917;
  wire _net_918;
  wire _net_919;
  wire _net_920;
  wire _net_921;
  wire _net_922;
  wire _net_923;
  wire _net_924;
  wire _net_925;
  wire _net_926;
  wire _net_927;
  wire _net_928;
  wire _net_929;
  wire _net_930;
  wire _net_931;
  wire _net_932;
  wire _net_933;
  wire _net_934;
  wire _net_935;
  wire _net_936;
  wire _net_937;
  wire _net_938;
  wire _net_939;
  wire _net_940;
  wire _net_941;
  wire _net_942;
  wire _net_943;
  wire _net_944;
  wire _net_945;
  wire _net_946;
  wire _net_947;
  wire _net_948;
  wire _net_949;
  wire _net_950;
  wire _net_951;
  wire _net_952;
  wire _net_953;
  wire _net_954;
  wire _net_955;
  wire _net_956;
  wire _net_957;
  wire _net_958;
  wire _net_959;
  wire _net_960;
  wire _net_961;
  wire _net_962;
  wire _net_963;
  wire _net_964;
  wire _net_965;
  wire _net_966;
  wire _net_967;
  wire _net_968;
  wire _net_969;
  wire _net_970;
  wire _net_971;
  wire _net_972;
  wire _net_973;
  wire _net_974;
  wire _net_975;
  wire _net_976;
  wire _net_977;
  wire _net_978;
  wire _net_979;
  wire _net_980;
  wire _net_981;
  wire _net_982;
  wire _net_983;
  wire _net_984;
  wire _net_985;
  wire _net_986;
  wire _net_987;
  wire _net_988;
  wire _net_989;
  wire _net_990;
  wire _net_991;
  wire _net_992;
  wire _net_993;
  wire _net_994;
  wire _net_995;
  wire _net_996;
  wire _net_997;
  wire _net_998;
  wire _net_999;
  wire _net_1000;
  wire _net_1001;
  wire _net_1002;
  wire _net_1003;
  wire _net_1004;
  wire _net_1005;
  wire _net_1006;
  wire _net_1007;
  wire _net_1008;
  wire _net_1009;
  wire _net_1010;
  wire _net_1011;
  wire _net_1012;
  wire _net_1013;
  wire _net_1014;
  wire _net_1015;
  wire _net_1016;
  wire _net_1017;
  wire _net_1018;
  wire _net_1019;
  wire _net_1020;
  wire _net_1021;
  wire _net_1022;
  wire _net_1023;
  wire _net_1024;
  wire _net_1025;
  wire _net_1026;
  wire _net_1027;
  wire _net_1028;
  wire _net_1029;
  wire _net_1030;
  wire _net_1031;
  wire _net_1032;
  wire _net_1033;
  wire _net_1034;
  wire _net_1035;
  wire _net_1036;
  wire _net_1037;
  wire _net_1038;
  wire _net_1039;
  wire _net_1040;
  wire _net_1041;
  wire _net_1042;
  wire _net_1043;
  wire _net_1044;
  wire _net_1045;
  wire _net_1046;
  wire _net_1047;
  wire _net_1048;
  wire _net_1049;
  wire _net_1050;
  wire _net_1051;
  wire _net_1052;
  wire _net_1053;
  wire _net_1054;
  wire _net_1055;
  wire _net_1056;
  wire _net_1057;
  wire _net_1058;
  wire _net_1059;
  wire _net_1060;
  wire _net_1061;
  wire _net_1062;
  wire _net_1063;
  wire _net_1064;
  wire _net_1065;
  wire _net_1066;
  wire _net_1067;
  wire _net_1068;
  wire _net_1069;
  wire _net_1070;
  wire _net_1071;
  wire _net_1072;
  wire _net_1073;
  wire _net_1074;
  wire _net_1075;
  wire _net_1076;
  wire _net_1077;
  wire _net_1078;
  wire _net_1079;
  wire _net_1080;
  wire _net_1081;
  wire _net_1082;
  wire _net_1083;
  wire _net_1084;
  wire _net_1085;
  wire _net_1086;
  wire _net_1087;
  wire _net_1088;
  wire _net_1089;
  wire _net_1090;
  wire _net_1091;
  wire _net_1092;
  wire _net_1093;
  wire _net_1094;
  wire _net_1095;
  wire _net_1096;
  wire _net_1097;
  wire _net_1098;
  wire _net_1099;
  wire _net_1100;
  wire _net_1101;
  wire _net_1102;
  wire _net_1103;
  wire _net_1104;
  wire _net_1105;
  wire _net_1106;
  wire _net_1107;
  wire _net_1108;
  wire _net_1109;
  wire _net_1110;
  wire _net_1111;
  wire _net_1112;
  wire _net_1113;
  wire _net_1114;
  wire _net_1115;
  wire _net_1116;
  wire _net_1117;
  wire _net_1118;
  wire _net_1119;
  wire _net_1120;
  wire _net_1121;
  wire _net_1122;
  wire _net_1123;
  wire _net_1124;
  wire _net_1125;
  wire _net_1126;
  wire _net_1127;
  wire _net_1128;
  wire _net_1129;
  wire _net_1130;
  wire _net_1131;
  wire _net_1132;
  wire _net_1133;
  wire _net_1134;
  wire _net_1135;
  wire _net_1136;
  wire _net_1137;
  wire _net_1138;
  wire _net_1139;
  wire _net_1140;
  wire _net_1141;
  wire _net_1142;
  wire _net_1143;
  wire _net_1144;
  wire _net_1145;
  wire _net_1146;
  wire _net_1147;
  wire _net_1148;
  wire _net_1149;
  wire _net_1150;
  wire _net_1151;
  wire _net_1152;
  wire _net_1153;
  wire _net_1154;
  wire _net_1155;
  wire _net_1156;
  wire _net_1157;
  wire _net_1158;
  wire _net_1159;
  wire _net_1160;
  wire _net_1161;
  wire _net_1162;
  wire _net_1163;
  wire _net_1164;
  wire _net_1165;
  wire _net_1166;
  wire _net_1167;
  wire _net_1168;
  wire _net_1169;
  wire _net_1170;
  wire _net_1171;
  wire _net_1172;
  wire _net_1173;
  wire _net_1174;
  wire _net_1175;
  wire _net_1176;
  wire _net_1177;
  wire _net_1178;
  wire _net_1179;
  wire _net_1180;
  wire _net_1181;
  wire _net_1182;
  wire _net_1183;
  wire _net_1184;
  wire _net_1185;
  wire _net_1186;
  wire _net_1187;
  wire _net_1188;
  wire _net_1189;
  wire _net_1190;
  wire _net_1191;
  wire _net_1192;
  wire _net_1193;
  wire _net_1194;
  wire _net_1195;
  wire _net_1196;
  wire _net_1197;
  wire _net_1198;
  wire _net_1199;
  wire _net_1200;
  wire _net_1201;
  wire _net_1202;
  wire _net_1203;
  wire _net_1204;
  wire _net_1205;
  wire _net_1206;
  wire _net_1207;
  wire _net_1208;
  wire _net_1209;
  wire _net_1210;
  wire _net_1211;
  wire _net_1212;
  wire _net_1213;
  wire _net_1214;
  wire _net_1215;
  wire _net_1216;
  wire _net_1217;
  wire _net_1218;
  wire _net_1219;
  wire _net_1220;
  wire _net_1221;
  wire _net_1222;
  wire _net_1223;
  wire _net_1224;
  wire _net_1225;
  wire _net_1226;
  wire _net_1227;
  wire _net_1228;
  wire _net_1229;
  wire _net_1230;
  wire _net_1231;
  wire _net_1232;
  wire _net_1233;
  wire _net_1234;
  wire _net_1235;
  wire _net_1236;
  wire _net_1237;
  wire _net_1238;
  wire _net_1239;
  wire _net_1240;
  wire _net_1241;
  wire _net_1242;
  wire _net_1243;
  wire _net_1244;
  wire _net_1245;
  wire _net_1246;
  wire _net_1247;
  wire _net_1248;
  wire _net_1249;
  wire _net_1250;
  wire _net_1251;
  wire _net_1252;
  wire _net_1253;
  wire _net_1254;
  wire _net_1255;
  wire _net_1256;
  wire _net_1257;
  wire _net_1258;
  wire _net_1259;
  wire _net_1260;
  wire _net_1261;
  wire _net_1262;
  wire _net_1263;
  wire _net_1264;
seach_block seach_blockx (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_in_do), .start(_seach_blockx_start), .goal(_seach_blockx_goal), .data_out(_seach_blockx_data_out), .map_block(_seach_blockx_map_block), .now(_seach_blockx_now));
seach_block seach_blockx_419 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_419_in_do), .start(_seach_blockx_419_start), .goal(_seach_blockx_419_goal), .data_out(_seach_blockx_419_data_out), .map_block(_seach_blockx_419_map_block), .now(_seach_blockx_419_now));
seach_block seach_blockx_418 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_418_in_do), .start(_seach_blockx_418_start), .goal(_seach_blockx_418_goal), .data_out(_seach_blockx_418_data_out), .map_block(_seach_blockx_418_map_block), .now(_seach_blockx_418_now));
seach_block seach_blockx_417 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_417_in_do), .start(_seach_blockx_417_start), .goal(_seach_blockx_417_goal), .data_out(_seach_blockx_417_data_out), .map_block(_seach_blockx_417_map_block), .now(_seach_blockx_417_now));
seach_block seach_blockx_416 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_416_in_do), .start(_seach_blockx_416_start), .goal(_seach_blockx_416_goal), .data_out(_seach_blockx_416_data_out), .map_block(_seach_blockx_416_map_block), .now(_seach_blockx_416_now));
seach_block seach_blockx_415 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_415_in_do), .start(_seach_blockx_415_start), .goal(_seach_blockx_415_goal), .data_out(_seach_blockx_415_data_out), .map_block(_seach_blockx_415_map_block), .now(_seach_blockx_415_now));
seach_block seach_blockx_414 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_414_in_do), .start(_seach_blockx_414_start), .goal(_seach_blockx_414_goal), .data_out(_seach_blockx_414_data_out), .map_block(_seach_blockx_414_map_block), .now(_seach_blockx_414_now));
seach_block seach_blockx_413 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_413_in_do), .start(_seach_blockx_413_start), .goal(_seach_blockx_413_goal), .data_out(_seach_blockx_413_data_out), .map_block(_seach_blockx_413_map_block), .now(_seach_blockx_413_now));
seach_block seach_blockx_412 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_412_in_do), .start(_seach_blockx_412_start), .goal(_seach_blockx_412_goal), .data_out(_seach_blockx_412_data_out), .map_block(_seach_blockx_412_map_block), .now(_seach_blockx_412_now));
seach_block seach_blockx_411 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_411_in_do), .start(_seach_blockx_411_start), .goal(_seach_blockx_411_goal), .data_out(_seach_blockx_411_data_out), .map_block(_seach_blockx_411_map_block), .now(_seach_blockx_411_now));
seach_block seach_blockx_410 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_410_in_do), .start(_seach_blockx_410_start), .goal(_seach_blockx_410_goal), .data_out(_seach_blockx_410_data_out), .map_block(_seach_blockx_410_map_block), .now(_seach_blockx_410_now));
seach_block seach_blockx_409 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_409_in_do), .start(_seach_blockx_409_start), .goal(_seach_blockx_409_goal), .data_out(_seach_blockx_409_data_out), .map_block(_seach_blockx_409_map_block), .now(_seach_blockx_409_now));
seach_block seach_blockx_408 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_408_in_do), .start(_seach_blockx_408_start), .goal(_seach_blockx_408_goal), .data_out(_seach_blockx_408_data_out), .map_block(_seach_blockx_408_map_block), .now(_seach_blockx_408_now));
seach_block seach_blockx_407 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_407_in_do), .start(_seach_blockx_407_start), .goal(_seach_blockx_407_goal), .data_out(_seach_blockx_407_data_out), .map_block(_seach_blockx_407_map_block), .now(_seach_blockx_407_now));
seach_block seach_blockx_406 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_406_in_do), .start(_seach_blockx_406_start), .goal(_seach_blockx_406_goal), .data_out(_seach_blockx_406_data_out), .map_block(_seach_blockx_406_map_block), .now(_seach_blockx_406_now));
seach_block seach_blockx_405 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_405_in_do), .start(_seach_blockx_405_start), .goal(_seach_blockx_405_goal), .data_out(_seach_blockx_405_data_out), .map_block(_seach_blockx_405_map_block), .now(_seach_blockx_405_now));
seach_block seach_blockx_404 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_404_in_do), .start(_seach_blockx_404_start), .goal(_seach_blockx_404_goal), .data_out(_seach_blockx_404_data_out), .map_block(_seach_blockx_404_map_block), .now(_seach_blockx_404_now));
seach_block seach_blockx_403 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_403_in_do), .start(_seach_blockx_403_start), .goal(_seach_blockx_403_goal), .data_out(_seach_blockx_403_data_out), .map_block(_seach_blockx_403_map_block), .now(_seach_blockx_403_now));
seach_block seach_blockx_402 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_402_in_do), .start(_seach_blockx_402_start), .goal(_seach_blockx_402_goal), .data_out(_seach_blockx_402_data_out), .map_block(_seach_blockx_402_map_block), .now(_seach_blockx_402_now));
seach_block seach_blockx_401 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_401_in_do), .start(_seach_blockx_401_start), .goal(_seach_blockx_401_goal), .data_out(_seach_blockx_401_data_out), .map_block(_seach_blockx_401_map_block), .now(_seach_blockx_401_now));
seach_block seach_blockx_400 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_400_in_do), .start(_seach_blockx_400_start), .goal(_seach_blockx_400_goal), .data_out(_seach_blockx_400_data_out), .map_block(_seach_blockx_400_map_block), .now(_seach_blockx_400_now));
seach_block seach_blockx_399 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_399_in_do), .start(_seach_blockx_399_start), .goal(_seach_blockx_399_goal), .data_out(_seach_blockx_399_data_out), .map_block(_seach_blockx_399_map_block), .now(_seach_blockx_399_now));
seach_block seach_blockx_398 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_398_in_do), .start(_seach_blockx_398_start), .goal(_seach_blockx_398_goal), .data_out(_seach_blockx_398_data_out), .map_block(_seach_blockx_398_map_block), .now(_seach_blockx_398_now));
seach_block seach_blockx_397 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_397_in_do), .start(_seach_blockx_397_start), .goal(_seach_blockx_397_goal), .data_out(_seach_blockx_397_data_out), .map_block(_seach_blockx_397_map_block), .now(_seach_blockx_397_now));
seach_block seach_blockx_396 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_396_in_do), .start(_seach_blockx_396_start), .goal(_seach_blockx_396_goal), .data_out(_seach_blockx_396_data_out), .map_block(_seach_blockx_396_map_block), .now(_seach_blockx_396_now));
seach_block seach_blockx_395 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_395_in_do), .start(_seach_blockx_395_start), .goal(_seach_blockx_395_goal), .data_out(_seach_blockx_395_data_out), .map_block(_seach_blockx_395_map_block), .now(_seach_blockx_395_now));
seach_block seach_blockx_394 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_394_in_do), .start(_seach_blockx_394_start), .goal(_seach_blockx_394_goal), .data_out(_seach_blockx_394_data_out), .map_block(_seach_blockx_394_map_block), .now(_seach_blockx_394_now));
seach_block seach_blockx_393 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_393_in_do), .start(_seach_blockx_393_start), .goal(_seach_blockx_393_goal), .data_out(_seach_blockx_393_data_out), .map_block(_seach_blockx_393_map_block), .now(_seach_blockx_393_now));
seach_block seach_blockx_392 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_392_in_do), .start(_seach_blockx_392_start), .goal(_seach_blockx_392_goal), .data_out(_seach_blockx_392_data_out), .map_block(_seach_blockx_392_map_block), .now(_seach_blockx_392_now));
seach_block seach_blockx_391 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_391_in_do), .start(_seach_blockx_391_start), .goal(_seach_blockx_391_goal), .data_out(_seach_blockx_391_data_out), .map_block(_seach_blockx_391_map_block), .now(_seach_blockx_391_now));
seach_block seach_blockx_390 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_390_in_do), .start(_seach_blockx_390_start), .goal(_seach_blockx_390_goal), .data_out(_seach_blockx_390_data_out), .map_block(_seach_blockx_390_map_block), .now(_seach_blockx_390_now));
seach_block seach_blockx_389 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_389_in_do), .start(_seach_blockx_389_start), .goal(_seach_blockx_389_goal), .data_out(_seach_blockx_389_data_out), .map_block(_seach_blockx_389_map_block), .now(_seach_blockx_389_now));
seach_block seach_blockx_388 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_388_in_do), .start(_seach_blockx_388_start), .goal(_seach_blockx_388_goal), .data_out(_seach_blockx_388_data_out), .map_block(_seach_blockx_388_map_block), .now(_seach_blockx_388_now));
seach_block seach_blockx_387 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_387_in_do), .start(_seach_blockx_387_start), .goal(_seach_blockx_387_goal), .data_out(_seach_blockx_387_data_out), .map_block(_seach_blockx_387_map_block), .now(_seach_blockx_387_now));
seach_block seach_blockx_386 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_386_in_do), .start(_seach_blockx_386_start), .goal(_seach_blockx_386_goal), .data_out(_seach_blockx_386_data_out), .map_block(_seach_blockx_386_map_block), .now(_seach_blockx_386_now));
seach_block seach_blockx_385 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_385_in_do), .start(_seach_blockx_385_start), .goal(_seach_blockx_385_goal), .data_out(_seach_blockx_385_data_out), .map_block(_seach_blockx_385_map_block), .now(_seach_blockx_385_now));
seach_block seach_blockx_384 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_384_in_do), .start(_seach_blockx_384_start), .goal(_seach_blockx_384_goal), .data_out(_seach_blockx_384_data_out), .map_block(_seach_blockx_384_map_block), .now(_seach_blockx_384_now));
seach_block seach_blockx_383 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_383_in_do), .start(_seach_blockx_383_start), .goal(_seach_blockx_383_goal), .data_out(_seach_blockx_383_data_out), .map_block(_seach_blockx_383_map_block), .now(_seach_blockx_383_now));
seach_block seach_blockx_382 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_382_in_do), .start(_seach_blockx_382_start), .goal(_seach_blockx_382_goal), .data_out(_seach_blockx_382_data_out), .map_block(_seach_blockx_382_map_block), .now(_seach_blockx_382_now));
seach_block seach_blockx_381 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_381_in_do), .start(_seach_blockx_381_start), .goal(_seach_blockx_381_goal), .data_out(_seach_blockx_381_data_out), .map_block(_seach_blockx_381_map_block), .now(_seach_blockx_381_now));
seach_block seach_blockx_380 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_380_in_do), .start(_seach_blockx_380_start), .goal(_seach_blockx_380_goal), .data_out(_seach_blockx_380_data_out), .map_block(_seach_blockx_380_map_block), .now(_seach_blockx_380_now));
seach_block seach_blockx_379 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_379_in_do), .start(_seach_blockx_379_start), .goal(_seach_blockx_379_goal), .data_out(_seach_blockx_379_data_out), .map_block(_seach_blockx_379_map_block), .now(_seach_blockx_379_now));
seach_block seach_blockx_378 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_378_in_do), .start(_seach_blockx_378_start), .goal(_seach_blockx_378_goal), .data_out(_seach_blockx_378_data_out), .map_block(_seach_blockx_378_map_block), .now(_seach_blockx_378_now));
seach_block seach_blockx_377 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_377_in_do), .start(_seach_blockx_377_start), .goal(_seach_blockx_377_goal), .data_out(_seach_blockx_377_data_out), .map_block(_seach_blockx_377_map_block), .now(_seach_blockx_377_now));
seach_block seach_blockx_376 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_376_in_do), .start(_seach_blockx_376_start), .goal(_seach_blockx_376_goal), .data_out(_seach_blockx_376_data_out), .map_block(_seach_blockx_376_map_block), .now(_seach_blockx_376_now));
seach_block seach_blockx_375 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_375_in_do), .start(_seach_blockx_375_start), .goal(_seach_blockx_375_goal), .data_out(_seach_blockx_375_data_out), .map_block(_seach_blockx_375_map_block), .now(_seach_blockx_375_now));
seach_block seach_blockx_374 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_374_in_do), .start(_seach_blockx_374_start), .goal(_seach_blockx_374_goal), .data_out(_seach_blockx_374_data_out), .map_block(_seach_blockx_374_map_block), .now(_seach_blockx_374_now));
seach_block seach_blockx_373 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_373_in_do), .start(_seach_blockx_373_start), .goal(_seach_blockx_373_goal), .data_out(_seach_blockx_373_data_out), .map_block(_seach_blockx_373_map_block), .now(_seach_blockx_373_now));
seach_block seach_blockx_372 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_372_in_do), .start(_seach_blockx_372_start), .goal(_seach_blockx_372_goal), .data_out(_seach_blockx_372_data_out), .map_block(_seach_blockx_372_map_block), .now(_seach_blockx_372_now));
seach_block seach_blockx_371 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_371_in_do), .start(_seach_blockx_371_start), .goal(_seach_blockx_371_goal), .data_out(_seach_blockx_371_data_out), .map_block(_seach_blockx_371_map_block), .now(_seach_blockx_371_now));
seach_block seach_blockx_370 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_370_in_do), .start(_seach_blockx_370_start), .goal(_seach_blockx_370_goal), .data_out(_seach_blockx_370_data_out), .map_block(_seach_blockx_370_map_block), .now(_seach_blockx_370_now));
seach_block seach_blockx_369 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_369_in_do), .start(_seach_blockx_369_start), .goal(_seach_blockx_369_goal), .data_out(_seach_blockx_369_data_out), .map_block(_seach_blockx_369_map_block), .now(_seach_blockx_369_now));
seach_block seach_blockx_368 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_368_in_do), .start(_seach_blockx_368_start), .goal(_seach_blockx_368_goal), .data_out(_seach_blockx_368_data_out), .map_block(_seach_blockx_368_map_block), .now(_seach_blockx_368_now));
seach_block seach_blockx_367 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_367_in_do), .start(_seach_blockx_367_start), .goal(_seach_blockx_367_goal), .data_out(_seach_blockx_367_data_out), .map_block(_seach_blockx_367_map_block), .now(_seach_blockx_367_now));
seach_block seach_blockx_366 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_366_in_do), .start(_seach_blockx_366_start), .goal(_seach_blockx_366_goal), .data_out(_seach_blockx_366_data_out), .map_block(_seach_blockx_366_map_block), .now(_seach_blockx_366_now));
seach_block seach_blockx_365 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_365_in_do), .start(_seach_blockx_365_start), .goal(_seach_blockx_365_goal), .data_out(_seach_blockx_365_data_out), .map_block(_seach_blockx_365_map_block), .now(_seach_blockx_365_now));
seach_block seach_blockx_364 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_364_in_do), .start(_seach_blockx_364_start), .goal(_seach_blockx_364_goal), .data_out(_seach_blockx_364_data_out), .map_block(_seach_blockx_364_map_block), .now(_seach_blockx_364_now));
seach_block seach_blockx_363 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_363_in_do), .start(_seach_blockx_363_start), .goal(_seach_blockx_363_goal), .data_out(_seach_blockx_363_data_out), .map_block(_seach_blockx_363_map_block), .now(_seach_blockx_363_now));
seach_block seach_blockx_362 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_362_in_do), .start(_seach_blockx_362_start), .goal(_seach_blockx_362_goal), .data_out(_seach_blockx_362_data_out), .map_block(_seach_blockx_362_map_block), .now(_seach_blockx_362_now));
seach_block seach_blockx_361 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_361_in_do), .start(_seach_blockx_361_start), .goal(_seach_blockx_361_goal), .data_out(_seach_blockx_361_data_out), .map_block(_seach_blockx_361_map_block), .now(_seach_blockx_361_now));
seach_block seach_blockx_360 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_360_in_do), .start(_seach_blockx_360_start), .goal(_seach_blockx_360_goal), .data_out(_seach_blockx_360_data_out), .map_block(_seach_blockx_360_map_block), .now(_seach_blockx_360_now));
seach_block seach_blockx_359 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_359_in_do), .start(_seach_blockx_359_start), .goal(_seach_blockx_359_goal), .data_out(_seach_blockx_359_data_out), .map_block(_seach_blockx_359_map_block), .now(_seach_blockx_359_now));
seach_block seach_blockx_358 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_358_in_do), .start(_seach_blockx_358_start), .goal(_seach_blockx_358_goal), .data_out(_seach_blockx_358_data_out), .map_block(_seach_blockx_358_map_block), .now(_seach_blockx_358_now));
seach_block seach_blockx_357 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_357_in_do), .start(_seach_blockx_357_start), .goal(_seach_blockx_357_goal), .data_out(_seach_blockx_357_data_out), .map_block(_seach_blockx_357_map_block), .now(_seach_blockx_357_now));
seach_block seach_blockx_356 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_356_in_do), .start(_seach_blockx_356_start), .goal(_seach_blockx_356_goal), .data_out(_seach_blockx_356_data_out), .map_block(_seach_blockx_356_map_block), .now(_seach_blockx_356_now));
seach_block seach_blockx_355 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_355_in_do), .start(_seach_blockx_355_start), .goal(_seach_blockx_355_goal), .data_out(_seach_blockx_355_data_out), .map_block(_seach_blockx_355_map_block), .now(_seach_blockx_355_now));
seach_block seach_blockx_354 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_354_in_do), .start(_seach_blockx_354_start), .goal(_seach_blockx_354_goal), .data_out(_seach_blockx_354_data_out), .map_block(_seach_blockx_354_map_block), .now(_seach_blockx_354_now));
seach_block seach_blockx_353 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_353_in_do), .start(_seach_blockx_353_start), .goal(_seach_blockx_353_goal), .data_out(_seach_blockx_353_data_out), .map_block(_seach_blockx_353_map_block), .now(_seach_blockx_353_now));
seach_block seach_blockx_352 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_352_in_do), .start(_seach_blockx_352_start), .goal(_seach_blockx_352_goal), .data_out(_seach_blockx_352_data_out), .map_block(_seach_blockx_352_map_block), .now(_seach_blockx_352_now));
seach_block seach_blockx_351 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_351_in_do), .start(_seach_blockx_351_start), .goal(_seach_blockx_351_goal), .data_out(_seach_blockx_351_data_out), .map_block(_seach_blockx_351_map_block), .now(_seach_blockx_351_now));
seach_block seach_blockx_350 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_350_in_do), .start(_seach_blockx_350_start), .goal(_seach_blockx_350_goal), .data_out(_seach_blockx_350_data_out), .map_block(_seach_blockx_350_map_block), .now(_seach_blockx_350_now));
seach_block seach_blockx_349 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_349_in_do), .start(_seach_blockx_349_start), .goal(_seach_blockx_349_goal), .data_out(_seach_blockx_349_data_out), .map_block(_seach_blockx_349_map_block), .now(_seach_blockx_349_now));
seach_block seach_blockx_348 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_348_in_do), .start(_seach_blockx_348_start), .goal(_seach_blockx_348_goal), .data_out(_seach_blockx_348_data_out), .map_block(_seach_blockx_348_map_block), .now(_seach_blockx_348_now));
seach_block seach_blockx_347 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_347_in_do), .start(_seach_blockx_347_start), .goal(_seach_blockx_347_goal), .data_out(_seach_blockx_347_data_out), .map_block(_seach_blockx_347_map_block), .now(_seach_blockx_347_now));
seach_block seach_blockx_346 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_346_in_do), .start(_seach_blockx_346_start), .goal(_seach_blockx_346_goal), .data_out(_seach_blockx_346_data_out), .map_block(_seach_blockx_346_map_block), .now(_seach_blockx_346_now));
seach_block seach_blockx_345 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_345_in_do), .start(_seach_blockx_345_start), .goal(_seach_blockx_345_goal), .data_out(_seach_blockx_345_data_out), .map_block(_seach_blockx_345_map_block), .now(_seach_blockx_345_now));
seach_block seach_blockx_344 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_344_in_do), .start(_seach_blockx_344_start), .goal(_seach_blockx_344_goal), .data_out(_seach_blockx_344_data_out), .map_block(_seach_blockx_344_map_block), .now(_seach_blockx_344_now));
seach_block seach_blockx_343 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_343_in_do), .start(_seach_blockx_343_start), .goal(_seach_blockx_343_goal), .data_out(_seach_blockx_343_data_out), .map_block(_seach_blockx_343_map_block), .now(_seach_blockx_343_now));
seach_block seach_blockx_342 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_342_in_do), .start(_seach_blockx_342_start), .goal(_seach_blockx_342_goal), .data_out(_seach_blockx_342_data_out), .map_block(_seach_blockx_342_map_block), .now(_seach_blockx_342_now));
seach_block seach_blockx_341 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_341_in_do), .start(_seach_blockx_341_start), .goal(_seach_blockx_341_goal), .data_out(_seach_blockx_341_data_out), .map_block(_seach_blockx_341_map_block), .now(_seach_blockx_341_now));
seach_block seach_blockx_340 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_340_in_do), .start(_seach_blockx_340_start), .goal(_seach_blockx_340_goal), .data_out(_seach_blockx_340_data_out), .map_block(_seach_blockx_340_map_block), .now(_seach_blockx_340_now));
seach_block seach_blockx_339 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_339_in_do), .start(_seach_blockx_339_start), .goal(_seach_blockx_339_goal), .data_out(_seach_blockx_339_data_out), .map_block(_seach_blockx_339_map_block), .now(_seach_blockx_339_now));
seach_block seach_blockx_338 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_338_in_do), .start(_seach_blockx_338_start), .goal(_seach_blockx_338_goal), .data_out(_seach_blockx_338_data_out), .map_block(_seach_blockx_338_map_block), .now(_seach_blockx_338_now));
seach_block seach_blockx_337 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_337_in_do), .start(_seach_blockx_337_start), .goal(_seach_blockx_337_goal), .data_out(_seach_blockx_337_data_out), .map_block(_seach_blockx_337_map_block), .now(_seach_blockx_337_now));
seach_block seach_blockx_336 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_336_in_do), .start(_seach_blockx_336_start), .goal(_seach_blockx_336_goal), .data_out(_seach_blockx_336_data_out), .map_block(_seach_blockx_336_map_block), .now(_seach_blockx_336_now));
seach_block seach_blockx_335 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_335_in_do), .start(_seach_blockx_335_start), .goal(_seach_blockx_335_goal), .data_out(_seach_blockx_335_data_out), .map_block(_seach_blockx_335_map_block), .now(_seach_blockx_335_now));
seach_block seach_blockx_334 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_334_in_do), .start(_seach_blockx_334_start), .goal(_seach_blockx_334_goal), .data_out(_seach_blockx_334_data_out), .map_block(_seach_blockx_334_map_block), .now(_seach_blockx_334_now));
seach_block seach_blockx_333 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_333_in_do), .start(_seach_blockx_333_start), .goal(_seach_blockx_333_goal), .data_out(_seach_blockx_333_data_out), .map_block(_seach_blockx_333_map_block), .now(_seach_blockx_333_now));
seach_block seach_blockx_332 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_332_in_do), .start(_seach_blockx_332_start), .goal(_seach_blockx_332_goal), .data_out(_seach_blockx_332_data_out), .map_block(_seach_blockx_332_map_block), .now(_seach_blockx_332_now));
seach_block seach_blockx_331 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_331_in_do), .start(_seach_blockx_331_start), .goal(_seach_blockx_331_goal), .data_out(_seach_blockx_331_data_out), .map_block(_seach_blockx_331_map_block), .now(_seach_blockx_331_now));
seach_block seach_blockx_330 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_330_in_do), .start(_seach_blockx_330_start), .goal(_seach_blockx_330_goal), .data_out(_seach_blockx_330_data_out), .map_block(_seach_blockx_330_map_block), .now(_seach_blockx_330_now));
seach_block seach_blockx_329 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_329_in_do), .start(_seach_blockx_329_start), .goal(_seach_blockx_329_goal), .data_out(_seach_blockx_329_data_out), .map_block(_seach_blockx_329_map_block), .now(_seach_blockx_329_now));
seach_block seach_blockx_328 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_328_in_do), .start(_seach_blockx_328_start), .goal(_seach_blockx_328_goal), .data_out(_seach_blockx_328_data_out), .map_block(_seach_blockx_328_map_block), .now(_seach_blockx_328_now));
seach_block seach_blockx_327 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_327_in_do), .start(_seach_blockx_327_start), .goal(_seach_blockx_327_goal), .data_out(_seach_blockx_327_data_out), .map_block(_seach_blockx_327_map_block), .now(_seach_blockx_327_now));
seach_block seach_blockx_326 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_326_in_do), .start(_seach_blockx_326_start), .goal(_seach_blockx_326_goal), .data_out(_seach_blockx_326_data_out), .map_block(_seach_blockx_326_map_block), .now(_seach_blockx_326_now));
seach_block seach_blockx_325 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_325_in_do), .start(_seach_blockx_325_start), .goal(_seach_blockx_325_goal), .data_out(_seach_blockx_325_data_out), .map_block(_seach_blockx_325_map_block), .now(_seach_blockx_325_now));
seach_block seach_blockx_324 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_324_in_do), .start(_seach_blockx_324_start), .goal(_seach_blockx_324_goal), .data_out(_seach_blockx_324_data_out), .map_block(_seach_blockx_324_map_block), .now(_seach_blockx_324_now));
seach_block seach_blockx_323 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_323_in_do), .start(_seach_blockx_323_start), .goal(_seach_blockx_323_goal), .data_out(_seach_blockx_323_data_out), .map_block(_seach_blockx_323_map_block), .now(_seach_blockx_323_now));
seach_block seach_blockx_322 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_322_in_do), .start(_seach_blockx_322_start), .goal(_seach_blockx_322_goal), .data_out(_seach_blockx_322_data_out), .map_block(_seach_blockx_322_map_block), .now(_seach_blockx_322_now));
seach_block seach_blockx_321 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_321_in_do), .start(_seach_blockx_321_start), .goal(_seach_blockx_321_goal), .data_out(_seach_blockx_321_data_out), .map_block(_seach_blockx_321_map_block), .now(_seach_blockx_321_now));
seach_block seach_blockx_320 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_320_in_do), .start(_seach_blockx_320_start), .goal(_seach_blockx_320_goal), .data_out(_seach_blockx_320_data_out), .map_block(_seach_blockx_320_map_block), .now(_seach_blockx_320_now));
seach_block seach_blockx_319 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_319_in_do), .start(_seach_blockx_319_start), .goal(_seach_blockx_319_goal), .data_out(_seach_blockx_319_data_out), .map_block(_seach_blockx_319_map_block), .now(_seach_blockx_319_now));
seach_block seach_blockx_318 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_318_in_do), .start(_seach_blockx_318_start), .goal(_seach_blockx_318_goal), .data_out(_seach_blockx_318_data_out), .map_block(_seach_blockx_318_map_block), .now(_seach_blockx_318_now));
seach_block seach_blockx_317 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_317_in_do), .start(_seach_blockx_317_start), .goal(_seach_blockx_317_goal), .data_out(_seach_blockx_317_data_out), .map_block(_seach_blockx_317_map_block), .now(_seach_blockx_317_now));
seach_block seach_blockx_316 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_316_in_do), .start(_seach_blockx_316_start), .goal(_seach_blockx_316_goal), .data_out(_seach_blockx_316_data_out), .map_block(_seach_blockx_316_map_block), .now(_seach_blockx_316_now));
seach_block seach_blockx_315 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_315_in_do), .start(_seach_blockx_315_start), .goal(_seach_blockx_315_goal), .data_out(_seach_blockx_315_data_out), .map_block(_seach_blockx_315_map_block), .now(_seach_blockx_315_now));
seach_block seach_blockx_314 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_314_in_do), .start(_seach_blockx_314_start), .goal(_seach_blockx_314_goal), .data_out(_seach_blockx_314_data_out), .map_block(_seach_blockx_314_map_block), .now(_seach_blockx_314_now));
seach_block seach_blockx_313 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_313_in_do), .start(_seach_blockx_313_start), .goal(_seach_blockx_313_goal), .data_out(_seach_blockx_313_data_out), .map_block(_seach_blockx_313_map_block), .now(_seach_blockx_313_now));
seach_block seach_blockx_312 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_312_in_do), .start(_seach_blockx_312_start), .goal(_seach_blockx_312_goal), .data_out(_seach_blockx_312_data_out), .map_block(_seach_blockx_312_map_block), .now(_seach_blockx_312_now));
seach_block seach_blockx_311 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_311_in_do), .start(_seach_blockx_311_start), .goal(_seach_blockx_311_goal), .data_out(_seach_blockx_311_data_out), .map_block(_seach_blockx_311_map_block), .now(_seach_blockx_311_now));
seach_block seach_blockx_310 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_310_in_do), .start(_seach_blockx_310_start), .goal(_seach_blockx_310_goal), .data_out(_seach_blockx_310_data_out), .map_block(_seach_blockx_310_map_block), .now(_seach_blockx_310_now));
seach_block seach_blockx_309 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_309_in_do), .start(_seach_blockx_309_start), .goal(_seach_blockx_309_goal), .data_out(_seach_blockx_309_data_out), .map_block(_seach_blockx_309_map_block), .now(_seach_blockx_309_now));
seach_block seach_blockx_308 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_308_in_do), .start(_seach_blockx_308_start), .goal(_seach_blockx_308_goal), .data_out(_seach_blockx_308_data_out), .map_block(_seach_blockx_308_map_block), .now(_seach_blockx_308_now));
seach_block seach_blockx_307 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_307_in_do), .start(_seach_blockx_307_start), .goal(_seach_blockx_307_goal), .data_out(_seach_blockx_307_data_out), .map_block(_seach_blockx_307_map_block), .now(_seach_blockx_307_now));
seach_block seach_blockx_306 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_306_in_do), .start(_seach_blockx_306_start), .goal(_seach_blockx_306_goal), .data_out(_seach_blockx_306_data_out), .map_block(_seach_blockx_306_map_block), .now(_seach_blockx_306_now));
seach_block seach_blockx_305 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_305_in_do), .start(_seach_blockx_305_start), .goal(_seach_blockx_305_goal), .data_out(_seach_blockx_305_data_out), .map_block(_seach_blockx_305_map_block), .now(_seach_blockx_305_now));
seach_block seach_blockx_304 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_304_in_do), .start(_seach_blockx_304_start), .goal(_seach_blockx_304_goal), .data_out(_seach_blockx_304_data_out), .map_block(_seach_blockx_304_map_block), .now(_seach_blockx_304_now));
seach_block seach_blockx_303 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_303_in_do), .start(_seach_blockx_303_start), .goal(_seach_blockx_303_goal), .data_out(_seach_blockx_303_data_out), .map_block(_seach_blockx_303_map_block), .now(_seach_blockx_303_now));
seach_block seach_blockx_302 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_302_in_do), .start(_seach_blockx_302_start), .goal(_seach_blockx_302_goal), .data_out(_seach_blockx_302_data_out), .map_block(_seach_blockx_302_map_block), .now(_seach_blockx_302_now));
seach_block seach_blockx_301 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_301_in_do), .start(_seach_blockx_301_start), .goal(_seach_blockx_301_goal), .data_out(_seach_blockx_301_data_out), .map_block(_seach_blockx_301_map_block), .now(_seach_blockx_301_now));
seach_block seach_blockx_300 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_300_in_do), .start(_seach_blockx_300_start), .goal(_seach_blockx_300_goal), .data_out(_seach_blockx_300_data_out), .map_block(_seach_blockx_300_map_block), .now(_seach_blockx_300_now));
seach_block seach_blockx_299 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_299_in_do), .start(_seach_blockx_299_start), .goal(_seach_blockx_299_goal), .data_out(_seach_blockx_299_data_out), .map_block(_seach_blockx_299_map_block), .now(_seach_blockx_299_now));
seach_block seach_blockx_298 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_298_in_do), .start(_seach_blockx_298_start), .goal(_seach_blockx_298_goal), .data_out(_seach_blockx_298_data_out), .map_block(_seach_blockx_298_map_block), .now(_seach_blockx_298_now));
seach_block seach_blockx_297 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_297_in_do), .start(_seach_blockx_297_start), .goal(_seach_blockx_297_goal), .data_out(_seach_blockx_297_data_out), .map_block(_seach_blockx_297_map_block), .now(_seach_blockx_297_now));
seach_block seach_blockx_296 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_296_in_do), .start(_seach_blockx_296_start), .goal(_seach_blockx_296_goal), .data_out(_seach_blockx_296_data_out), .map_block(_seach_blockx_296_map_block), .now(_seach_blockx_296_now));
seach_block seach_blockx_295 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_295_in_do), .start(_seach_blockx_295_start), .goal(_seach_blockx_295_goal), .data_out(_seach_blockx_295_data_out), .map_block(_seach_blockx_295_map_block), .now(_seach_blockx_295_now));
seach_block seach_blockx_294 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_294_in_do), .start(_seach_blockx_294_start), .goal(_seach_blockx_294_goal), .data_out(_seach_blockx_294_data_out), .map_block(_seach_blockx_294_map_block), .now(_seach_blockx_294_now));
seach_block seach_blockx_293 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_293_in_do), .start(_seach_blockx_293_start), .goal(_seach_blockx_293_goal), .data_out(_seach_blockx_293_data_out), .map_block(_seach_blockx_293_map_block), .now(_seach_blockx_293_now));
seach_block seach_blockx_292 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_292_in_do), .start(_seach_blockx_292_start), .goal(_seach_blockx_292_goal), .data_out(_seach_blockx_292_data_out), .map_block(_seach_blockx_292_map_block), .now(_seach_blockx_292_now));
seach_block seach_blockx_291 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_291_in_do), .start(_seach_blockx_291_start), .goal(_seach_blockx_291_goal), .data_out(_seach_blockx_291_data_out), .map_block(_seach_blockx_291_map_block), .now(_seach_blockx_291_now));
seach_block seach_blockx_290 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_290_in_do), .start(_seach_blockx_290_start), .goal(_seach_blockx_290_goal), .data_out(_seach_blockx_290_data_out), .map_block(_seach_blockx_290_map_block), .now(_seach_blockx_290_now));
seach_block seach_blockx_289 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_289_in_do), .start(_seach_blockx_289_start), .goal(_seach_blockx_289_goal), .data_out(_seach_blockx_289_data_out), .map_block(_seach_blockx_289_map_block), .now(_seach_blockx_289_now));
seach_block seach_blockx_288 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_288_in_do), .start(_seach_blockx_288_start), .goal(_seach_blockx_288_goal), .data_out(_seach_blockx_288_data_out), .map_block(_seach_blockx_288_map_block), .now(_seach_blockx_288_now));
seach_block seach_blockx_287 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_287_in_do), .start(_seach_blockx_287_start), .goal(_seach_blockx_287_goal), .data_out(_seach_blockx_287_data_out), .map_block(_seach_blockx_287_map_block), .now(_seach_blockx_287_now));
seach_block seach_blockx_286 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_286_in_do), .start(_seach_blockx_286_start), .goal(_seach_blockx_286_goal), .data_out(_seach_blockx_286_data_out), .map_block(_seach_blockx_286_map_block), .now(_seach_blockx_286_now));
seach_block seach_blockx_285 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_285_in_do), .start(_seach_blockx_285_start), .goal(_seach_blockx_285_goal), .data_out(_seach_blockx_285_data_out), .map_block(_seach_blockx_285_map_block), .now(_seach_blockx_285_now));
seach_block seach_blockx_284 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_284_in_do), .start(_seach_blockx_284_start), .goal(_seach_blockx_284_goal), .data_out(_seach_blockx_284_data_out), .map_block(_seach_blockx_284_map_block), .now(_seach_blockx_284_now));
seach_block seach_blockx_283 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_283_in_do), .start(_seach_blockx_283_start), .goal(_seach_blockx_283_goal), .data_out(_seach_blockx_283_data_out), .map_block(_seach_blockx_283_map_block), .now(_seach_blockx_283_now));
seach_block seach_blockx_282 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_282_in_do), .start(_seach_blockx_282_start), .goal(_seach_blockx_282_goal), .data_out(_seach_blockx_282_data_out), .map_block(_seach_blockx_282_map_block), .now(_seach_blockx_282_now));
seach_block seach_blockx_281 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_281_in_do), .start(_seach_blockx_281_start), .goal(_seach_blockx_281_goal), .data_out(_seach_blockx_281_data_out), .map_block(_seach_blockx_281_map_block), .now(_seach_blockx_281_now));
seach_block seach_blockx_280 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_280_in_do), .start(_seach_blockx_280_start), .goal(_seach_blockx_280_goal), .data_out(_seach_blockx_280_data_out), .map_block(_seach_blockx_280_map_block), .now(_seach_blockx_280_now));
seach_block seach_blockx_279 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_279_in_do), .start(_seach_blockx_279_start), .goal(_seach_blockx_279_goal), .data_out(_seach_blockx_279_data_out), .map_block(_seach_blockx_279_map_block), .now(_seach_blockx_279_now));
seach_block seach_blockx_278 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_278_in_do), .start(_seach_blockx_278_start), .goal(_seach_blockx_278_goal), .data_out(_seach_blockx_278_data_out), .map_block(_seach_blockx_278_map_block), .now(_seach_blockx_278_now));
seach_block seach_blockx_277 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_277_in_do), .start(_seach_blockx_277_start), .goal(_seach_blockx_277_goal), .data_out(_seach_blockx_277_data_out), .map_block(_seach_blockx_277_map_block), .now(_seach_blockx_277_now));
seach_block seach_blockx_276 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_276_in_do), .start(_seach_blockx_276_start), .goal(_seach_blockx_276_goal), .data_out(_seach_blockx_276_data_out), .map_block(_seach_blockx_276_map_block), .now(_seach_blockx_276_now));
seach_block seach_blockx_275 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_275_in_do), .start(_seach_blockx_275_start), .goal(_seach_blockx_275_goal), .data_out(_seach_blockx_275_data_out), .map_block(_seach_blockx_275_map_block), .now(_seach_blockx_275_now));
seach_block seach_blockx_274 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_274_in_do), .start(_seach_blockx_274_start), .goal(_seach_blockx_274_goal), .data_out(_seach_blockx_274_data_out), .map_block(_seach_blockx_274_map_block), .now(_seach_blockx_274_now));
seach_block seach_blockx_273 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_273_in_do), .start(_seach_blockx_273_start), .goal(_seach_blockx_273_goal), .data_out(_seach_blockx_273_data_out), .map_block(_seach_blockx_273_map_block), .now(_seach_blockx_273_now));
seach_block seach_blockx_272 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_272_in_do), .start(_seach_blockx_272_start), .goal(_seach_blockx_272_goal), .data_out(_seach_blockx_272_data_out), .map_block(_seach_blockx_272_map_block), .now(_seach_blockx_272_now));
seach_block seach_blockx_271 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_271_in_do), .start(_seach_blockx_271_start), .goal(_seach_blockx_271_goal), .data_out(_seach_blockx_271_data_out), .map_block(_seach_blockx_271_map_block), .now(_seach_blockx_271_now));
seach_block seach_blockx_270 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_270_in_do), .start(_seach_blockx_270_start), .goal(_seach_blockx_270_goal), .data_out(_seach_blockx_270_data_out), .map_block(_seach_blockx_270_map_block), .now(_seach_blockx_270_now));
seach_block seach_blockx_269 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_269_in_do), .start(_seach_blockx_269_start), .goal(_seach_blockx_269_goal), .data_out(_seach_blockx_269_data_out), .map_block(_seach_blockx_269_map_block), .now(_seach_blockx_269_now));
seach_block seach_blockx_268 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_268_in_do), .start(_seach_blockx_268_start), .goal(_seach_blockx_268_goal), .data_out(_seach_blockx_268_data_out), .map_block(_seach_blockx_268_map_block), .now(_seach_blockx_268_now));
seach_block seach_blockx_267 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_267_in_do), .start(_seach_blockx_267_start), .goal(_seach_blockx_267_goal), .data_out(_seach_blockx_267_data_out), .map_block(_seach_blockx_267_map_block), .now(_seach_blockx_267_now));
seach_block seach_blockx_266 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_266_in_do), .start(_seach_blockx_266_start), .goal(_seach_blockx_266_goal), .data_out(_seach_blockx_266_data_out), .map_block(_seach_blockx_266_map_block), .now(_seach_blockx_266_now));
seach_block seach_blockx_265 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_265_in_do), .start(_seach_blockx_265_start), .goal(_seach_blockx_265_goal), .data_out(_seach_blockx_265_data_out), .map_block(_seach_blockx_265_map_block), .now(_seach_blockx_265_now));
seach_block seach_blockx_264 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_264_in_do), .start(_seach_blockx_264_start), .goal(_seach_blockx_264_goal), .data_out(_seach_blockx_264_data_out), .map_block(_seach_blockx_264_map_block), .now(_seach_blockx_264_now));
seach_block seach_blockx_263 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_263_in_do), .start(_seach_blockx_263_start), .goal(_seach_blockx_263_goal), .data_out(_seach_blockx_263_data_out), .map_block(_seach_blockx_263_map_block), .now(_seach_blockx_263_now));
seach_block seach_blockx_262 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_262_in_do), .start(_seach_blockx_262_start), .goal(_seach_blockx_262_goal), .data_out(_seach_blockx_262_data_out), .map_block(_seach_blockx_262_map_block), .now(_seach_blockx_262_now));
seach_block seach_blockx_261 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_261_in_do), .start(_seach_blockx_261_start), .goal(_seach_blockx_261_goal), .data_out(_seach_blockx_261_data_out), .map_block(_seach_blockx_261_map_block), .now(_seach_blockx_261_now));
seach_block seach_blockx_260 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_260_in_do), .start(_seach_blockx_260_start), .goal(_seach_blockx_260_goal), .data_out(_seach_blockx_260_data_out), .map_block(_seach_blockx_260_map_block), .now(_seach_blockx_260_now));
seach_block seach_blockx_259 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_259_in_do), .start(_seach_blockx_259_start), .goal(_seach_blockx_259_goal), .data_out(_seach_blockx_259_data_out), .map_block(_seach_blockx_259_map_block), .now(_seach_blockx_259_now));
seach_block seach_blockx_258 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_258_in_do), .start(_seach_blockx_258_start), .goal(_seach_blockx_258_goal), .data_out(_seach_blockx_258_data_out), .map_block(_seach_blockx_258_map_block), .now(_seach_blockx_258_now));
seach_block seach_blockx_257 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_257_in_do), .start(_seach_blockx_257_start), .goal(_seach_blockx_257_goal), .data_out(_seach_blockx_257_data_out), .map_block(_seach_blockx_257_map_block), .now(_seach_blockx_257_now));
seach_block seach_blockx_256 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_256_in_do), .start(_seach_blockx_256_start), .goal(_seach_blockx_256_goal), .data_out(_seach_blockx_256_data_out), .map_block(_seach_blockx_256_map_block), .now(_seach_blockx_256_now));
seach_block seach_blockx_255 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_255_in_do), .start(_seach_blockx_255_start), .goal(_seach_blockx_255_goal), .data_out(_seach_blockx_255_data_out), .map_block(_seach_blockx_255_map_block), .now(_seach_blockx_255_now));
seach_block seach_blockx_254 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_254_in_do), .start(_seach_blockx_254_start), .goal(_seach_blockx_254_goal), .data_out(_seach_blockx_254_data_out), .map_block(_seach_blockx_254_map_block), .now(_seach_blockx_254_now));
seach_block seach_blockx_253 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_253_in_do), .start(_seach_blockx_253_start), .goal(_seach_blockx_253_goal), .data_out(_seach_blockx_253_data_out), .map_block(_seach_blockx_253_map_block), .now(_seach_blockx_253_now));
seach_block seach_blockx_252 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_252_in_do), .start(_seach_blockx_252_start), .goal(_seach_blockx_252_goal), .data_out(_seach_blockx_252_data_out), .map_block(_seach_blockx_252_map_block), .now(_seach_blockx_252_now));
seach_block seach_blockx_251 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_251_in_do), .start(_seach_blockx_251_start), .goal(_seach_blockx_251_goal), .data_out(_seach_blockx_251_data_out), .map_block(_seach_blockx_251_map_block), .now(_seach_blockx_251_now));
seach_block seach_blockx_250 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_250_in_do), .start(_seach_blockx_250_start), .goal(_seach_blockx_250_goal), .data_out(_seach_blockx_250_data_out), .map_block(_seach_blockx_250_map_block), .now(_seach_blockx_250_now));
seach_block seach_blockx_249 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_249_in_do), .start(_seach_blockx_249_start), .goal(_seach_blockx_249_goal), .data_out(_seach_blockx_249_data_out), .map_block(_seach_blockx_249_map_block), .now(_seach_blockx_249_now));
seach_block seach_blockx_248 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_248_in_do), .start(_seach_blockx_248_start), .goal(_seach_blockx_248_goal), .data_out(_seach_blockx_248_data_out), .map_block(_seach_blockx_248_map_block), .now(_seach_blockx_248_now));
seach_block seach_blockx_247 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_247_in_do), .start(_seach_blockx_247_start), .goal(_seach_blockx_247_goal), .data_out(_seach_blockx_247_data_out), .map_block(_seach_blockx_247_map_block), .now(_seach_blockx_247_now));
seach_block seach_blockx_246 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_246_in_do), .start(_seach_blockx_246_start), .goal(_seach_blockx_246_goal), .data_out(_seach_blockx_246_data_out), .map_block(_seach_blockx_246_map_block), .now(_seach_blockx_246_now));
seach_block seach_blockx_245 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_245_in_do), .start(_seach_blockx_245_start), .goal(_seach_blockx_245_goal), .data_out(_seach_blockx_245_data_out), .map_block(_seach_blockx_245_map_block), .now(_seach_blockx_245_now));
seach_block seach_blockx_244 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_244_in_do), .start(_seach_blockx_244_start), .goal(_seach_blockx_244_goal), .data_out(_seach_blockx_244_data_out), .map_block(_seach_blockx_244_map_block), .now(_seach_blockx_244_now));
seach_block seach_blockx_243 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_243_in_do), .start(_seach_blockx_243_start), .goal(_seach_blockx_243_goal), .data_out(_seach_blockx_243_data_out), .map_block(_seach_blockx_243_map_block), .now(_seach_blockx_243_now));
seach_block seach_blockx_242 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_242_in_do), .start(_seach_blockx_242_start), .goal(_seach_blockx_242_goal), .data_out(_seach_blockx_242_data_out), .map_block(_seach_blockx_242_map_block), .now(_seach_blockx_242_now));
seach_block seach_blockx_241 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_241_in_do), .start(_seach_blockx_241_start), .goal(_seach_blockx_241_goal), .data_out(_seach_blockx_241_data_out), .map_block(_seach_blockx_241_map_block), .now(_seach_blockx_241_now));
seach_block seach_blockx_240 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_240_in_do), .start(_seach_blockx_240_start), .goal(_seach_blockx_240_goal), .data_out(_seach_blockx_240_data_out), .map_block(_seach_blockx_240_map_block), .now(_seach_blockx_240_now));
seach_block seach_blockx_239 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_239_in_do), .start(_seach_blockx_239_start), .goal(_seach_blockx_239_goal), .data_out(_seach_blockx_239_data_out), .map_block(_seach_blockx_239_map_block), .now(_seach_blockx_239_now));
seach_block seach_blockx_238 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_238_in_do), .start(_seach_blockx_238_start), .goal(_seach_blockx_238_goal), .data_out(_seach_blockx_238_data_out), .map_block(_seach_blockx_238_map_block), .now(_seach_blockx_238_now));
seach_block seach_blockx_237 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_237_in_do), .start(_seach_blockx_237_start), .goal(_seach_blockx_237_goal), .data_out(_seach_blockx_237_data_out), .map_block(_seach_blockx_237_map_block), .now(_seach_blockx_237_now));
seach_block seach_blockx_236 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_236_in_do), .start(_seach_blockx_236_start), .goal(_seach_blockx_236_goal), .data_out(_seach_blockx_236_data_out), .map_block(_seach_blockx_236_map_block), .now(_seach_blockx_236_now));
seach_block seach_blockx_235 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_235_in_do), .start(_seach_blockx_235_start), .goal(_seach_blockx_235_goal), .data_out(_seach_blockx_235_data_out), .map_block(_seach_blockx_235_map_block), .now(_seach_blockx_235_now));
seach_block seach_blockx_234 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_234_in_do), .start(_seach_blockx_234_start), .goal(_seach_blockx_234_goal), .data_out(_seach_blockx_234_data_out), .map_block(_seach_blockx_234_map_block), .now(_seach_blockx_234_now));
seach_block seach_blockx_233 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_233_in_do), .start(_seach_blockx_233_start), .goal(_seach_blockx_233_goal), .data_out(_seach_blockx_233_data_out), .map_block(_seach_blockx_233_map_block), .now(_seach_blockx_233_now));
seach_block seach_blockx_232 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_232_in_do), .start(_seach_blockx_232_start), .goal(_seach_blockx_232_goal), .data_out(_seach_blockx_232_data_out), .map_block(_seach_blockx_232_map_block), .now(_seach_blockx_232_now));
seach_block seach_blockx_231 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_231_in_do), .start(_seach_blockx_231_start), .goal(_seach_blockx_231_goal), .data_out(_seach_blockx_231_data_out), .map_block(_seach_blockx_231_map_block), .now(_seach_blockx_231_now));
seach_block seach_blockx_230 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_230_in_do), .start(_seach_blockx_230_start), .goal(_seach_blockx_230_goal), .data_out(_seach_blockx_230_data_out), .map_block(_seach_blockx_230_map_block), .now(_seach_blockx_230_now));
seach_block seach_blockx_229 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_229_in_do), .start(_seach_blockx_229_start), .goal(_seach_blockx_229_goal), .data_out(_seach_blockx_229_data_out), .map_block(_seach_blockx_229_map_block), .now(_seach_blockx_229_now));
seach_block seach_blockx_228 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_228_in_do), .start(_seach_blockx_228_start), .goal(_seach_blockx_228_goal), .data_out(_seach_blockx_228_data_out), .map_block(_seach_blockx_228_map_block), .now(_seach_blockx_228_now));
seach_block seach_blockx_227 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_227_in_do), .start(_seach_blockx_227_start), .goal(_seach_blockx_227_goal), .data_out(_seach_blockx_227_data_out), .map_block(_seach_blockx_227_map_block), .now(_seach_blockx_227_now));
seach_block seach_blockx_226 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_226_in_do), .start(_seach_blockx_226_start), .goal(_seach_blockx_226_goal), .data_out(_seach_blockx_226_data_out), .map_block(_seach_blockx_226_map_block), .now(_seach_blockx_226_now));
seach_block seach_blockx_225 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_225_in_do), .start(_seach_blockx_225_start), .goal(_seach_blockx_225_goal), .data_out(_seach_blockx_225_data_out), .map_block(_seach_blockx_225_map_block), .now(_seach_blockx_225_now));
seach_block seach_blockx_224 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_224_in_do), .start(_seach_blockx_224_start), .goal(_seach_blockx_224_goal), .data_out(_seach_blockx_224_data_out), .map_block(_seach_blockx_224_map_block), .now(_seach_blockx_224_now));
seach_block seach_blockx_223 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_223_in_do), .start(_seach_blockx_223_start), .goal(_seach_blockx_223_goal), .data_out(_seach_blockx_223_data_out), .map_block(_seach_blockx_223_map_block), .now(_seach_blockx_223_now));
seach_block seach_blockx_222 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_222_in_do), .start(_seach_blockx_222_start), .goal(_seach_blockx_222_goal), .data_out(_seach_blockx_222_data_out), .map_block(_seach_blockx_222_map_block), .now(_seach_blockx_222_now));
seach_block seach_blockx_221 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_221_in_do), .start(_seach_blockx_221_start), .goal(_seach_blockx_221_goal), .data_out(_seach_blockx_221_data_out), .map_block(_seach_blockx_221_map_block), .now(_seach_blockx_221_now));
seach_block seach_blockx_220 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_220_in_do), .start(_seach_blockx_220_start), .goal(_seach_blockx_220_goal), .data_out(_seach_blockx_220_data_out), .map_block(_seach_blockx_220_map_block), .now(_seach_blockx_220_now));
seach_block seach_blockx_219 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_219_in_do), .start(_seach_blockx_219_start), .goal(_seach_blockx_219_goal), .data_out(_seach_blockx_219_data_out), .map_block(_seach_blockx_219_map_block), .now(_seach_blockx_219_now));
seach_block seach_blockx_218 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_218_in_do), .start(_seach_blockx_218_start), .goal(_seach_blockx_218_goal), .data_out(_seach_blockx_218_data_out), .map_block(_seach_blockx_218_map_block), .now(_seach_blockx_218_now));
seach_block seach_blockx_217 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_217_in_do), .start(_seach_blockx_217_start), .goal(_seach_blockx_217_goal), .data_out(_seach_blockx_217_data_out), .map_block(_seach_blockx_217_map_block), .now(_seach_blockx_217_now));
seach_block seach_blockx_216 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_216_in_do), .start(_seach_blockx_216_start), .goal(_seach_blockx_216_goal), .data_out(_seach_blockx_216_data_out), .map_block(_seach_blockx_216_map_block), .now(_seach_blockx_216_now));
seach_block seach_blockx_215 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_215_in_do), .start(_seach_blockx_215_start), .goal(_seach_blockx_215_goal), .data_out(_seach_blockx_215_data_out), .map_block(_seach_blockx_215_map_block), .now(_seach_blockx_215_now));
seach_block seach_blockx_214 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_214_in_do), .start(_seach_blockx_214_start), .goal(_seach_blockx_214_goal), .data_out(_seach_blockx_214_data_out), .map_block(_seach_blockx_214_map_block), .now(_seach_blockx_214_now));
seach_block seach_blockx_213 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_213_in_do), .start(_seach_blockx_213_start), .goal(_seach_blockx_213_goal), .data_out(_seach_blockx_213_data_out), .map_block(_seach_blockx_213_map_block), .now(_seach_blockx_213_now));
seach_block seach_blockx_212 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_212_in_do), .start(_seach_blockx_212_start), .goal(_seach_blockx_212_goal), .data_out(_seach_blockx_212_data_out), .map_block(_seach_blockx_212_map_block), .now(_seach_blockx_212_now));
seach_block seach_blockx_211 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_211_in_do), .start(_seach_blockx_211_start), .goal(_seach_blockx_211_goal), .data_out(_seach_blockx_211_data_out), .map_block(_seach_blockx_211_map_block), .now(_seach_blockx_211_now));
seach_block seach_blockx_210 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_210_in_do), .start(_seach_blockx_210_start), .goal(_seach_blockx_210_goal), .data_out(_seach_blockx_210_data_out), .map_block(_seach_blockx_210_map_block), .now(_seach_blockx_210_now));
seach_block seach_blockx_209 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_209_in_do), .start(_seach_blockx_209_start), .goal(_seach_blockx_209_goal), .data_out(_seach_blockx_209_data_out), .map_block(_seach_blockx_209_map_block), .now(_seach_blockx_209_now));
seach_block seach_blockx_208 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_208_in_do), .start(_seach_blockx_208_start), .goal(_seach_blockx_208_goal), .data_out(_seach_blockx_208_data_out), .map_block(_seach_blockx_208_map_block), .now(_seach_blockx_208_now));
seach_block seach_blockx_207 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_207_in_do), .start(_seach_blockx_207_start), .goal(_seach_blockx_207_goal), .data_out(_seach_blockx_207_data_out), .map_block(_seach_blockx_207_map_block), .now(_seach_blockx_207_now));
seach_block seach_blockx_206 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_206_in_do), .start(_seach_blockx_206_start), .goal(_seach_blockx_206_goal), .data_out(_seach_blockx_206_data_out), .map_block(_seach_blockx_206_map_block), .now(_seach_blockx_206_now));
seach_block seach_blockx_205 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_205_in_do), .start(_seach_blockx_205_start), .goal(_seach_blockx_205_goal), .data_out(_seach_blockx_205_data_out), .map_block(_seach_blockx_205_map_block), .now(_seach_blockx_205_now));
seach_block seach_blockx_204 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_204_in_do), .start(_seach_blockx_204_start), .goal(_seach_blockx_204_goal), .data_out(_seach_blockx_204_data_out), .map_block(_seach_blockx_204_map_block), .now(_seach_blockx_204_now));
seach_block seach_blockx_203 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_203_in_do), .start(_seach_blockx_203_start), .goal(_seach_blockx_203_goal), .data_out(_seach_blockx_203_data_out), .map_block(_seach_blockx_203_map_block), .now(_seach_blockx_203_now));
seach_block seach_blockx_202 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_202_in_do), .start(_seach_blockx_202_start), .goal(_seach_blockx_202_goal), .data_out(_seach_blockx_202_data_out), .map_block(_seach_blockx_202_map_block), .now(_seach_blockx_202_now));
seach_block seach_blockx_201 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_201_in_do), .start(_seach_blockx_201_start), .goal(_seach_blockx_201_goal), .data_out(_seach_blockx_201_data_out), .map_block(_seach_blockx_201_map_block), .now(_seach_blockx_201_now));
seach_block seach_blockx_200 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_200_in_do), .start(_seach_blockx_200_start), .goal(_seach_blockx_200_goal), .data_out(_seach_blockx_200_data_out), .map_block(_seach_blockx_200_map_block), .now(_seach_blockx_200_now));
seach_block seach_blockx_199 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_199_in_do), .start(_seach_blockx_199_start), .goal(_seach_blockx_199_goal), .data_out(_seach_blockx_199_data_out), .map_block(_seach_blockx_199_map_block), .now(_seach_blockx_199_now));
seach_block seach_blockx_198 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_198_in_do), .start(_seach_blockx_198_start), .goal(_seach_blockx_198_goal), .data_out(_seach_blockx_198_data_out), .map_block(_seach_blockx_198_map_block), .now(_seach_blockx_198_now));
seach_block seach_blockx_197 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_197_in_do), .start(_seach_blockx_197_start), .goal(_seach_blockx_197_goal), .data_out(_seach_blockx_197_data_out), .map_block(_seach_blockx_197_map_block), .now(_seach_blockx_197_now));
seach_block seach_blockx_196 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_196_in_do), .start(_seach_blockx_196_start), .goal(_seach_blockx_196_goal), .data_out(_seach_blockx_196_data_out), .map_block(_seach_blockx_196_map_block), .now(_seach_blockx_196_now));
seach_block seach_blockx_195 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_195_in_do), .start(_seach_blockx_195_start), .goal(_seach_blockx_195_goal), .data_out(_seach_blockx_195_data_out), .map_block(_seach_blockx_195_map_block), .now(_seach_blockx_195_now));
seach_block seach_blockx_194 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_194_in_do), .start(_seach_blockx_194_start), .goal(_seach_blockx_194_goal), .data_out(_seach_blockx_194_data_out), .map_block(_seach_blockx_194_map_block), .now(_seach_blockx_194_now));
seach_block seach_blockx_193 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_193_in_do), .start(_seach_blockx_193_start), .goal(_seach_blockx_193_goal), .data_out(_seach_blockx_193_data_out), .map_block(_seach_blockx_193_map_block), .now(_seach_blockx_193_now));
seach_block seach_blockx_192 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_192_in_do), .start(_seach_blockx_192_start), .goal(_seach_blockx_192_goal), .data_out(_seach_blockx_192_data_out), .map_block(_seach_blockx_192_map_block), .now(_seach_blockx_192_now));
seach_block seach_blockx_191 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_191_in_do), .start(_seach_blockx_191_start), .goal(_seach_blockx_191_goal), .data_out(_seach_blockx_191_data_out), .map_block(_seach_blockx_191_map_block), .now(_seach_blockx_191_now));
seach_block seach_blockx_190 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_190_in_do), .start(_seach_blockx_190_start), .goal(_seach_blockx_190_goal), .data_out(_seach_blockx_190_data_out), .map_block(_seach_blockx_190_map_block), .now(_seach_blockx_190_now));
seach_block seach_blockx_189 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_189_in_do), .start(_seach_blockx_189_start), .goal(_seach_blockx_189_goal), .data_out(_seach_blockx_189_data_out), .map_block(_seach_blockx_189_map_block), .now(_seach_blockx_189_now));
seach_block seach_blockx_188 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_188_in_do), .start(_seach_blockx_188_start), .goal(_seach_blockx_188_goal), .data_out(_seach_blockx_188_data_out), .map_block(_seach_blockx_188_map_block), .now(_seach_blockx_188_now));
seach_block seach_blockx_187 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_187_in_do), .start(_seach_blockx_187_start), .goal(_seach_blockx_187_goal), .data_out(_seach_blockx_187_data_out), .map_block(_seach_blockx_187_map_block), .now(_seach_blockx_187_now));
seach_block seach_blockx_186 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_186_in_do), .start(_seach_blockx_186_start), .goal(_seach_blockx_186_goal), .data_out(_seach_blockx_186_data_out), .map_block(_seach_blockx_186_map_block), .now(_seach_blockx_186_now));
seach_block seach_blockx_185 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_185_in_do), .start(_seach_blockx_185_start), .goal(_seach_blockx_185_goal), .data_out(_seach_blockx_185_data_out), .map_block(_seach_blockx_185_map_block), .now(_seach_blockx_185_now));
seach_block seach_blockx_184 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_184_in_do), .start(_seach_blockx_184_start), .goal(_seach_blockx_184_goal), .data_out(_seach_blockx_184_data_out), .map_block(_seach_blockx_184_map_block), .now(_seach_blockx_184_now));
seach_block seach_blockx_183 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_183_in_do), .start(_seach_blockx_183_start), .goal(_seach_blockx_183_goal), .data_out(_seach_blockx_183_data_out), .map_block(_seach_blockx_183_map_block), .now(_seach_blockx_183_now));
seach_block seach_blockx_182 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_182_in_do), .start(_seach_blockx_182_start), .goal(_seach_blockx_182_goal), .data_out(_seach_blockx_182_data_out), .map_block(_seach_blockx_182_map_block), .now(_seach_blockx_182_now));
seach_block seach_blockx_181 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_181_in_do), .start(_seach_blockx_181_start), .goal(_seach_blockx_181_goal), .data_out(_seach_blockx_181_data_out), .map_block(_seach_blockx_181_map_block), .now(_seach_blockx_181_now));
seach_block seach_blockx_180 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_180_in_do), .start(_seach_blockx_180_start), .goal(_seach_blockx_180_goal), .data_out(_seach_blockx_180_data_out), .map_block(_seach_blockx_180_map_block), .now(_seach_blockx_180_now));
seach_block seach_blockx_179 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_179_in_do), .start(_seach_blockx_179_start), .goal(_seach_blockx_179_goal), .data_out(_seach_blockx_179_data_out), .map_block(_seach_blockx_179_map_block), .now(_seach_blockx_179_now));
seach_block seach_blockx_178 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_178_in_do), .start(_seach_blockx_178_start), .goal(_seach_blockx_178_goal), .data_out(_seach_blockx_178_data_out), .map_block(_seach_blockx_178_map_block), .now(_seach_blockx_178_now));
seach_block seach_blockx_177 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_177_in_do), .start(_seach_blockx_177_start), .goal(_seach_blockx_177_goal), .data_out(_seach_blockx_177_data_out), .map_block(_seach_blockx_177_map_block), .now(_seach_blockx_177_now));
seach_block seach_blockx_176 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_176_in_do), .start(_seach_blockx_176_start), .goal(_seach_blockx_176_goal), .data_out(_seach_blockx_176_data_out), .map_block(_seach_blockx_176_map_block), .now(_seach_blockx_176_now));
seach_block seach_blockx_175 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_175_in_do), .start(_seach_blockx_175_start), .goal(_seach_blockx_175_goal), .data_out(_seach_blockx_175_data_out), .map_block(_seach_blockx_175_map_block), .now(_seach_blockx_175_now));
seach_block seach_blockx_174 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_174_in_do), .start(_seach_blockx_174_start), .goal(_seach_blockx_174_goal), .data_out(_seach_blockx_174_data_out), .map_block(_seach_blockx_174_map_block), .now(_seach_blockx_174_now));
seach_block seach_blockx_173 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_173_in_do), .start(_seach_blockx_173_start), .goal(_seach_blockx_173_goal), .data_out(_seach_blockx_173_data_out), .map_block(_seach_blockx_173_map_block), .now(_seach_blockx_173_now));
seach_block seach_blockx_172 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_172_in_do), .start(_seach_blockx_172_start), .goal(_seach_blockx_172_goal), .data_out(_seach_blockx_172_data_out), .map_block(_seach_blockx_172_map_block), .now(_seach_blockx_172_now));
seach_block seach_blockx_171 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_171_in_do), .start(_seach_blockx_171_start), .goal(_seach_blockx_171_goal), .data_out(_seach_blockx_171_data_out), .map_block(_seach_blockx_171_map_block), .now(_seach_blockx_171_now));
seach_block seach_blockx_170 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_170_in_do), .start(_seach_blockx_170_start), .goal(_seach_blockx_170_goal), .data_out(_seach_blockx_170_data_out), .map_block(_seach_blockx_170_map_block), .now(_seach_blockx_170_now));
seach_block seach_blockx_169 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_169_in_do), .start(_seach_blockx_169_start), .goal(_seach_blockx_169_goal), .data_out(_seach_blockx_169_data_out), .map_block(_seach_blockx_169_map_block), .now(_seach_blockx_169_now));
seach_block seach_blockx_168 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_168_in_do), .start(_seach_blockx_168_start), .goal(_seach_blockx_168_goal), .data_out(_seach_blockx_168_data_out), .map_block(_seach_blockx_168_map_block), .now(_seach_blockx_168_now));
seach_block seach_blockx_167 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_167_in_do), .start(_seach_blockx_167_start), .goal(_seach_blockx_167_goal), .data_out(_seach_blockx_167_data_out), .map_block(_seach_blockx_167_map_block), .now(_seach_blockx_167_now));
seach_block seach_blockx_166 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_166_in_do), .start(_seach_blockx_166_start), .goal(_seach_blockx_166_goal), .data_out(_seach_blockx_166_data_out), .map_block(_seach_blockx_166_map_block), .now(_seach_blockx_166_now));
seach_block seach_blockx_165 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_165_in_do), .start(_seach_blockx_165_start), .goal(_seach_blockx_165_goal), .data_out(_seach_blockx_165_data_out), .map_block(_seach_blockx_165_map_block), .now(_seach_blockx_165_now));
seach_block seach_blockx_164 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_164_in_do), .start(_seach_blockx_164_start), .goal(_seach_blockx_164_goal), .data_out(_seach_blockx_164_data_out), .map_block(_seach_blockx_164_map_block), .now(_seach_blockx_164_now));
seach_block seach_blockx_163 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_163_in_do), .start(_seach_blockx_163_start), .goal(_seach_blockx_163_goal), .data_out(_seach_blockx_163_data_out), .map_block(_seach_blockx_163_map_block), .now(_seach_blockx_163_now));
seach_block seach_blockx_162 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_162_in_do), .start(_seach_blockx_162_start), .goal(_seach_blockx_162_goal), .data_out(_seach_blockx_162_data_out), .map_block(_seach_blockx_162_map_block), .now(_seach_blockx_162_now));
seach_block seach_blockx_161 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_161_in_do), .start(_seach_blockx_161_start), .goal(_seach_blockx_161_goal), .data_out(_seach_blockx_161_data_out), .map_block(_seach_blockx_161_map_block), .now(_seach_blockx_161_now));
seach_block seach_blockx_160 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_160_in_do), .start(_seach_blockx_160_start), .goal(_seach_blockx_160_goal), .data_out(_seach_blockx_160_data_out), .map_block(_seach_blockx_160_map_block), .now(_seach_blockx_160_now));
seach_block seach_blockx_159 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_159_in_do), .start(_seach_blockx_159_start), .goal(_seach_blockx_159_goal), .data_out(_seach_blockx_159_data_out), .map_block(_seach_blockx_159_map_block), .now(_seach_blockx_159_now));
seach_block seach_blockx_158 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_158_in_do), .start(_seach_blockx_158_start), .goal(_seach_blockx_158_goal), .data_out(_seach_blockx_158_data_out), .map_block(_seach_blockx_158_map_block), .now(_seach_blockx_158_now));
seach_block seach_blockx_157 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_157_in_do), .start(_seach_blockx_157_start), .goal(_seach_blockx_157_goal), .data_out(_seach_blockx_157_data_out), .map_block(_seach_blockx_157_map_block), .now(_seach_blockx_157_now));
seach_block seach_blockx_156 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_156_in_do), .start(_seach_blockx_156_start), .goal(_seach_blockx_156_goal), .data_out(_seach_blockx_156_data_out), .map_block(_seach_blockx_156_map_block), .now(_seach_blockx_156_now));
seach_block seach_blockx_155 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_155_in_do), .start(_seach_blockx_155_start), .goal(_seach_blockx_155_goal), .data_out(_seach_blockx_155_data_out), .map_block(_seach_blockx_155_map_block), .now(_seach_blockx_155_now));
seach_block seach_blockx_154 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_154_in_do), .start(_seach_blockx_154_start), .goal(_seach_blockx_154_goal), .data_out(_seach_blockx_154_data_out), .map_block(_seach_blockx_154_map_block), .now(_seach_blockx_154_now));
seach_block seach_blockx_153 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_153_in_do), .start(_seach_blockx_153_start), .goal(_seach_blockx_153_goal), .data_out(_seach_blockx_153_data_out), .map_block(_seach_blockx_153_map_block), .now(_seach_blockx_153_now));
seach_block seach_blockx_152 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_152_in_do), .start(_seach_blockx_152_start), .goal(_seach_blockx_152_goal), .data_out(_seach_blockx_152_data_out), .map_block(_seach_blockx_152_map_block), .now(_seach_blockx_152_now));
seach_block seach_blockx_151 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_151_in_do), .start(_seach_blockx_151_start), .goal(_seach_blockx_151_goal), .data_out(_seach_blockx_151_data_out), .map_block(_seach_blockx_151_map_block), .now(_seach_blockx_151_now));
seach_block seach_blockx_150 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_150_in_do), .start(_seach_blockx_150_start), .goal(_seach_blockx_150_goal), .data_out(_seach_blockx_150_data_out), .map_block(_seach_blockx_150_map_block), .now(_seach_blockx_150_now));
seach_block seach_blockx_149 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_149_in_do), .start(_seach_blockx_149_start), .goal(_seach_blockx_149_goal), .data_out(_seach_blockx_149_data_out), .map_block(_seach_blockx_149_map_block), .now(_seach_blockx_149_now));
seach_block seach_blockx_148 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_148_in_do), .start(_seach_blockx_148_start), .goal(_seach_blockx_148_goal), .data_out(_seach_blockx_148_data_out), .map_block(_seach_blockx_148_map_block), .now(_seach_blockx_148_now));
seach_block seach_blockx_147 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_147_in_do), .start(_seach_blockx_147_start), .goal(_seach_blockx_147_goal), .data_out(_seach_blockx_147_data_out), .map_block(_seach_blockx_147_map_block), .now(_seach_blockx_147_now));
seach_block seach_blockx_146 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_146_in_do), .start(_seach_blockx_146_start), .goal(_seach_blockx_146_goal), .data_out(_seach_blockx_146_data_out), .map_block(_seach_blockx_146_map_block), .now(_seach_blockx_146_now));
seach_block seach_blockx_145 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_145_in_do), .start(_seach_blockx_145_start), .goal(_seach_blockx_145_goal), .data_out(_seach_blockx_145_data_out), .map_block(_seach_blockx_145_map_block), .now(_seach_blockx_145_now));
seach_block seach_blockx_144 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_144_in_do), .start(_seach_blockx_144_start), .goal(_seach_blockx_144_goal), .data_out(_seach_blockx_144_data_out), .map_block(_seach_blockx_144_map_block), .now(_seach_blockx_144_now));
seach_block seach_blockx_143 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_143_in_do), .start(_seach_blockx_143_start), .goal(_seach_blockx_143_goal), .data_out(_seach_blockx_143_data_out), .map_block(_seach_blockx_143_map_block), .now(_seach_blockx_143_now));
seach_block seach_blockx_142 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_142_in_do), .start(_seach_blockx_142_start), .goal(_seach_blockx_142_goal), .data_out(_seach_blockx_142_data_out), .map_block(_seach_blockx_142_map_block), .now(_seach_blockx_142_now));
seach_block seach_blockx_141 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_141_in_do), .start(_seach_blockx_141_start), .goal(_seach_blockx_141_goal), .data_out(_seach_blockx_141_data_out), .map_block(_seach_blockx_141_map_block), .now(_seach_blockx_141_now));
seach_block seach_blockx_140 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_140_in_do), .start(_seach_blockx_140_start), .goal(_seach_blockx_140_goal), .data_out(_seach_blockx_140_data_out), .map_block(_seach_blockx_140_map_block), .now(_seach_blockx_140_now));
seach_block seach_blockx_139 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_139_in_do), .start(_seach_blockx_139_start), .goal(_seach_blockx_139_goal), .data_out(_seach_blockx_139_data_out), .map_block(_seach_blockx_139_map_block), .now(_seach_blockx_139_now));
seach_block seach_blockx_138 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_138_in_do), .start(_seach_blockx_138_start), .goal(_seach_blockx_138_goal), .data_out(_seach_blockx_138_data_out), .map_block(_seach_blockx_138_map_block), .now(_seach_blockx_138_now));
seach_block seach_blockx_137 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_137_in_do), .start(_seach_blockx_137_start), .goal(_seach_blockx_137_goal), .data_out(_seach_blockx_137_data_out), .map_block(_seach_blockx_137_map_block), .now(_seach_blockx_137_now));
seach_block seach_blockx_136 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_136_in_do), .start(_seach_blockx_136_start), .goal(_seach_blockx_136_goal), .data_out(_seach_blockx_136_data_out), .map_block(_seach_blockx_136_map_block), .now(_seach_blockx_136_now));
seach_block seach_blockx_135 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_135_in_do), .start(_seach_blockx_135_start), .goal(_seach_blockx_135_goal), .data_out(_seach_blockx_135_data_out), .map_block(_seach_blockx_135_map_block), .now(_seach_blockx_135_now));
seach_block seach_blockx_134 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_134_in_do), .start(_seach_blockx_134_start), .goal(_seach_blockx_134_goal), .data_out(_seach_blockx_134_data_out), .map_block(_seach_blockx_134_map_block), .now(_seach_blockx_134_now));
seach_block seach_blockx_133 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_133_in_do), .start(_seach_blockx_133_start), .goal(_seach_blockx_133_goal), .data_out(_seach_blockx_133_data_out), .map_block(_seach_blockx_133_map_block), .now(_seach_blockx_133_now));
seach_block seach_blockx_132 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_132_in_do), .start(_seach_blockx_132_start), .goal(_seach_blockx_132_goal), .data_out(_seach_blockx_132_data_out), .map_block(_seach_blockx_132_map_block), .now(_seach_blockx_132_now));
seach_block seach_blockx_131 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_131_in_do), .start(_seach_blockx_131_start), .goal(_seach_blockx_131_goal), .data_out(_seach_blockx_131_data_out), .map_block(_seach_blockx_131_map_block), .now(_seach_blockx_131_now));
seach_block seach_blockx_130 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_130_in_do), .start(_seach_blockx_130_start), .goal(_seach_blockx_130_goal), .data_out(_seach_blockx_130_data_out), .map_block(_seach_blockx_130_map_block), .now(_seach_blockx_130_now));
seach_block seach_blockx_129 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_129_in_do), .start(_seach_blockx_129_start), .goal(_seach_blockx_129_goal), .data_out(_seach_blockx_129_data_out), .map_block(_seach_blockx_129_map_block), .now(_seach_blockx_129_now));
seach_block seach_blockx_128 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_128_in_do), .start(_seach_blockx_128_start), .goal(_seach_blockx_128_goal), .data_out(_seach_blockx_128_data_out), .map_block(_seach_blockx_128_map_block), .now(_seach_blockx_128_now));
seach_block seach_blockx_127 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_127_in_do), .start(_seach_blockx_127_start), .goal(_seach_blockx_127_goal), .data_out(_seach_blockx_127_data_out), .map_block(_seach_blockx_127_map_block), .now(_seach_blockx_127_now));
seach_block seach_blockx_126 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_126_in_do), .start(_seach_blockx_126_start), .goal(_seach_blockx_126_goal), .data_out(_seach_blockx_126_data_out), .map_block(_seach_blockx_126_map_block), .now(_seach_blockx_126_now));
seach_block seach_blockx_125 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_125_in_do), .start(_seach_blockx_125_start), .goal(_seach_blockx_125_goal), .data_out(_seach_blockx_125_data_out), .map_block(_seach_blockx_125_map_block), .now(_seach_blockx_125_now));
seach_block seach_blockx_124 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_124_in_do), .start(_seach_blockx_124_start), .goal(_seach_blockx_124_goal), .data_out(_seach_blockx_124_data_out), .map_block(_seach_blockx_124_map_block), .now(_seach_blockx_124_now));
seach_block seach_blockx_123 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_123_in_do), .start(_seach_blockx_123_start), .goal(_seach_blockx_123_goal), .data_out(_seach_blockx_123_data_out), .map_block(_seach_blockx_123_map_block), .now(_seach_blockx_123_now));
seach_block seach_blockx_122 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_122_in_do), .start(_seach_blockx_122_start), .goal(_seach_blockx_122_goal), .data_out(_seach_blockx_122_data_out), .map_block(_seach_blockx_122_map_block), .now(_seach_blockx_122_now));
seach_block seach_blockx_121 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_121_in_do), .start(_seach_blockx_121_start), .goal(_seach_blockx_121_goal), .data_out(_seach_blockx_121_data_out), .map_block(_seach_blockx_121_map_block), .now(_seach_blockx_121_now));
seach_block seach_blockx_120 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_120_in_do), .start(_seach_blockx_120_start), .goal(_seach_blockx_120_goal), .data_out(_seach_blockx_120_data_out), .map_block(_seach_blockx_120_map_block), .now(_seach_blockx_120_now));
seach_block seach_blockx_119 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_119_in_do), .start(_seach_blockx_119_start), .goal(_seach_blockx_119_goal), .data_out(_seach_blockx_119_data_out), .map_block(_seach_blockx_119_map_block), .now(_seach_blockx_119_now));
seach_block seach_blockx_118 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_118_in_do), .start(_seach_blockx_118_start), .goal(_seach_blockx_118_goal), .data_out(_seach_blockx_118_data_out), .map_block(_seach_blockx_118_map_block), .now(_seach_blockx_118_now));
seach_block seach_blockx_117 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_117_in_do), .start(_seach_blockx_117_start), .goal(_seach_blockx_117_goal), .data_out(_seach_blockx_117_data_out), .map_block(_seach_blockx_117_map_block), .now(_seach_blockx_117_now));
seach_block seach_blockx_116 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_116_in_do), .start(_seach_blockx_116_start), .goal(_seach_blockx_116_goal), .data_out(_seach_blockx_116_data_out), .map_block(_seach_blockx_116_map_block), .now(_seach_blockx_116_now));
seach_block seach_blockx_115 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_115_in_do), .start(_seach_blockx_115_start), .goal(_seach_blockx_115_goal), .data_out(_seach_blockx_115_data_out), .map_block(_seach_blockx_115_map_block), .now(_seach_blockx_115_now));
seach_block seach_blockx_114 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_114_in_do), .start(_seach_blockx_114_start), .goal(_seach_blockx_114_goal), .data_out(_seach_blockx_114_data_out), .map_block(_seach_blockx_114_map_block), .now(_seach_blockx_114_now));
seach_block seach_blockx_113 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_113_in_do), .start(_seach_blockx_113_start), .goal(_seach_blockx_113_goal), .data_out(_seach_blockx_113_data_out), .map_block(_seach_blockx_113_map_block), .now(_seach_blockx_113_now));
seach_block seach_blockx_112 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_112_in_do), .start(_seach_blockx_112_start), .goal(_seach_blockx_112_goal), .data_out(_seach_blockx_112_data_out), .map_block(_seach_blockx_112_map_block), .now(_seach_blockx_112_now));
seach_block seach_blockx_111 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_111_in_do), .start(_seach_blockx_111_start), .goal(_seach_blockx_111_goal), .data_out(_seach_blockx_111_data_out), .map_block(_seach_blockx_111_map_block), .now(_seach_blockx_111_now));
seach_block seach_blockx_110 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_110_in_do), .start(_seach_blockx_110_start), .goal(_seach_blockx_110_goal), .data_out(_seach_blockx_110_data_out), .map_block(_seach_blockx_110_map_block), .now(_seach_blockx_110_now));
seach_block seach_blockx_109 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_109_in_do), .start(_seach_blockx_109_start), .goal(_seach_blockx_109_goal), .data_out(_seach_blockx_109_data_out), .map_block(_seach_blockx_109_map_block), .now(_seach_blockx_109_now));
seach_block seach_blockx_108 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_108_in_do), .start(_seach_blockx_108_start), .goal(_seach_blockx_108_goal), .data_out(_seach_blockx_108_data_out), .map_block(_seach_blockx_108_map_block), .now(_seach_blockx_108_now));
seach_block seach_blockx_107 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_107_in_do), .start(_seach_blockx_107_start), .goal(_seach_blockx_107_goal), .data_out(_seach_blockx_107_data_out), .map_block(_seach_blockx_107_map_block), .now(_seach_blockx_107_now));
seach_block seach_blockx_106 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_106_in_do), .start(_seach_blockx_106_start), .goal(_seach_blockx_106_goal), .data_out(_seach_blockx_106_data_out), .map_block(_seach_blockx_106_map_block), .now(_seach_blockx_106_now));
seach_block seach_blockx_105 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_105_in_do), .start(_seach_blockx_105_start), .goal(_seach_blockx_105_goal), .data_out(_seach_blockx_105_data_out), .map_block(_seach_blockx_105_map_block), .now(_seach_blockx_105_now));
seach_block seach_blockx_104 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_104_in_do), .start(_seach_blockx_104_start), .goal(_seach_blockx_104_goal), .data_out(_seach_blockx_104_data_out), .map_block(_seach_blockx_104_map_block), .now(_seach_blockx_104_now));
seach_block seach_blockx_103 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_103_in_do), .start(_seach_blockx_103_start), .goal(_seach_blockx_103_goal), .data_out(_seach_blockx_103_data_out), .map_block(_seach_blockx_103_map_block), .now(_seach_blockx_103_now));
seach_block seach_blockx_102 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_102_in_do), .start(_seach_blockx_102_start), .goal(_seach_blockx_102_goal), .data_out(_seach_blockx_102_data_out), .map_block(_seach_blockx_102_map_block), .now(_seach_blockx_102_now));
seach_block seach_blockx_101 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_101_in_do), .start(_seach_blockx_101_start), .goal(_seach_blockx_101_goal), .data_out(_seach_blockx_101_data_out), .map_block(_seach_blockx_101_map_block), .now(_seach_blockx_101_now));
seach_block seach_blockx_100 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_100_in_do), .start(_seach_blockx_100_start), .goal(_seach_blockx_100_goal), .data_out(_seach_blockx_100_data_out), .map_block(_seach_blockx_100_map_block), .now(_seach_blockx_100_now));
seach_block seach_blockx_99 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_99_in_do), .start(_seach_blockx_99_start), .goal(_seach_blockx_99_goal), .data_out(_seach_blockx_99_data_out), .map_block(_seach_blockx_99_map_block), .now(_seach_blockx_99_now));
seach_block seach_blockx_98 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_98_in_do), .start(_seach_blockx_98_start), .goal(_seach_blockx_98_goal), .data_out(_seach_blockx_98_data_out), .map_block(_seach_blockx_98_map_block), .now(_seach_blockx_98_now));
seach_block seach_blockx_97 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_97_in_do), .start(_seach_blockx_97_start), .goal(_seach_blockx_97_goal), .data_out(_seach_blockx_97_data_out), .map_block(_seach_blockx_97_map_block), .now(_seach_blockx_97_now));
seach_block seach_blockx_96 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_96_in_do), .start(_seach_blockx_96_start), .goal(_seach_blockx_96_goal), .data_out(_seach_blockx_96_data_out), .map_block(_seach_blockx_96_map_block), .now(_seach_blockx_96_now));
seach_block seach_blockx_95 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_95_in_do), .start(_seach_blockx_95_start), .goal(_seach_blockx_95_goal), .data_out(_seach_blockx_95_data_out), .map_block(_seach_blockx_95_map_block), .now(_seach_blockx_95_now));
seach_block seach_blockx_94 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_94_in_do), .start(_seach_blockx_94_start), .goal(_seach_blockx_94_goal), .data_out(_seach_blockx_94_data_out), .map_block(_seach_blockx_94_map_block), .now(_seach_blockx_94_now));
seach_block seach_blockx_93 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_93_in_do), .start(_seach_blockx_93_start), .goal(_seach_blockx_93_goal), .data_out(_seach_blockx_93_data_out), .map_block(_seach_blockx_93_map_block), .now(_seach_blockx_93_now));
seach_block seach_blockx_92 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_92_in_do), .start(_seach_blockx_92_start), .goal(_seach_blockx_92_goal), .data_out(_seach_blockx_92_data_out), .map_block(_seach_blockx_92_map_block), .now(_seach_blockx_92_now));
seach_block seach_blockx_91 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_91_in_do), .start(_seach_blockx_91_start), .goal(_seach_blockx_91_goal), .data_out(_seach_blockx_91_data_out), .map_block(_seach_blockx_91_map_block), .now(_seach_blockx_91_now));
seach_block seach_blockx_90 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_90_in_do), .start(_seach_blockx_90_start), .goal(_seach_blockx_90_goal), .data_out(_seach_blockx_90_data_out), .map_block(_seach_blockx_90_map_block), .now(_seach_blockx_90_now));
seach_block seach_blockx_89 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_89_in_do), .start(_seach_blockx_89_start), .goal(_seach_blockx_89_goal), .data_out(_seach_blockx_89_data_out), .map_block(_seach_blockx_89_map_block), .now(_seach_blockx_89_now));
seach_block seach_blockx_88 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_88_in_do), .start(_seach_blockx_88_start), .goal(_seach_blockx_88_goal), .data_out(_seach_blockx_88_data_out), .map_block(_seach_blockx_88_map_block), .now(_seach_blockx_88_now));
seach_block seach_blockx_87 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_87_in_do), .start(_seach_blockx_87_start), .goal(_seach_blockx_87_goal), .data_out(_seach_blockx_87_data_out), .map_block(_seach_blockx_87_map_block), .now(_seach_blockx_87_now));
seach_block seach_blockx_86 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_86_in_do), .start(_seach_blockx_86_start), .goal(_seach_blockx_86_goal), .data_out(_seach_blockx_86_data_out), .map_block(_seach_blockx_86_map_block), .now(_seach_blockx_86_now));
seach_block seach_blockx_85 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_85_in_do), .start(_seach_blockx_85_start), .goal(_seach_blockx_85_goal), .data_out(_seach_blockx_85_data_out), .map_block(_seach_blockx_85_map_block), .now(_seach_blockx_85_now));
seach_block seach_blockx_84 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_84_in_do), .start(_seach_blockx_84_start), .goal(_seach_blockx_84_goal), .data_out(_seach_blockx_84_data_out), .map_block(_seach_blockx_84_map_block), .now(_seach_blockx_84_now));
seach_block seach_blockx_83 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_83_in_do), .start(_seach_blockx_83_start), .goal(_seach_blockx_83_goal), .data_out(_seach_blockx_83_data_out), .map_block(_seach_blockx_83_map_block), .now(_seach_blockx_83_now));
seach_block seach_blockx_82 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_82_in_do), .start(_seach_blockx_82_start), .goal(_seach_blockx_82_goal), .data_out(_seach_blockx_82_data_out), .map_block(_seach_blockx_82_map_block), .now(_seach_blockx_82_now));
seach_block seach_blockx_81 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_81_in_do), .start(_seach_blockx_81_start), .goal(_seach_blockx_81_goal), .data_out(_seach_blockx_81_data_out), .map_block(_seach_blockx_81_map_block), .now(_seach_blockx_81_now));
seach_block seach_blockx_80 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_80_in_do), .start(_seach_blockx_80_start), .goal(_seach_blockx_80_goal), .data_out(_seach_blockx_80_data_out), .map_block(_seach_blockx_80_map_block), .now(_seach_blockx_80_now));
seach_block seach_blockx_79 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_79_in_do), .start(_seach_blockx_79_start), .goal(_seach_blockx_79_goal), .data_out(_seach_blockx_79_data_out), .map_block(_seach_blockx_79_map_block), .now(_seach_blockx_79_now));
seach_block seach_blockx_78 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_78_in_do), .start(_seach_blockx_78_start), .goal(_seach_blockx_78_goal), .data_out(_seach_blockx_78_data_out), .map_block(_seach_blockx_78_map_block), .now(_seach_blockx_78_now));
seach_block seach_blockx_77 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_77_in_do), .start(_seach_blockx_77_start), .goal(_seach_blockx_77_goal), .data_out(_seach_blockx_77_data_out), .map_block(_seach_blockx_77_map_block), .now(_seach_blockx_77_now));
seach_block seach_blockx_76 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_76_in_do), .start(_seach_blockx_76_start), .goal(_seach_blockx_76_goal), .data_out(_seach_blockx_76_data_out), .map_block(_seach_blockx_76_map_block), .now(_seach_blockx_76_now));
seach_block seach_blockx_75 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_75_in_do), .start(_seach_blockx_75_start), .goal(_seach_blockx_75_goal), .data_out(_seach_blockx_75_data_out), .map_block(_seach_blockx_75_map_block), .now(_seach_blockx_75_now));
seach_block seach_blockx_74 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_74_in_do), .start(_seach_blockx_74_start), .goal(_seach_blockx_74_goal), .data_out(_seach_blockx_74_data_out), .map_block(_seach_blockx_74_map_block), .now(_seach_blockx_74_now));
seach_block seach_blockx_73 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_73_in_do), .start(_seach_blockx_73_start), .goal(_seach_blockx_73_goal), .data_out(_seach_blockx_73_data_out), .map_block(_seach_blockx_73_map_block), .now(_seach_blockx_73_now));
seach_block seach_blockx_72 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_72_in_do), .start(_seach_blockx_72_start), .goal(_seach_blockx_72_goal), .data_out(_seach_blockx_72_data_out), .map_block(_seach_blockx_72_map_block), .now(_seach_blockx_72_now));
seach_block seach_blockx_71 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_71_in_do), .start(_seach_blockx_71_start), .goal(_seach_blockx_71_goal), .data_out(_seach_blockx_71_data_out), .map_block(_seach_blockx_71_map_block), .now(_seach_blockx_71_now));
seach_block seach_blockx_70 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_70_in_do), .start(_seach_blockx_70_start), .goal(_seach_blockx_70_goal), .data_out(_seach_blockx_70_data_out), .map_block(_seach_blockx_70_map_block), .now(_seach_blockx_70_now));
seach_block seach_blockx_69 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_69_in_do), .start(_seach_blockx_69_start), .goal(_seach_blockx_69_goal), .data_out(_seach_blockx_69_data_out), .map_block(_seach_blockx_69_map_block), .now(_seach_blockx_69_now));
seach_block seach_blockx_68 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_68_in_do), .start(_seach_blockx_68_start), .goal(_seach_blockx_68_goal), .data_out(_seach_blockx_68_data_out), .map_block(_seach_blockx_68_map_block), .now(_seach_blockx_68_now));
seach_block seach_blockx_67 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_67_in_do), .start(_seach_blockx_67_start), .goal(_seach_blockx_67_goal), .data_out(_seach_blockx_67_data_out), .map_block(_seach_blockx_67_map_block), .now(_seach_blockx_67_now));
seach_block seach_blockx_66 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_66_in_do), .start(_seach_blockx_66_start), .goal(_seach_blockx_66_goal), .data_out(_seach_blockx_66_data_out), .map_block(_seach_blockx_66_map_block), .now(_seach_blockx_66_now));
seach_block seach_blockx_65 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_65_in_do), .start(_seach_blockx_65_start), .goal(_seach_blockx_65_goal), .data_out(_seach_blockx_65_data_out), .map_block(_seach_blockx_65_map_block), .now(_seach_blockx_65_now));
seach_block seach_blockx_64 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_64_in_do), .start(_seach_blockx_64_start), .goal(_seach_blockx_64_goal), .data_out(_seach_blockx_64_data_out), .map_block(_seach_blockx_64_map_block), .now(_seach_blockx_64_now));
seach_block seach_blockx_63 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_63_in_do), .start(_seach_blockx_63_start), .goal(_seach_blockx_63_goal), .data_out(_seach_blockx_63_data_out), .map_block(_seach_blockx_63_map_block), .now(_seach_blockx_63_now));
seach_block seach_blockx_62 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_62_in_do), .start(_seach_blockx_62_start), .goal(_seach_blockx_62_goal), .data_out(_seach_blockx_62_data_out), .map_block(_seach_blockx_62_map_block), .now(_seach_blockx_62_now));
seach_block seach_blockx_61 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_61_in_do), .start(_seach_blockx_61_start), .goal(_seach_blockx_61_goal), .data_out(_seach_blockx_61_data_out), .map_block(_seach_blockx_61_map_block), .now(_seach_blockx_61_now));
seach_block seach_blockx_60 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_60_in_do), .start(_seach_blockx_60_start), .goal(_seach_blockx_60_goal), .data_out(_seach_blockx_60_data_out), .map_block(_seach_blockx_60_map_block), .now(_seach_blockx_60_now));
seach_block seach_blockx_59 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_59_in_do), .start(_seach_blockx_59_start), .goal(_seach_blockx_59_goal), .data_out(_seach_blockx_59_data_out), .map_block(_seach_blockx_59_map_block), .now(_seach_blockx_59_now));
seach_block seach_blockx_58 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_58_in_do), .start(_seach_blockx_58_start), .goal(_seach_blockx_58_goal), .data_out(_seach_blockx_58_data_out), .map_block(_seach_blockx_58_map_block), .now(_seach_blockx_58_now));
seach_block seach_blockx_57 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_57_in_do), .start(_seach_blockx_57_start), .goal(_seach_blockx_57_goal), .data_out(_seach_blockx_57_data_out), .map_block(_seach_blockx_57_map_block), .now(_seach_blockx_57_now));
seach_block seach_blockx_56 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_56_in_do), .start(_seach_blockx_56_start), .goal(_seach_blockx_56_goal), .data_out(_seach_blockx_56_data_out), .map_block(_seach_blockx_56_map_block), .now(_seach_blockx_56_now));
seach_block seach_blockx_55 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_55_in_do), .start(_seach_blockx_55_start), .goal(_seach_blockx_55_goal), .data_out(_seach_blockx_55_data_out), .map_block(_seach_blockx_55_map_block), .now(_seach_blockx_55_now));
seach_block seach_blockx_54 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_54_in_do), .start(_seach_blockx_54_start), .goal(_seach_blockx_54_goal), .data_out(_seach_blockx_54_data_out), .map_block(_seach_blockx_54_map_block), .now(_seach_blockx_54_now));
seach_block seach_blockx_53 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_53_in_do), .start(_seach_blockx_53_start), .goal(_seach_blockx_53_goal), .data_out(_seach_blockx_53_data_out), .map_block(_seach_blockx_53_map_block), .now(_seach_blockx_53_now));
seach_block seach_blockx_52 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_52_in_do), .start(_seach_blockx_52_start), .goal(_seach_blockx_52_goal), .data_out(_seach_blockx_52_data_out), .map_block(_seach_blockx_52_map_block), .now(_seach_blockx_52_now));
seach_block seach_blockx_51 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_51_in_do), .start(_seach_blockx_51_start), .goal(_seach_blockx_51_goal), .data_out(_seach_blockx_51_data_out), .map_block(_seach_blockx_51_map_block), .now(_seach_blockx_51_now));
seach_block seach_blockx_50 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_50_in_do), .start(_seach_blockx_50_start), .goal(_seach_blockx_50_goal), .data_out(_seach_blockx_50_data_out), .map_block(_seach_blockx_50_map_block), .now(_seach_blockx_50_now));
seach_block seach_blockx_49 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_49_in_do), .start(_seach_blockx_49_start), .goal(_seach_blockx_49_goal), .data_out(_seach_blockx_49_data_out), .map_block(_seach_blockx_49_map_block), .now(_seach_blockx_49_now));
seach_block seach_blockx_48 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_48_in_do), .start(_seach_blockx_48_start), .goal(_seach_blockx_48_goal), .data_out(_seach_blockx_48_data_out), .map_block(_seach_blockx_48_map_block), .now(_seach_blockx_48_now));
seach_block seach_blockx_47 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_47_in_do), .start(_seach_blockx_47_start), .goal(_seach_blockx_47_goal), .data_out(_seach_blockx_47_data_out), .map_block(_seach_blockx_47_map_block), .now(_seach_blockx_47_now));
seach_block seach_blockx_46 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_46_in_do), .start(_seach_blockx_46_start), .goal(_seach_blockx_46_goal), .data_out(_seach_blockx_46_data_out), .map_block(_seach_blockx_46_map_block), .now(_seach_blockx_46_now));
seach_block seach_blockx_45 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_45_in_do), .start(_seach_blockx_45_start), .goal(_seach_blockx_45_goal), .data_out(_seach_blockx_45_data_out), .map_block(_seach_blockx_45_map_block), .now(_seach_blockx_45_now));
seach_block seach_blockx_44 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_44_in_do), .start(_seach_blockx_44_start), .goal(_seach_blockx_44_goal), .data_out(_seach_blockx_44_data_out), .map_block(_seach_blockx_44_map_block), .now(_seach_blockx_44_now));
seach_block seach_blockx_43 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_43_in_do), .start(_seach_blockx_43_start), .goal(_seach_blockx_43_goal), .data_out(_seach_blockx_43_data_out), .map_block(_seach_blockx_43_map_block), .now(_seach_blockx_43_now));
seach_block seach_blockx_42 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_42_in_do), .start(_seach_blockx_42_start), .goal(_seach_blockx_42_goal), .data_out(_seach_blockx_42_data_out), .map_block(_seach_blockx_42_map_block), .now(_seach_blockx_42_now));
seach_block seach_blockx_41 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_41_in_do), .start(_seach_blockx_41_start), .goal(_seach_blockx_41_goal), .data_out(_seach_blockx_41_data_out), .map_block(_seach_blockx_41_map_block), .now(_seach_blockx_41_now));
seach_block seach_blockx_40 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_40_in_do), .start(_seach_blockx_40_start), .goal(_seach_blockx_40_goal), .data_out(_seach_blockx_40_data_out), .map_block(_seach_blockx_40_map_block), .now(_seach_blockx_40_now));
seach_block seach_blockx_39 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_39_in_do), .start(_seach_blockx_39_start), .goal(_seach_blockx_39_goal), .data_out(_seach_blockx_39_data_out), .map_block(_seach_blockx_39_map_block), .now(_seach_blockx_39_now));
seach_block seach_blockx_38 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_38_in_do), .start(_seach_blockx_38_start), .goal(_seach_blockx_38_goal), .data_out(_seach_blockx_38_data_out), .map_block(_seach_blockx_38_map_block), .now(_seach_blockx_38_now));
seach_block seach_blockx_37 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_37_in_do), .start(_seach_blockx_37_start), .goal(_seach_blockx_37_goal), .data_out(_seach_blockx_37_data_out), .map_block(_seach_blockx_37_map_block), .now(_seach_blockx_37_now));
seach_block seach_blockx_36 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_36_in_do), .start(_seach_blockx_36_start), .goal(_seach_blockx_36_goal), .data_out(_seach_blockx_36_data_out), .map_block(_seach_blockx_36_map_block), .now(_seach_blockx_36_now));
seach_block seach_blockx_35 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_35_in_do), .start(_seach_blockx_35_start), .goal(_seach_blockx_35_goal), .data_out(_seach_blockx_35_data_out), .map_block(_seach_blockx_35_map_block), .now(_seach_blockx_35_now));
seach_block seach_blockx_34 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_34_in_do), .start(_seach_blockx_34_start), .goal(_seach_blockx_34_goal), .data_out(_seach_blockx_34_data_out), .map_block(_seach_blockx_34_map_block), .now(_seach_blockx_34_now));
seach_block seach_blockx_33 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_33_in_do), .start(_seach_blockx_33_start), .goal(_seach_blockx_33_goal), .data_out(_seach_blockx_33_data_out), .map_block(_seach_blockx_33_map_block), .now(_seach_blockx_33_now));
seach_block seach_blockx_32 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_32_in_do), .start(_seach_blockx_32_start), .goal(_seach_blockx_32_goal), .data_out(_seach_blockx_32_data_out), .map_block(_seach_blockx_32_map_block), .now(_seach_blockx_32_now));
seach_block seach_blockx_31 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_31_in_do), .start(_seach_blockx_31_start), .goal(_seach_blockx_31_goal), .data_out(_seach_blockx_31_data_out), .map_block(_seach_blockx_31_map_block), .now(_seach_blockx_31_now));
seach_block seach_blockx_30 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_30_in_do), .start(_seach_blockx_30_start), .goal(_seach_blockx_30_goal), .data_out(_seach_blockx_30_data_out), .map_block(_seach_blockx_30_map_block), .now(_seach_blockx_30_now));
seach_block seach_blockx_29 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_29_in_do), .start(_seach_blockx_29_start), .goal(_seach_blockx_29_goal), .data_out(_seach_blockx_29_data_out), .map_block(_seach_blockx_29_map_block), .now(_seach_blockx_29_now));
seach_block seach_blockx_28 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_28_in_do), .start(_seach_blockx_28_start), .goal(_seach_blockx_28_goal), .data_out(_seach_blockx_28_data_out), .map_block(_seach_blockx_28_map_block), .now(_seach_blockx_28_now));
seach_block seach_blockx_27 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_27_in_do), .start(_seach_blockx_27_start), .goal(_seach_blockx_27_goal), .data_out(_seach_blockx_27_data_out), .map_block(_seach_blockx_27_map_block), .now(_seach_blockx_27_now));
seach_block seach_blockx_26 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_26_in_do), .start(_seach_blockx_26_start), .goal(_seach_blockx_26_goal), .data_out(_seach_blockx_26_data_out), .map_block(_seach_blockx_26_map_block), .now(_seach_blockx_26_now));
seach_block seach_blockx_25 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_25_in_do), .start(_seach_blockx_25_start), .goal(_seach_blockx_25_goal), .data_out(_seach_blockx_25_data_out), .map_block(_seach_blockx_25_map_block), .now(_seach_blockx_25_now));
seach_block seach_blockx_24 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_24_in_do), .start(_seach_blockx_24_start), .goal(_seach_blockx_24_goal), .data_out(_seach_blockx_24_data_out), .map_block(_seach_blockx_24_map_block), .now(_seach_blockx_24_now));
seach_block seach_blockx_23 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_23_in_do), .start(_seach_blockx_23_start), .goal(_seach_blockx_23_goal), .data_out(_seach_blockx_23_data_out), .map_block(_seach_blockx_23_map_block), .now(_seach_blockx_23_now));
seach_block seach_blockx_22 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_22_in_do), .start(_seach_blockx_22_start), .goal(_seach_blockx_22_goal), .data_out(_seach_blockx_22_data_out), .map_block(_seach_blockx_22_map_block), .now(_seach_blockx_22_now));
seach_block seach_blockx_21 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_21_in_do), .start(_seach_blockx_21_start), .goal(_seach_blockx_21_goal), .data_out(_seach_blockx_21_data_out), .map_block(_seach_blockx_21_map_block), .now(_seach_blockx_21_now));
seach_block seach_blockx_20 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_20_in_do), .start(_seach_blockx_20_start), .goal(_seach_blockx_20_goal), .data_out(_seach_blockx_20_data_out), .map_block(_seach_blockx_20_map_block), .now(_seach_blockx_20_now));
seach_block seach_blockx_19 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_19_in_do), .start(_seach_blockx_19_start), .goal(_seach_blockx_19_goal), .data_out(_seach_blockx_19_data_out), .map_block(_seach_blockx_19_map_block), .now(_seach_blockx_19_now));
seach_block seach_blockx_18 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_18_in_do), .start(_seach_blockx_18_start), .goal(_seach_blockx_18_goal), .data_out(_seach_blockx_18_data_out), .map_block(_seach_blockx_18_map_block), .now(_seach_blockx_18_now));
seach_block seach_blockx_17 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_17_in_do), .start(_seach_blockx_17_start), .goal(_seach_blockx_17_goal), .data_out(_seach_blockx_17_data_out), .map_block(_seach_blockx_17_map_block), .now(_seach_blockx_17_now));
seach_block seach_blockx_16 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_16_in_do), .start(_seach_blockx_16_start), .goal(_seach_blockx_16_goal), .data_out(_seach_blockx_16_data_out), .map_block(_seach_blockx_16_map_block), .now(_seach_blockx_16_now));
seach_block seach_blockx_15 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_15_in_do), .start(_seach_blockx_15_start), .goal(_seach_blockx_15_goal), .data_out(_seach_blockx_15_data_out), .map_block(_seach_blockx_15_map_block), .now(_seach_blockx_15_now));
seach_block seach_blockx_14 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_14_in_do), .start(_seach_blockx_14_start), .goal(_seach_blockx_14_goal), .data_out(_seach_blockx_14_data_out), .map_block(_seach_blockx_14_map_block), .now(_seach_blockx_14_now));
seach_block seach_blockx_13 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_13_in_do), .start(_seach_blockx_13_start), .goal(_seach_blockx_13_goal), .data_out(_seach_blockx_13_data_out), .map_block(_seach_blockx_13_map_block), .now(_seach_blockx_13_now));
seach_block seach_blockx_12 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_12_in_do), .start(_seach_blockx_12_start), .goal(_seach_blockx_12_goal), .data_out(_seach_blockx_12_data_out), .map_block(_seach_blockx_12_map_block), .now(_seach_blockx_12_now));
seach_block seach_blockx_11 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_11_in_do), .start(_seach_blockx_11_start), .goal(_seach_blockx_11_goal), .data_out(_seach_blockx_11_data_out), .map_block(_seach_blockx_11_map_block), .now(_seach_blockx_11_now));
seach_block seach_blockx_10 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_10_in_do), .start(_seach_blockx_10_start), .goal(_seach_blockx_10_goal), .data_out(_seach_blockx_10_data_out), .map_block(_seach_blockx_10_map_block), .now(_seach_blockx_10_now));
seach_block seach_blockx_9 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_9_in_do), .start(_seach_blockx_9_start), .goal(_seach_blockx_9_goal), .data_out(_seach_blockx_9_data_out), .map_block(_seach_blockx_9_map_block), .now(_seach_blockx_9_now));
seach_block seach_blockx_8 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_8_in_do), .start(_seach_blockx_8_start), .goal(_seach_blockx_8_goal), .data_out(_seach_blockx_8_data_out), .map_block(_seach_blockx_8_map_block), .now(_seach_blockx_8_now));
seach_block seach_blockx_7 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_7_in_do), .start(_seach_blockx_7_start), .goal(_seach_blockx_7_goal), .data_out(_seach_blockx_7_data_out), .map_block(_seach_blockx_7_map_block), .now(_seach_blockx_7_now));
seach_block seach_blockx_6 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_6_in_do), .start(_seach_blockx_6_start), .goal(_seach_blockx_6_goal), .data_out(_seach_blockx_6_data_out), .map_block(_seach_blockx_6_map_block), .now(_seach_blockx_6_now));
seach_block seach_blockx_5 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_5_in_do), .start(_seach_blockx_5_start), .goal(_seach_blockx_5_goal), .data_out(_seach_blockx_5_data_out), .map_block(_seach_blockx_5_map_block), .now(_seach_blockx_5_now));
seach_block seach_blockx_4 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_4_in_do), .start(_seach_blockx_4_start), .goal(_seach_blockx_4_goal), .data_out(_seach_blockx_4_data_out), .map_block(_seach_blockx_4_map_block), .now(_seach_blockx_4_now));
seach_block seach_blockx_3 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_3_in_do), .start(_seach_blockx_3_start), .goal(_seach_blockx_3_goal), .data_out(_seach_blockx_3_data_out), .map_block(_seach_blockx_3_map_block), .now(_seach_blockx_3_now));
seach_block seach_blockx_2 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_2_in_do), .start(_seach_blockx_2_start), .goal(_seach_blockx_2_goal), .data_out(_seach_blockx_2_data_out), .map_block(_seach_blockx_2_map_block), .now(_seach_blockx_2_now));
seach_block seach_blockx_1 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_1_in_do), .start(_seach_blockx_1_start), .goal(_seach_blockx_1_goal), .data_out(_seach_blockx_1_data_out), .map_block(_seach_blockx_1_map_block), .now(_seach_blockx_1_now));

   assign  _seach_blockx_map_block = data_in33;
   assign  _seach_blockx_now = 10'b0000100001;
   assign  _seach_blockx_in_do = _net_2;
   assign  _seach_blockx_p_reset = p_reset;
   assign  _seach_blockx_m_clock = m_clock;
   assign  _seach_blockx_419_map_block = data_in478;
   assign  _seach_blockx_419_now = 10'b0111011110;
   assign  _seach_blockx_419_in_do = _net_1259;
   assign  _seach_blockx_419_p_reset = p_reset;
   assign  _seach_blockx_419_m_clock = m_clock;
   assign  _seach_blockx_418_map_block = data_in477;
   assign  _seach_blockx_418_now = 10'b0111011101;
   assign  _seach_blockx_418_in_do = _net_1256;
   assign  _seach_blockx_418_p_reset = p_reset;
   assign  _seach_blockx_418_m_clock = m_clock;
   assign  _seach_blockx_417_map_block = data_in476;
   assign  _seach_blockx_417_now = 10'b0111011100;
   assign  _seach_blockx_417_in_do = _net_1253;
   assign  _seach_blockx_417_p_reset = p_reset;
   assign  _seach_blockx_417_m_clock = m_clock;
   assign  _seach_blockx_416_map_block = data_in475;
   assign  _seach_blockx_416_now = 10'b0111011011;
   assign  _seach_blockx_416_in_do = _net_1250;
   assign  _seach_blockx_416_p_reset = p_reset;
   assign  _seach_blockx_416_m_clock = m_clock;
   assign  _seach_blockx_415_map_block = data_in474;
   assign  _seach_blockx_415_now = 10'b0111011010;
   assign  _seach_blockx_415_in_do = _net_1247;
   assign  _seach_blockx_415_p_reset = p_reset;
   assign  _seach_blockx_415_m_clock = m_clock;
   assign  _seach_blockx_414_map_block = data_in473;
   assign  _seach_blockx_414_now = 10'b0111011001;
   assign  _seach_blockx_414_in_do = _net_1244;
   assign  _seach_blockx_414_p_reset = p_reset;
   assign  _seach_blockx_414_m_clock = m_clock;
   assign  _seach_blockx_413_map_block = data_in472;
   assign  _seach_blockx_413_now = 10'b0111011000;
   assign  _seach_blockx_413_in_do = _net_1241;
   assign  _seach_blockx_413_p_reset = p_reset;
   assign  _seach_blockx_413_m_clock = m_clock;
   assign  _seach_blockx_412_map_block = data_in471;
   assign  _seach_blockx_412_now = 10'b0111010111;
   assign  _seach_blockx_412_in_do = _net_1238;
   assign  _seach_blockx_412_p_reset = p_reset;
   assign  _seach_blockx_412_m_clock = m_clock;
   assign  _seach_blockx_411_map_block = data_in470;
   assign  _seach_blockx_411_now = 10'b0111010110;
   assign  _seach_blockx_411_in_do = _net_1235;
   assign  _seach_blockx_411_p_reset = p_reset;
   assign  _seach_blockx_411_m_clock = m_clock;
   assign  _seach_blockx_410_map_block = data_in469;
   assign  _seach_blockx_410_now = 10'b0111010101;
   assign  _seach_blockx_410_in_do = _net_1232;
   assign  _seach_blockx_410_p_reset = p_reset;
   assign  _seach_blockx_410_m_clock = m_clock;
   assign  _seach_blockx_409_map_block = data_in468;
   assign  _seach_blockx_409_now = 10'b0111010100;
   assign  _seach_blockx_409_in_do = _net_1229;
   assign  _seach_blockx_409_p_reset = p_reset;
   assign  _seach_blockx_409_m_clock = m_clock;
   assign  _seach_blockx_408_map_block = data_in467;
   assign  _seach_blockx_408_now = 10'b0111010011;
   assign  _seach_blockx_408_in_do = _net_1226;
   assign  _seach_blockx_408_p_reset = p_reset;
   assign  _seach_blockx_408_m_clock = m_clock;
   assign  _seach_blockx_407_map_block = data_in466;
   assign  _seach_blockx_407_now = 10'b0111010010;
   assign  _seach_blockx_407_in_do = _net_1223;
   assign  _seach_blockx_407_p_reset = p_reset;
   assign  _seach_blockx_407_m_clock = m_clock;
   assign  _seach_blockx_406_map_block = data_in465;
   assign  _seach_blockx_406_now = 10'b0111010001;
   assign  _seach_blockx_406_in_do = _net_1220;
   assign  _seach_blockx_406_p_reset = p_reset;
   assign  _seach_blockx_406_m_clock = m_clock;
   assign  _seach_blockx_405_map_block = data_in464;
   assign  _seach_blockx_405_now = 10'b0111010000;
   assign  _seach_blockx_405_in_do = _net_1217;
   assign  _seach_blockx_405_p_reset = p_reset;
   assign  _seach_blockx_405_m_clock = m_clock;
   assign  _seach_blockx_404_map_block = data_in463;
   assign  _seach_blockx_404_now = 10'b0111001111;
   assign  _seach_blockx_404_in_do = _net_1214;
   assign  _seach_blockx_404_p_reset = p_reset;
   assign  _seach_blockx_404_m_clock = m_clock;
   assign  _seach_blockx_403_map_block = data_in462;
   assign  _seach_blockx_403_now = 10'b0111001110;
   assign  _seach_blockx_403_in_do = _net_1211;
   assign  _seach_blockx_403_p_reset = p_reset;
   assign  _seach_blockx_403_m_clock = m_clock;
   assign  _seach_blockx_402_map_block = data_in461;
   assign  _seach_blockx_402_now = 10'b0111001101;
   assign  _seach_blockx_402_in_do = _net_1208;
   assign  _seach_blockx_402_p_reset = p_reset;
   assign  _seach_blockx_402_m_clock = m_clock;
   assign  _seach_blockx_401_map_block = data_in460;
   assign  _seach_blockx_401_now = 10'b0111001100;
   assign  _seach_blockx_401_in_do = _net_1205;
   assign  _seach_blockx_401_p_reset = p_reset;
   assign  _seach_blockx_401_m_clock = m_clock;
   assign  _seach_blockx_400_map_block = data_in459;
   assign  _seach_blockx_400_now = 10'b0111001011;
   assign  _seach_blockx_400_in_do = _net_1202;
   assign  _seach_blockx_400_p_reset = p_reset;
   assign  _seach_blockx_400_m_clock = m_clock;
   assign  _seach_blockx_399_map_block = data_in458;
   assign  _seach_blockx_399_now = 10'b0111001010;
   assign  _seach_blockx_399_in_do = _net_1199;
   assign  _seach_blockx_399_p_reset = p_reset;
   assign  _seach_blockx_399_m_clock = m_clock;
   assign  _seach_blockx_398_map_block = data_in457;
   assign  _seach_blockx_398_now = 10'b0111001001;
   assign  _seach_blockx_398_in_do = _net_1196;
   assign  _seach_blockx_398_p_reset = p_reset;
   assign  _seach_blockx_398_m_clock = m_clock;
   assign  _seach_blockx_397_map_block = data_in456;
   assign  _seach_blockx_397_now = 10'b0111001000;
   assign  _seach_blockx_397_in_do = _net_1193;
   assign  _seach_blockx_397_p_reset = p_reset;
   assign  _seach_blockx_397_m_clock = m_clock;
   assign  _seach_blockx_396_map_block = data_in455;
   assign  _seach_blockx_396_now = 10'b0111000111;
   assign  _seach_blockx_396_in_do = _net_1190;
   assign  _seach_blockx_396_p_reset = p_reset;
   assign  _seach_blockx_396_m_clock = m_clock;
   assign  _seach_blockx_395_map_block = data_in454;
   assign  _seach_blockx_395_now = 10'b0111000110;
   assign  _seach_blockx_395_in_do = _net_1187;
   assign  _seach_blockx_395_p_reset = p_reset;
   assign  _seach_blockx_395_m_clock = m_clock;
   assign  _seach_blockx_394_map_block = data_in453;
   assign  _seach_blockx_394_now = 10'b0111000101;
   assign  _seach_blockx_394_in_do = _net_1184;
   assign  _seach_blockx_394_p_reset = p_reset;
   assign  _seach_blockx_394_m_clock = m_clock;
   assign  _seach_blockx_393_map_block = data_in452;
   assign  _seach_blockx_393_now = 10'b0111000100;
   assign  _seach_blockx_393_in_do = _net_1181;
   assign  _seach_blockx_393_p_reset = p_reset;
   assign  _seach_blockx_393_m_clock = m_clock;
   assign  _seach_blockx_392_map_block = data_in451;
   assign  _seach_blockx_392_now = 10'b0111000011;
   assign  _seach_blockx_392_in_do = _net_1178;
   assign  _seach_blockx_392_p_reset = p_reset;
   assign  _seach_blockx_392_m_clock = m_clock;
   assign  _seach_blockx_391_map_block = data_in450;
   assign  _seach_blockx_391_now = 10'b0111000010;
   assign  _seach_blockx_391_in_do = _net_1175;
   assign  _seach_blockx_391_p_reset = p_reset;
   assign  _seach_blockx_391_m_clock = m_clock;
   assign  _seach_blockx_390_map_block = data_in449;
   assign  _seach_blockx_390_now = 10'b0111000001;
   assign  _seach_blockx_390_in_do = _net_1172;
   assign  _seach_blockx_390_p_reset = p_reset;
   assign  _seach_blockx_390_m_clock = m_clock;
   assign  _seach_blockx_389_map_block = data_in446;
   assign  _seach_blockx_389_now = 10'b0110111110;
   assign  _seach_blockx_389_in_do = _net_1169;
   assign  _seach_blockx_389_p_reset = p_reset;
   assign  _seach_blockx_389_m_clock = m_clock;
   assign  _seach_blockx_388_map_block = data_in445;
   assign  _seach_blockx_388_now = 10'b0110111101;
   assign  _seach_blockx_388_in_do = _net_1166;
   assign  _seach_blockx_388_p_reset = p_reset;
   assign  _seach_blockx_388_m_clock = m_clock;
   assign  _seach_blockx_387_map_block = data_in444;
   assign  _seach_blockx_387_now = 10'b0110111100;
   assign  _seach_blockx_387_in_do = _net_1163;
   assign  _seach_blockx_387_p_reset = p_reset;
   assign  _seach_blockx_387_m_clock = m_clock;
   assign  _seach_blockx_386_map_block = data_in443;
   assign  _seach_blockx_386_now = 10'b0110111011;
   assign  _seach_blockx_386_in_do = _net_1160;
   assign  _seach_blockx_386_p_reset = p_reset;
   assign  _seach_blockx_386_m_clock = m_clock;
   assign  _seach_blockx_385_map_block = data_in442;
   assign  _seach_blockx_385_now = 10'b0110111010;
   assign  _seach_blockx_385_in_do = _net_1157;
   assign  _seach_blockx_385_p_reset = p_reset;
   assign  _seach_blockx_385_m_clock = m_clock;
   assign  _seach_blockx_384_map_block = data_in441;
   assign  _seach_blockx_384_now = 10'b0110111001;
   assign  _seach_blockx_384_in_do = _net_1154;
   assign  _seach_blockx_384_p_reset = p_reset;
   assign  _seach_blockx_384_m_clock = m_clock;
   assign  _seach_blockx_383_map_block = data_in440;
   assign  _seach_blockx_383_now = 10'b0110111000;
   assign  _seach_blockx_383_in_do = _net_1151;
   assign  _seach_blockx_383_p_reset = p_reset;
   assign  _seach_blockx_383_m_clock = m_clock;
   assign  _seach_blockx_382_map_block = data_in439;
   assign  _seach_blockx_382_now = 10'b0110110111;
   assign  _seach_blockx_382_in_do = _net_1148;
   assign  _seach_blockx_382_p_reset = p_reset;
   assign  _seach_blockx_382_m_clock = m_clock;
   assign  _seach_blockx_381_map_block = data_in438;
   assign  _seach_blockx_381_now = 10'b0110110110;
   assign  _seach_blockx_381_in_do = _net_1145;
   assign  _seach_blockx_381_p_reset = p_reset;
   assign  _seach_blockx_381_m_clock = m_clock;
   assign  _seach_blockx_380_map_block = data_in437;
   assign  _seach_blockx_380_now = 10'b0110110101;
   assign  _seach_blockx_380_in_do = _net_1142;
   assign  _seach_blockx_380_p_reset = p_reset;
   assign  _seach_blockx_380_m_clock = m_clock;
   assign  _seach_blockx_379_map_block = data_in436;
   assign  _seach_blockx_379_now = 10'b0110110100;
   assign  _seach_blockx_379_in_do = _net_1139;
   assign  _seach_blockx_379_p_reset = p_reset;
   assign  _seach_blockx_379_m_clock = m_clock;
   assign  _seach_blockx_378_map_block = data_in435;
   assign  _seach_blockx_378_now = 10'b0110110011;
   assign  _seach_blockx_378_in_do = _net_1136;
   assign  _seach_blockx_378_p_reset = p_reset;
   assign  _seach_blockx_378_m_clock = m_clock;
   assign  _seach_blockx_377_map_block = data_in434;
   assign  _seach_blockx_377_now = 10'b0110110010;
   assign  _seach_blockx_377_in_do = _net_1133;
   assign  _seach_blockx_377_p_reset = p_reset;
   assign  _seach_blockx_377_m_clock = m_clock;
   assign  _seach_blockx_376_map_block = data_in433;
   assign  _seach_blockx_376_now = 10'b0110110001;
   assign  _seach_blockx_376_in_do = _net_1130;
   assign  _seach_blockx_376_p_reset = p_reset;
   assign  _seach_blockx_376_m_clock = m_clock;
   assign  _seach_blockx_375_map_block = data_in432;
   assign  _seach_blockx_375_now = 10'b0110110000;
   assign  _seach_blockx_375_in_do = _net_1127;
   assign  _seach_blockx_375_p_reset = p_reset;
   assign  _seach_blockx_375_m_clock = m_clock;
   assign  _seach_blockx_374_map_block = data_in431;
   assign  _seach_blockx_374_now = 10'b0110101111;
   assign  _seach_blockx_374_in_do = _net_1124;
   assign  _seach_blockx_374_p_reset = p_reset;
   assign  _seach_blockx_374_m_clock = m_clock;
   assign  _seach_blockx_373_map_block = data_in430;
   assign  _seach_blockx_373_now = 10'b0110101110;
   assign  _seach_blockx_373_in_do = _net_1121;
   assign  _seach_blockx_373_p_reset = p_reset;
   assign  _seach_blockx_373_m_clock = m_clock;
   assign  _seach_blockx_372_map_block = data_in429;
   assign  _seach_blockx_372_now = 10'b0110101101;
   assign  _seach_blockx_372_in_do = _net_1118;
   assign  _seach_blockx_372_p_reset = p_reset;
   assign  _seach_blockx_372_m_clock = m_clock;
   assign  _seach_blockx_371_map_block = data_in428;
   assign  _seach_blockx_371_now = 10'b0110101100;
   assign  _seach_blockx_371_in_do = _net_1115;
   assign  _seach_blockx_371_p_reset = p_reset;
   assign  _seach_blockx_371_m_clock = m_clock;
   assign  _seach_blockx_370_map_block = data_in427;
   assign  _seach_blockx_370_now = 10'b0110101011;
   assign  _seach_blockx_370_in_do = _net_1112;
   assign  _seach_blockx_370_p_reset = p_reset;
   assign  _seach_blockx_370_m_clock = m_clock;
   assign  _seach_blockx_369_map_block = data_in426;
   assign  _seach_blockx_369_now = 10'b0110101010;
   assign  _seach_blockx_369_in_do = _net_1109;
   assign  _seach_blockx_369_p_reset = p_reset;
   assign  _seach_blockx_369_m_clock = m_clock;
   assign  _seach_blockx_368_map_block = data_in425;
   assign  _seach_blockx_368_now = 10'b0110101001;
   assign  _seach_blockx_368_in_do = _net_1106;
   assign  _seach_blockx_368_p_reset = p_reset;
   assign  _seach_blockx_368_m_clock = m_clock;
   assign  _seach_blockx_367_map_block = data_in424;
   assign  _seach_blockx_367_now = 10'b0110101000;
   assign  _seach_blockx_367_in_do = _net_1103;
   assign  _seach_blockx_367_p_reset = p_reset;
   assign  _seach_blockx_367_m_clock = m_clock;
   assign  _seach_blockx_366_map_block = data_in423;
   assign  _seach_blockx_366_now = 10'b0110100111;
   assign  _seach_blockx_366_in_do = _net_1100;
   assign  _seach_blockx_366_p_reset = p_reset;
   assign  _seach_blockx_366_m_clock = m_clock;
   assign  _seach_blockx_365_map_block = data_in422;
   assign  _seach_blockx_365_now = 10'b0110100110;
   assign  _seach_blockx_365_in_do = _net_1097;
   assign  _seach_blockx_365_p_reset = p_reset;
   assign  _seach_blockx_365_m_clock = m_clock;
   assign  _seach_blockx_364_map_block = data_in421;
   assign  _seach_blockx_364_now = 10'b0110100101;
   assign  _seach_blockx_364_in_do = _net_1094;
   assign  _seach_blockx_364_p_reset = p_reset;
   assign  _seach_blockx_364_m_clock = m_clock;
   assign  _seach_blockx_363_map_block = data_in420;
   assign  _seach_blockx_363_now = 10'b0110100100;
   assign  _seach_blockx_363_in_do = _net_1091;
   assign  _seach_blockx_363_p_reset = p_reset;
   assign  _seach_blockx_363_m_clock = m_clock;
   assign  _seach_blockx_362_map_block = data_in419;
   assign  _seach_blockx_362_now = 10'b0110100011;
   assign  _seach_blockx_362_in_do = _net_1088;
   assign  _seach_blockx_362_p_reset = p_reset;
   assign  _seach_blockx_362_m_clock = m_clock;
   assign  _seach_blockx_361_map_block = data_in418;
   assign  _seach_blockx_361_now = 10'b0110100010;
   assign  _seach_blockx_361_in_do = _net_1085;
   assign  _seach_blockx_361_p_reset = p_reset;
   assign  _seach_blockx_361_m_clock = m_clock;
   assign  _seach_blockx_360_map_block = data_in417;
   assign  _seach_blockx_360_now = 10'b0110100001;
   assign  _seach_blockx_360_in_do = _net_1082;
   assign  _seach_blockx_360_p_reset = p_reset;
   assign  _seach_blockx_360_m_clock = m_clock;
   assign  _seach_blockx_359_map_block = data_in414;
   assign  _seach_blockx_359_now = 10'b0110011110;
   assign  _seach_blockx_359_in_do = _net_1079;
   assign  _seach_blockx_359_p_reset = p_reset;
   assign  _seach_blockx_359_m_clock = m_clock;
   assign  _seach_blockx_358_map_block = data_in413;
   assign  _seach_blockx_358_now = 10'b0110011101;
   assign  _seach_blockx_358_in_do = _net_1076;
   assign  _seach_blockx_358_p_reset = p_reset;
   assign  _seach_blockx_358_m_clock = m_clock;
   assign  _seach_blockx_357_map_block = data_in412;
   assign  _seach_blockx_357_now = 10'b0110011100;
   assign  _seach_blockx_357_in_do = _net_1073;
   assign  _seach_blockx_357_p_reset = p_reset;
   assign  _seach_blockx_357_m_clock = m_clock;
   assign  _seach_blockx_356_map_block = data_in411;
   assign  _seach_blockx_356_now = 10'b0110011011;
   assign  _seach_blockx_356_in_do = _net_1070;
   assign  _seach_blockx_356_p_reset = p_reset;
   assign  _seach_blockx_356_m_clock = m_clock;
   assign  _seach_blockx_355_map_block = data_in410;
   assign  _seach_blockx_355_now = 10'b0110011010;
   assign  _seach_blockx_355_in_do = _net_1067;
   assign  _seach_blockx_355_p_reset = p_reset;
   assign  _seach_blockx_355_m_clock = m_clock;
   assign  _seach_blockx_354_map_block = data_in409;
   assign  _seach_blockx_354_now = 10'b0110011001;
   assign  _seach_blockx_354_in_do = _net_1064;
   assign  _seach_blockx_354_p_reset = p_reset;
   assign  _seach_blockx_354_m_clock = m_clock;
   assign  _seach_blockx_353_map_block = data_in408;
   assign  _seach_blockx_353_now = 10'b0110011000;
   assign  _seach_blockx_353_in_do = _net_1061;
   assign  _seach_blockx_353_p_reset = p_reset;
   assign  _seach_blockx_353_m_clock = m_clock;
   assign  _seach_blockx_352_map_block = data_in407;
   assign  _seach_blockx_352_now = 10'b0110010111;
   assign  _seach_blockx_352_in_do = _net_1058;
   assign  _seach_blockx_352_p_reset = p_reset;
   assign  _seach_blockx_352_m_clock = m_clock;
   assign  _seach_blockx_351_map_block = data_in406;
   assign  _seach_blockx_351_now = 10'b0110010110;
   assign  _seach_blockx_351_in_do = _net_1055;
   assign  _seach_blockx_351_p_reset = p_reset;
   assign  _seach_blockx_351_m_clock = m_clock;
   assign  _seach_blockx_350_map_block = data_in405;
   assign  _seach_blockx_350_now = 10'b0110010101;
   assign  _seach_blockx_350_in_do = _net_1052;
   assign  _seach_blockx_350_p_reset = p_reset;
   assign  _seach_blockx_350_m_clock = m_clock;
   assign  _seach_blockx_349_map_block = data_in404;
   assign  _seach_blockx_349_now = 10'b0110010100;
   assign  _seach_blockx_349_in_do = _net_1049;
   assign  _seach_blockx_349_p_reset = p_reset;
   assign  _seach_blockx_349_m_clock = m_clock;
   assign  _seach_blockx_348_map_block = data_in403;
   assign  _seach_blockx_348_now = 10'b0110010011;
   assign  _seach_blockx_348_in_do = _net_1046;
   assign  _seach_blockx_348_p_reset = p_reset;
   assign  _seach_blockx_348_m_clock = m_clock;
   assign  _seach_blockx_347_map_block = data_in402;
   assign  _seach_blockx_347_now = 10'b0110010010;
   assign  _seach_blockx_347_in_do = _net_1043;
   assign  _seach_blockx_347_p_reset = p_reset;
   assign  _seach_blockx_347_m_clock = m_clock;
   assign  _seach_blockx_346_map_block = data_in401;
   assign  _seach_blockx_346_now = 10'b0110010001;
   assign  _seach_blockx_346_in_do = _net_1040;
   assign  _seach_blockx_346_p_reset = p_reset;
   assign  _seach_blockx_346_m_clock = m_clock;
   assign  _seach_blockx_345_map_block = data_in400;
   assign  _seach_blockx_345_now = 10'b0110010000;
   assign  _seach_blockx_345_in_do = _net_1037;
   assign  _seach_blockx_345_p_reset = p_reset;
   assign  _seach_blockx_345_m_clock = m_clock;
   assign  _seach_blockx_344_map_block = data_in399;
   assign  _seach_blockx_344_now = 10'b0110001111;
   assign  _seach_blockx_344_in_do = _net_1034;
   assign  _seach_blockx_344_p_reset = p_reset;
   assign  _seach_blockx_344_m_clock = m_clock;
   assign  _seach_blockx_343_map_block = data_in398;
   assign  _seach_blockx_343_now = 10'b0110001110;
   assign  _seach_blockx_343_in_do = _net_1031;
   assign  _seach_blockx_343_p_reset = p_reset;
   assign  _seach_blockx_343_m_clock = m_clock;
   assign  _seach_blockx_342_map_block = data_in397;
   assign  _seach_blockx_342_now = 10'b0110001101;
   assign  _seach_blockx_342_in_do = _net_1028;
   assign  _seach_blockx_342_p_reset = p_reset;
   assign  _seach_blockx_342_m_clock = m_clock;
   assign  _seach_blockx_341_map_block = data_in396;
   assign  _seach_blockx_341_now = 10'b0110001100;
   assign  _seach_blockx_341_in_do = _net_1025;
   assign  _seach_blockx_341_p_reset = p_reset;
   assign  _seach_blockx_341_m_clock = m_clock;
   assign  _seach_blockx_340_map_block = data_in395;
   assign  _seach_blockx_340_now = 10'b0110001011;
   assign  _seach_blockx_340_in_do = _net_1022;
   assign  _seach_blockx_340_p_reset = p_reset;
   assign  _seach_blockx_340_m_clock = m_clock;
   assign  _seach_blockx_339_map_block = data_in394;
   assign  _seach_blockx_339_now = 10'b0110001010;
   assign  _seach_blockx_339_in_do = _net_1019;
   assign  _seach_blockx_339_p_reset = p_reset;
   assign  _seach_blockx_339_m_clock = m_clock;
   assign  _seach_blockx_338_map_block = data_in393;
   assign  _seach_blockx_338_now = 10'b0110001001;
   assign  _seach_blockx_338_in_do = _net_1016;
   assign  _seach_blockx_338_p_reset = p_reset;
   assign  _seach_blockx_338_m_clock = m_clock;
   assign  _seach_blockx_337_map_block = data_in392;
   assign  _seach_blockx_337_now = 10'b0110001000;
   assign  _seach_blockx_337_in_do = _net_1013;
   assign  _seach_blockx_337_p_reset = p_reset;
   assign  _seach_blockx_337_m_clock = m_clock;
   assign  _seach_blockx_336_map_block = data_in391;
   assign  _seach_blockx_336_now = 10'b0110000111;
   assign  _seach_blockx_336_in_do = _net_1010;
   assign  _seach_blockx_336_p_reset = p_reset;
   assign  _seach_blockx_336_m_clock = m_clock;
   assign  _seach_blockx_335_map_block = data_in390;
   assign  _seach_blockx_335_now = 10'b0110000110;
   assign  _seach_blockx_335_in_do = _net_1007;
   assign  _seach_blockx_335_p_reset = p_reset;
   assign  _seach_blockx_335_m_clock = m_clock;
   assign  _seach_blockx_334_map_block = data_in389;
   assign  _seach_blockx_334_now = 10'b0110000101;
   assign  _seach_blockx_334_in_do = _net_1004;
   assign  _seach_blockx_334_p_reset = p_reset;
   assign  _seach_blockx_334_m_clock = m_clock;
   assign  _seach_blockx_333_map_block = data_in388;
   assign  _seach_blockx_333_now = 10'b0110000100;
   assign  _seach_blockx_333_in_do = _net_1001;
   assign  _seach_blockx_333_p_reset = p_reset;
   assign  _seach_blockx_333_m_clock = m_clock;
   assign  _seach_blockx_332_map_block = data_in387;
   assign  _seach_blockx_332_now = 10'b0110000011;
   assign  _seach_blockx_332_in_do = _net_998;
   assign  _seach_blockx_332_p_reset = p_reset;
   assign  _seach_blockx_332_m_clock = m_clock;
   assign  _seach_blockx_331_map_block = data_in386;
   assign  _seach_blockx_331_now = 10'b0110000010;
   assign  _seach_blockx_331_in_do = _net_995;
   assign  _seach_blockx_331_p_reset = p_reset;
   assign  _seach_blockx_331_m_clock = m_clock;
   assign  _seach_blockx_330_map_block = data_in385;
   assign  _seach_blockx_330_now = 10'b0110000001;
   assign  _seach_blockx_330_in_do = _net_992;
   assign  _seach_blockx_330_p_reset = p_reset;
   assign  _seach_blockx_330_m_clock = m_clock;
   assign  _seach_blockx_329_map_block = data_in382;
   assign  _seach_blockx_329_now = 10'b0101111110;
   assign  _seach_blockx_329_in_do = _net_989;
   assign  _seach_blockx_329_p_reset = p_reset;
   assign  _seach_blockx_329_m_clock = m_clock;
   assign  _seach_blockx_328_map_block = data_in381;
   assign  _seach_blockx_328_now = 10'b0101111101;
   assign  _seach_blockx_328_in_do = _net_986;
   assign  _seach_blockx_328_p_reset = p_reset;
   assign  _seach_blockx_328_m_clock = m_clock;
   assign  _seach_blockx_327_map_block = data_in380;
   assign  _seach_blockx_327_now = 10'b0101111100;
   assign  _seach_blockx_327_in_do = _net_983;
   assign  _seach_blockx_327_p_reset = p_reset;
   assign  _seach_blockx_327_m_clock = m_clock;
   assign  _seach_blockx_326_map_block = data_in379;
   assign  _seach_blockx_326_now = 10'b0101111011;
   assign  _seach_blockx_326_in_do = _net_980;
   assign  _seach_blockx_326_p_reset = p_reset;
   assign  _seach_blockx_326_m_clock = m_clock;
   assign  _seach_blockx_325_map_block = data_in378;
   assign  _seach_blockx_325_now = 10'b0101111010;
   assign  _seach_blockx_325_in_do = _net_977;
   assign  _seach_blockx_325_p_reset = p_reset;
   assign  _seach_blockx_325_m_clock = m_clock;
   assign  _seach_blockx_324_map_block = data_in377;
   assign  _seach_blockx_324_now = 10'b0101111001;
   assign  _seach_blockx_324_in_do = _net_974;
   assign  _seach_blockx_324_p_reset = p_reset;
   assign  _seach_blockx_324_m_clock = m_clock;
   assign  _seach_blockx_323_map_block = data_in376;
   assign  _seach_blockx_323_now = 10'b0101111000;
   assign  _seach_blockx_323_in_do = _net_971;
   assign  _seach_blockx_323_p_reset = p_reset;
   assign  _seach_blockx_323_m_clock = m_clock;
   assign  _seach_blockx_322_map_block = data_in375;
   assign  _seach_blockx_322_now = 10'b0101110111;
   assign  _seach_blockx_322_in_do = _net_968;
   assign  _seach_blockx_322_p_reset = p_reset;
   assign  _seach_blockx_322_m_clock = m_clock;
   assign  _seach_blockx_321_map_block = data_in374;
   assign  _seach_blockx_321_now = 10'b0101110110;
   assign  _seach_blockx_321_in_do = _net_965;
   assign  _seach_blockx_321_p_reset = p_reset;
   assign  _seach_blockx_321_m_clock = m_clock;
   assign  _seach_blockx_320_map_block = data_in373;
   assign  _seach_blockx_320_now = 10'b0101110101;
   assign  _seach_blockx_320_in_do = _net_962;
   assign  _seach_blockx_320_p_reset = p_reset;
   assign  _seach_blockx_320_m_clock = m_clock;
   assign  _seach_blockx_319_map_block = data_in372;
   assign  _seach_blockx_319_now = 10'b0101110100;
   assign  _seach_blockx_319_in_do = _net_959;
   assign  _seach_blockx_319_p_reset = p_reset;
   assign  _seach_blockx_319_m_clock = m_clock;
   assign  _seach_blockx_318_map_block = data_in371;
   assign  _seach_blockx_318_now = 10'b0101110011;
   assign  _seach_blockx_318_in_do = _net_956;
   assign  _seach_blockx_318_p_reset = p_reset;
   assign  _seach_blockx_318_m_clock = m_clock;
   assign  _seach_blockx_317_map_block = data_in370;
   assign  _seach_blockx_317_now = 10'b0101110010;
   assign  _seach_blockx_317_in_do = _net_953;
   assign  _seach_blockx_317_p_reset = p_reset;
   assign  _seach_blockx_317_m_clock = m_clock;
   assign  _seach_blockx_316_map_block = data_in369;
   assign  _seach_blockx_316_now = 10'b0101110001;
   assign  _seach_blockx_316_in_do = _net_950;
   assign  _seach_blockx_316_p_reset = p_reset;
   assign  _seach_blockx_316_m_clock = m_clock;
   assign  _seach_blockx_315_map_block = data_in368;
   assign  _seach_blockx_315_now = 10'b0101110000;
   assign  _seach_blockx_315_in_do = _net_947;
   assign  _seach_blockx_315_p_reset = p_reset;
   assign  _seach_blockx_315_m_clock = m_clock;
   assign  _seach_blockx_314_map_block = data_in367;
   assign  _seach_blockx_314_now = 10'b0101101111;
   assign  _seach_blockx_314_in_do = _net_944;
   assign  _seach_blockx_314_p_reset = p_reset;
   assign  _seach_blockx_314_m_clock = m_clock;
   assign  _seach_blockx_313_map_block = data_in366;
   assign  _seach_blockx_313_now = 10'b0101101110;
   assign  _seach_blockx_313_in_do = _net_941;
   assign  _seach_blockx_313_p_reset = p_reset;
   assign  _seach_blockx_313_m_clock = m_clock;
   assign  _seach_blockx_312_map_block = data_in365;
   assign  _seach_blockx_312_now = 10'b0101101101;
   assign  _seach_blockx_312_in_do = _net_938;
   assign  _seach_blockx_312_p_reset = p_reset;
   assign  _seach_blockx_312_m_clock = m_clock;
   assign  _seach_blockx_311_map_block = data_in364;
   assign  _seach_blockx_311_now = 10'b0101101100;
   assign  _seach_blockx_311_in_do = _net_935;
   assign  _seach_blockx_311_p_reset = p_reset;
   assign  _seach_blockx_311_m_clock = m_clock;
   assign  _seach_blockx_310_map_block = data_in363;
   assign  _seach_blockx_310_now = 10'b0101101011;
   assign  _seach_blockx_310_in_do = _net_932;
   assign  _seach_blockx_310_p_reset = p_reset;
   assign  _seach_blockx_310_m_clock = m_clock;
   assign  _seach_blockx_309_map_block = data_in362;
   assign  _seach_blockx_309_now = 10'b0101101010;
   assign  _seach_blockx_309_in_do = _net_929;
   assign  _seach_blockx_309_p_reset = p_reset;
   assign  _seach_blockx_309_m_clock = m_clock;
   assign  _seach_blockx_308_map_block = data_in361;
   assign  _seach_blockx_308_now = 10'b0101101001;
   assign  _seach_blockx_308_in_do = _net_926;
   assign  _seach_blockx_308_p_reset = p_reset;
   assign  _seach_blockx_308_m_clock = m_clock;
   assign  _seach_blockx_307_map_block = data_in360;
   assign  _seach_blockx_307_now = 10'b0101101000;
   assign  _seach_blockx_307_in_do = _net_923;
   assign  _seach_blockx_307_p_reset = p_reset;
   assign  _seach_blockx_307_m_clock = m_clock;
   assign  _seach_blockx_306_map_block = data_in359;
   assign  _seach_blockx_306_now = 10'b0101100111;
   assign  _seach_blockx_306_in_do = _net_920;
   assign  _seach_blockx_306_p_reset = p_reset;
   assign  _seach_blockx_306_m_clock = m_clock;
   assign  _seach_blockx_305_map_block = data_in358;
   assign  _seach_blockx_305_now = 10'b0101100110;
   assign  _seach_blockx_305_in_do = _net_917;
   assign  _seach_blockx_305_p_reset = p_reset;
   assign  _seach_blockx_305_m_clock = m_clock;
   assign  _seach_blockx_304_map_block = data_in357;
   assign  _seach_blockx_304_now = 10'b0101100101;
   assign  _seach_blockx_304_in_do = _net_914;
   assign  _seach_blockx_304_p_reset = p_reset;
   assign  _seach_blockx_304_m_clock = m_clock;
   assign  _seach_blockx_303_map_block = data_in356;
   assign  _seach_blockx_303_now = 10'b0101100100;
   assign  _seach_blockx_303_in_do = _net_911;
   assign  _seach_blockx_303_p_reset = p_reset;
   assign  _seach_blockx_303_m_clock = m_clock;
   assign  _seach_blockx_302_map_block = data_in355;
   assign  _seach_blockx_302_now = 10'b0101100011;
   assign  _seach_blockx_302_in_do = _net_908;
   assign  _seach_blockx_302_p_reset = p_reset;
   assign  _seach_blockx_302_m_clock = m_clock;
   assign  _seach_blockx_301_map_block = data_in354;
   assign  _seach_blockx_301_now = 10'b0101100010;
   assign  _seach_blockx_301_in_do = _net_905;
   assign  _seach_blockx_301_p_reset = p_reset;
   assign  _seach_blockx_301_m_clock = m_clock;
   assign  _seach_blockx_300_map_block = data_in353;
   assign  _seach_blockx_300_now = 10'b0101100001;
   assign  _seach_blockx_300_in_do = _net_902;
   assign  _seach_blockx_300_p_reset = p_reset;
   assign  _seach_blockx_300_m_clock = m_clock;
   assign  _seach_blockx_299_map_block = data_in350;
   assign  _seach_blockx_299_now = 10'b0101011110;
   assign  _seach_blockx_299_in_do = _net_899;
   assign  _seach_blockx_299_p_reset = p_reset;
   assign  _seach_blockx_299_m_clock = m_clock;
   assign  _seach_blockx_298_map_block = data_in349;
   assign  _seach_blockx_298_now = 10'b0101011101;
   assign  _seach_blockx_298_in_do = _net_896;
   assign  _seach_blockx_298_p_reset = p_reset;
   assign  _seach_blockx_298_m_clock = m_clock;
   assign  _seach_blockx_297_map_block = data_in348;
   assign  _seach_blockx_297_now = 10'b0101011100;
   assign  _seach_blockx_297_in_do = _net_893;
   assign  _seach_blockx_297_p_reset = p_reset;
   assign  _seach_blockx_297_m_clock = m_clock;
   assign  _seach_blockx_296_map_block = data_in347;
   assign  _seach_blockx_296_now = 10'b0101011011;
   assign  _seach_blockx_296_in_do = _net_890;
   assign  _seach_blockx_296_p_reset = p_reset;
   assign  _seach_blockx_296_m_clock = m_clock;
   assign  _seach_blockx_295_map_block = data_in346;
   assign  _seach_blockx_295_now = 10'b0101011010;
   assign  _seach_blockx_295_in_do = _net_887;
   assign  _seach_blockx_295_p_reset = p_reset;
   assign  _seach_blockx_295_m_clock = m_clock;
   assign  _seach_blockx_294_map_block = data_in345;
   assign  _seach_blockx_294_now = 10'b0101011001;
   assign  _seach_blockx_294_in_do = _net_884;
   assign  _seach_blockx_294_p_reset = p_reset;
   assign  _seach_blockx_294_m_clock = m_clock;
   assign  _seach_blockx_293_map_block = data_in344;
   assign  _seach_blockx_293_now = 10'b0101011000;
   assign  _seach_blockx_293_in_do = _net_881;
   assign  _seach_blockx_293_p_reset = p_reset;
   assign  _seach_blockx_293_m_clock = m_clock;
   assign  _seach_blockx_292_map_block = data_in343;
   assign  _seach_blockx_292_now = 10'b0101010111;
   assign  _seach_blockx_292_in_do = _net_878;
   assign  _seach_blockx_292_p_reset = p_reset;
   assign  _seach_blockx_292_m_clock = m_clock;
   assign  _seach_blockx_291_map_block = data_in342;
   assign  _seach_blockx_291_now = 10'b0101010110;
   assign  _seach_blockx_291_in_do = _net_875;
   assign  _seach_blockx_291_p_reset = p_reset;
   assign  _seach_blockx_291_m_clock = m_clock;
   assign  _seach_blockx_290_map_block = data_in341;
   assign  _seach_blockx_290_now = 10'b0101010101;
   assign  _seach_blockx_290_in_do = _net_872;
   assign  _seach_blockx_290_p_reset = p_reset;
   assign  _seach_blockx_290_m_clock = m_clock;
   assign  _seach_blockx_289_map_block = data_in340;
   assign  _seach_blockx_289_now = 10'b0101010100;
   assign  _seach_blockx_289_in_do = _net_869;
   assign  _seach_blockx_289_p_reset = p_reset;
   assign  _seach_blockx_289_m_clock = m_clock;
   assign  _seach_blockx_288_map_block = data_in339;
   assign  _seach_blockx_288_now = 10'b0101010011;
   assign  _seach_blockx_288_in_do = _net_866;
   assign  _seach_blockx_288_p_reset = p_reset;
   assign  _seach_blockx_288_m_clock = m_clock;
   assign  _seach_blockx_287_map_block = data_in338;
   assign  _seach_blockx_287_now = 10'b0101010010;
   assign  _seach_blockx_287_in_do = _net_863;
   assign  _seach_blockx_287_p_reset = p_reset;
   assign  _seach_blockx_287_m_clock = m_clock;
   assign  _seach_blockx_286_map_block = data_in337;
   assign  _seach_blockx_286_now = 10'b0101010001;
   assign  _seach_blockx_286_in_do = _net_860;
   assign  _seach_blockx_286_p_reset = p_reset;
   assign  _seach_blockx_286_m_clock = m_clock;
   assign  _seach_blockx_285_map_block = data_in336;
   assign  _seach_blockx_285_now = 10'b0101010000;
   assign  _seach_blockx_285_in_do = _net_857;
   assign  _seach_blockx_285_p_reset = p_reset;
   assign  _seach_blockx_285_m_clock = m_clock;
   assign  _seach_blockx_284_map_block = data_in335;
   assign  _seach_blockx_284_now = 10'b0101001111;
   assign  _seach_blockx_284_in_do = _net_854;
   assign  _seach_blockx_284_p_reset = p_reset;
   assign  _seach_blockx_284_m_clock = m_clock;
   assign  _seach_blockx_283_map_block = data_in334;
   assign  _seach_blockx_283_now = 10'b0101001110;
   assign  _seach_blockx_283_in_do = _net_851;
   assign  _seach_blockx_283_p_reset = p_reset;
   assign  _seach_blockx_283_m_clock = m_clock;
   assign  _seach_blockx_282_map_block = data_in333;
   assign  _seach_blockx_282_now = 10'b0101001101;
   assign  _seach_blockx_282_in_do = _net_848;
   assign  _seach_blockx_282_p_reset = p_reset;
   assign  _seach_blockx_282_m_clock = m_clock;
   assign  _seach_blockx_281_map_block = data_in332;
   assign  _seach_blockx_281_now = 10'b0101001100;
   assign  _seach_blockx_281_in_do = _net_845;
   assign  _seach_blockx_281_p_reset = p_reset;
   assign  _seach_blockx_281_m_clock = m_clock;
   assign  _seach_blockx_280_map_block = data_in331;
   assign  _seach_blockx_280_now = 10'b0101001011;
   assign  _seach_blockx_280_in_do = _net_842;
   assign  _seach_blockx_280_p_reset = p_reset;
   assign  _seach_blockx_280_m_clock = m_clock;
   assign  _seach_blockx_279_map_block = data_in330;
   assign  _seach_blockx_279_now = 10'b0101001010;
   assign  _seach_blockx_279_in_do = _net_839;
   assign  _seach_blockx_279_p_reset = p_reset;
   assign  _seach_blockx_279_m_clock = m_clock;
   assign  _seach_blockx_278_map_block = data_in329;
   assign  _seach_blockx_278_now = 10'b0101001001;
   assign  _seach_blockx_278_in_do = _net_836;
   assign  _seach_blockx_278_p_reset = p_reset;
   assign  _seach_blockx_278_m_clock = m_clock;
   assign  _seach_blockx_277_map_block = data_in328;
   assign  _seach_blockx_277_now = 10'b0101001000;
   assign  _seach_blockx_277_in_do = _net_833;
   assign  _seach_blockx_277_p_reset = p_reset;
   assign  _seach_blockx_277_m_clock = m_clock;
   assign  _seach_blockx_276_map_block = data_in327;
   assign  _seach_blockx_276_now = 10'b0101000111;
   assign  _seach_blockx_276_in_do = _net_830;
   assign  _seach_blockx_276_p_reset = p_reset;
   assign  _seach_blockx_276_m_clock = m_clock;
   assign  _seach_blockx_275_map_block = data_in326;
   assign  _seach_blockx_275_now = 10'b0101000110;
   assign  _seach_blockx_275_in_do = _net_827;
   assign  _seach_blockx_275_p_reset = p_reset;
   assign  _seach_blockx_275_m_clock = m_clock;
   assign  _seach_blockx_274_map_block = data_in325;
   assign  _seach_blockx_274_now = 10'b0101000101;
   assign  _seach_blockx_274_in_do = _net_824;
   assign  _seach_blockx_274_p_reset = p_reset;
   assign  _seach_blockx_274_m_clock = m_clock;
   assign  _seach_blockx_273_map_block = data_in324;
   assign  _seach_blockx_273_now = 10'b0101000100;
   assign  _seach_blockx_273_in_do = _net_821;
   assign  _seach_blockx_273_p_reset = p_reset;
   assign  _seach_blockx_273_m_clock = m_clock;
   assign  _seach_blockx_272_map_block = data_in323;
   assign  _seach_blockx_272_now = 10'b0101000011;
   assign  _seach_blockx_272_in_do = _net_818;
   assign  _seach_blockx_272_p_reset = p_reset;
   assign  _seach_blockx_272_m_clock = m_clock;
   assign  _seach_blockx_271_map_block = data_in322;
   assign  _seach_blockx_271_now = 10'b0101000010;
   assign  _seach_blockx_271_in_do = _net_815;
   assign  _seach_blockx_271_p_reset = p_reset;
   assign  _seach_blockx_271_m_clock = m_clock;
   assign  _seach_blockx_270_map_block = data_in321;
   assign  _seach_blockx_270_now = 10'b0101000001;
   assign  _seach_blockx_270_in_do = _net_812;
   assign  _seach_blockx_270_p_reset = p_reset;
   assign  _seach_blockx_270_m_clock = m_clock;
   assign  _seach_blockx_269_map_block = data_in318;
   assign  _seach_blockx_269_now = 10'b0100111110;
   assign  _seach_blockx_269_in_do = _net_809;
   assign  _seach_blockx_269_p_reset = p_reset;
   assign  _seach_blockx_269_m_clock = m_clock;
   assign  _seach_blockx_268_map_block = data_in317;
   assign  _seach_blockx_268_now = 10'b0100111101;
   assign  _seach_blockx_268_in_do = _net_806;
   assign  _seach_blockx_268_p_reset = p_reset;
   assign  _seach_blockx_268_m_clock = m_clock;
   assign  _seach_blockx_267_map_block = data_in316;
   assign  _seach_blockx_267_now = 10'b0100111100;
   assign  _seach_blockx_267_in_do = _net_803;
   assign  _seach_blockx_267_p_reset = p_reset;
   assign  _seach_blockx_267_m_clock = m_clock;
   assign  _seach_blockx_266_map_block = data_in315;
   assign  _seach_blockx_266_now = 10'b0100111011;
   assign  _seach_blockx_266_in_do = _net_800;
   assign  _seach_blockx_266_p_reset = p_reset;
   assign  _seach_blockx_266_m_clock = m_clock;
   assign  _seach_blockx_265_map_block = data_in314;
   assign  _seach_blockx_265_now = 10'b0100111010;
   assign  _seach_blockx_265_in_do = _net_797;
   assign  _seach_blockx_265_p_reset = p_reset;
   assign  _seach_blockx_265_m_clock = m_clock;
   assign  _seach_blockx_264_map_block = data_in313;
   assign  _seach_blockx_264_now = 10'b0100111001;
   assign  _seach_blockx_264_in_do = _net_794;
   assign  _seach_blockx_264_p_reset = p_reset;
   assign  _seach_blockx_264_m_clock = m_clock;
   assign  _seach_blockx_263_map_block = data_in312;
   assign  _seach_blockx_263_now = 10'b0100111000;
   assign  _seach_blockx_263_in_do = _net_791;
   assign  _seach_blockx_263_p_reset = p_reset;
   assign  _seach_blockx_263_m_clock = m_clock;
   assign  _seach_blockx_262_map_block = data_in311;
   assign  _seach_blockx_262_now = 10'b0100110111;
   assign  _seach_blockx_262_in_do = _net_788;
   assign  _seach_blockx_262_p_reset = p_reset;
   assign  _seach_blockx_262_m_clock = m_clock;
   assign  _seach_blockx_261_map_block = data_in310;
   assign  _seach_blockx_261_now = 10'b0100110110;
   assign  _seach_blockx_261_in_do = _net_785;
   assign  _seach_blockx_261_p_reset = p_reset;
   assign  _seach_blockx_261_m_clock = m_clock;
   assign  _seach_blockx_260_map_block = data_in309;
   assign  _seach_blockx_260_now = 10'b0100110101;
   assign  _seach_blockx_260_in_do = _net_782;
   assign  _seach_blockx_260_p_reset = p_reset;
   assign  _seach_blockx_260_m_clock = m_clock;
   assign  _seach_blockx_259_map_block = data_in308;
   assign  _seach_blockx_259_now = 10'b0100110100;
   assign  _seach_blockx_259_in_do = _net_779;
   assign  _seach_blockx_259_p_reset = p_reset;
   assign  _seach_blockx_259_m_clock = m_clock;
   assign  _seach_blockx_258_map_block = data_in307;
   assign  _seach_blockx_258_now = 10'b0100110011;
   assign  _seach_blockx_258_in_do = _net_776;
   assign  _seach_blockx_258_p_reset = p_reset;
   assign  _seach_blockx_258_m_clock = m_clock;
   assign  _seach_blockx_257_map_block = data_in306;
   assign  _seach_blockx_257_now = 10'b0100110010;
   assign  _seach_blockx_257_in_do = _net_773;
   assign  _seach_blockx_257_p_reset = p_reset;
   assign  _seach_blockx_257_m_clock = m_clock;
   assign  _seach_blockx_256_map_block = data_in305;
   assign  _seach_blockx_256_now = 10'b0100110001;
   assign  _seach_blockx_256_in_do = _net_770;
   assign  _seach_blockx_256_p_reset = p_reset;
   assign  _seach_blockx_256_m_clock = m_clock;
   assign  _seach_blockx_255_map_block = data_in304;
   assign  _seach_blockx_255_now = 10'b0100110000;
   assign  _seach_blockx_255_in_do = _net_767;
   assign  _seach_blockx_255_p_reset = p_reset;
   assign  _seach_blockx_255_m_clock = m_clock;
   assign  _seach_blockx_254_map_block = data_in303;
   assign  _seach_blockx_254_now = 10'b0100101111;
   assign  _seach_blockx_254_in_do = _net_764;
   assign  _seach_blockx_254_p_reset = p_reset;
   assign  _seach_blockx_254_m_clock = m_clock;
   assign  _seach_blockx_253_map_block = data_in302;
   assign  _seach_blockx_253_now = 10'b0100101110;
   assign  _seach_blockx_253_in_do = _net_761;
   assign  _seach_blockx_253_p_reset = p_reset;
   assign  _seach_blockx_253_m_clock = m_clock;
   assign  _seach_blockx_252_map_block = data_in301;
   assign  _seach_blockx_252_now = 10'b0100101101;
   assign  _seach_blockx_252_in_do = _net_758;
   assign  _seach_blockx_252_p_reset = p_reset;
   assign  _seach_blockx_252_m_clock = m_clock;
   assign  _seach_blockx_251_map_block = data_in300;
   assign  _seach_blockx_251_now = 10'b0100101100;
   assign  _seach_blockx_251_in_do = _net_755;
   assign  _seach_blockx_251_p_reset = p_reset;
   assign  _seach_blockx_251_m_clock = m_clock;
   assign  _seach_blockx_250_map_block = data_in299;
   assign  _seach_blockx_250_now = 10'b0100101011;
   assign  _seach_blockx_250_in_do = _net_752;
   assign  _seach_blockx_250_p_reset = p_reset;
   assign  _seach_blockx_250_m_clock = m_clock;
   assign  _seach_blockx_249_map_block = data_in298;
   assign  _seach_blockx_249_now = 10'b0100101010;
   assign  _seach_blockx_249_in_do = _net_749;
   assign  _seach_blockx_249_p_reset = p_reset;
   assign  _seach_blockx_249_m_clock = m_clock;
   assign  _seach_blockx_248_map_block = data_in297;
   assign  _seach_blockx_248_now = 10'b0100101001;
   assign  _seach_blockx_248_in_do = _net_746;
   assign  _seach_blockx_248_p_reset = p_reset;
   assign  _seach_blockx_248_m_clock = m_clock;
   assign  _seach_blockx_247_map_block = data_in296;
   assign  _seach_blockx_247_now = 10'b0100101000;
   assign  _seach_blockx_247_in_do = _net_743;
   assign  _seach_blockx_247_p_reset = p_reset;
   assign  _seach_blockx_247_m_clock = m_clock;
   assign  _seach_blockx_246_map_block = data_in295;
   assign  _seach_blockx_246_now = 10'b0100100111;
   assign  _seach_blockx_246_in_do = _net_740;
   assign  _seach_blockx_246_p_reset = p_reset;
   assign  _seach_blockx_246_m_clock = m_clock;
   assign  _seach_blockx_245_map_block = data_in294;
   assign  _seach_blockx_245_now = 10'b0100100110;
   assign  _seach_blockx_245_in_do = _net_737;
   assign  _seach_blockx_245_p_reset = p_reset;
   assign  _seach_blockx_245_m_clock = m_clock;
   assign  _seach_blockx_244_map_block = data_in293;
   assign  _seach_blockx_244_now = 10'b0100100101;
   assign  _seach_blockx_244_in_do = _net_734;
   assign  _seach_blockx_244_p_reset = p_reset;
   assign  _seach_blockx_244_m_clock = m_clock;
   assign  _seach_blockx_243_map_block = data_in292;
   assign  _seach_blockx_243_now = 10'b0100100100;
   assign  _seach_blockx_243_in_do = _net_731;
   assign  _seach_blockx_243_p_reset = p_reset;
   assign  _seach_blockx_243_m_clock = m_clock;
   assign  _seach_blockx_242_map_block = data_in291;
   assign  _seach_blockx_242_now = 10'b0100100011;
   assign  _seach_blockx_242_in_do = _net_728;
   assign  _seach_blockx_242_p_reset = p_reset;
   assign  _seach_blockx_242_m_clock = m_clock;
   assign  _seach_blockx_241_map_block = data_in290;
   assign  _seach_blockx_241_now = 10'b0100100010;
   assign  _seach_blockx_241_in_do = _net_725;
   assign  _seach_blockx_241_p_reset = p_reset;
   assign  _seach_blockx_241_m_clock = m_clock;
   assign  _seach_blockx_240_map_block = data_in289;
   assign  _seach_blockx_240_now = 10'b0100100001;
   assign  _seach_blockx_240_in_do = _net_722;
   assign  _seach_blockx_240_p_reset = p_reset;
   assign  _seach_blockx_240_m_clock = m_clock;
   assign  _seach_blockx_239_map_block = data_in286;
   assign  _seach_blockx_239_now = 10'b0100011110;
   assign  _seach_blockx_239_in_do = _net_719;
   assign  _seach_blockx_239_p_reset = p_reset;
   assign  _seach_blockx_239_m_clock = m_clock;
   assign  _seach_blockx_238_map_block = data_in285;
   assign  _seach_blockx_238_now = 10'b0100011101;
   assign  _seach_blockx_238_in_do = _net_716;
   assign  _seach_blockx_238_p_reset = p_reset;
   assign  _seach_blockx_238_m_clock = m_clock;
   assign  _seach_blockx_237_map_block = data_in284;
   assign  _seach_blockx_237_now = 10'b0100011100;
   assign  _seach_blockx_237_in_do = _net_713;
   assign  _seach_blockx_237_p_reset = p_reset;
   assign  _seach_blockx_237_m_clock = m_clock;
   assign  _seach_blockx_236_map_block = data_in283;
   assign  _seach_blockx_236_now = 10'b0100011011;
   assign  _seach_blockx_236_in_do = _net_710;
   assign  _seach_blockx_236_p_reset = p_reset;
   assign  _seach_blockx_236_m_clock = m_clock;
   assign  _seach_blockx_235_map_block = data_in282;
   assign  _seach_blockx_235_now = 10'b0100011010;
   assign  _seach_blockx_235_in_do = _net_707;
   assign  _seach_blockx_235_p_reset = p_reset;
   assign  _seach_blockx_235_m_clock = m_clock;
   assign  _seach_blockx_234_map_block = data_in281;
   assign  _seach_blockx_234_now = 10'b0100011001;
   assign  _seach_blockx_234_in_do = _net_704;
   assign  _seach_blockx_234_p_reset = p_reset;
   assign  _seach_blockx_234_m_clock = m_clock;
   assign  _seach_blockx_233_map_block = data_in280;
   assign  _seach_blockx_233_now = 10'b0100011000;
   assign  _seach_blockx_233_in_do = _net_701;
   assign  _seach_blockx_233_p_reset = p_reset;
   assign  _seach_blockx_233_m_clock = m_clock;
   assign  _seach_blockx_232_map_block = data_in279;
   assign  _seach_blockx_232_now = 10'b0100010111;
   assign  _seach_blockx_232_in_do = _net_698;
   assign  _seach_blockx_232_p_reset = p_reset;
   assign  _seach_blockx_232_m_clock = m_clock;
   assign  _seach_blockx_231_map_block = data_in278;
   assign  _seach_blockx_231_now = 10'b0100010110;
   assign  _seach_blockx_231_in_do = _net_695;
   assign  _seach_blockx_231_p_reset = p_reset;
   assign  _seach_blockx_231_m_clock = m_clock;
   assign  _seach_blockx_230_map_block = data_in277;
   assign  _seach_blockx_230_now = 10'b0100010101;
   assign  _seach_blockx_230_in_do = _net_692;
   assign  _seach_blockx_230_p_reset = p_reset;
   assign  _seach_blockx_230_m_clock = m_clock;
   assign  _seach_blockx_229_map_block = data_in276;
   assign  _seach_blockx_229_now = 10'b0100010100;
   assign  _seach_blockx_229_in_do = _net_689;
   assign  _seach_blockx_229_p_reset = p_reset;
   assign  _seach_blockx_229_m_clock = m_clock;
   assign  _seach_blockx_228_map_block = data_in275;
   assign  _seach_blockx_228_now = 10'b0100010011;
   assign  _seach_blockx_228_in_do = _net_686;
   assign  _seach_blockx_228_p_reset = p_reset;
   assign  _seach_blockx_228_m_clock = m_clock;
   assign  _seach_blockx_227_map_block = data_in274;
   assign  _seach_blockx_227_now = 10'b0100010010;
   assign  _seach_blockx_227_in_do = _net_683;
   assign  _seach_blockx_227_p_reset = p_reset;
   assign  _seach_blockx_227_m_clock = m_clock;
   assign  _seach_blockx_226_map_block = data_in273;
   assign  _seach_blockx_226_now = 10'b0100010001;
   assign  _seach_blockx_226_in_do = _net_680;
   assign  _seach_blockx_226_p_reset = p_reset;
   assign  _seach_blockx_226_m_clock = m_clock;
   assign  _seach_blockx_225_map_block = data_in272;
   assign  _seach_blockx_225_now = 10'b0100010000;
   assign  _seach_blockx_225_in_do = _net_677;
   assign  _seach_blockx_225_p_reset = p_reset;
   assign  _seach_blockx_225_m_clock = m_clock;
   assign  _seach_blockx_224_map_block = data_in271;
   assign  _seach_blockx_224_now = 10'b0100001111;
   assign  _seach_blockx_224_in_do = _net_674;
   assign  _seach_blockx_224_p_reset = p_reset;
   assign  _seach_blockx_224_m_clock = m_clock;
   assign  _seach_blockx_223_map_block = data_in270;
   assign  _seach_blockx_223_now = 10'b0100001110;
   assign  _seach_blockx_223_in_do = _net_671;
   assign  _seach_blockx_223_p_reset = p_reset;
   assign  _seach_blockx_223_m_clock = m_clock;
   assign  _seach_blockx_222_map_block = data_in269;
   assign  _seach_blockx_222_now = 10'b0100001101;
   assign  _seach_blockx_222_in_do = _net_668;
   assign  _seach_blockx_222_p_reset = p_reset;
   assign  _seach_blockx_222_m_clock = m_clock;
   assign  _seach_blockx_221_map_block = data_in268;
   assign  _seach_blockx_221_now = 10'b0100001100;
   assign  _seach_blockx_221_in_do = _net_665;
   assign  _seach_blockx_221_p_reset = p_reset;
   assign  _seach_blockx_221_m_clock = m_clock;
   assign  _seach_blockx_220_map_block = data_in267;
   assign  _seach_blockx_220_now = 10'b0100001011;
   assign  _seach_blockx_220_in_do = _net_662;
   assign  _seach_blockx_220_p_reset = p_reset;
   assign  _seach_blockx_220_m_clock = m_clock;
   assign  _seach_blockx_219_map_block = data_in266;
   assign  _seach_blockx_219_now = 10'b0100001010;
   assign  _seach_blockx_219_in_do = _net_659;
   assign  _seach_blockx_219_p_reset = p_reset;
   assign  _seach_blockx_219_m_clock = m_clock;
   assign  _seach_blockx_218_map_block = data_in265;
   assign  _seach_blockx_218_now = 10'b0100001001;
   assign  _seach_blockx_218_in_do = _net_656;
   assign  _seach_blockx_218_p_reset = p_reset;
   assign  _seach_blockx_218_m_clock = m_clock;
   assign  _seach_blockx_217_map_block = data_in264;
   assign  _seach_blockx_217_now = 10'b0100001000;
   assign  _seach_blockx_217_in_do = _net_653;
   assign  _seach_blockx_217_p_reset = p_reset;
   assign  _seach_blockx_217_m_clock = m_clock;
   assign  _seach_blockx_216_map_block = data_in263;
   assign  _seach_blockx_216_now = 10'b0100000111;
   assign  _seach_blockx_216_in_do = _net_650;
   assign  _seach_blockx_216_p_reset = p_reset;
   assign  _seach_blockx_216_m_clock = m_clock;
   assign  _seach_blockx_215_map_block = data_in262;
   assign  _seach_blockx_215_now = 10'b0100000110;
   assign  _seach_blockx_215_in_do = _net_647;
   assign  _seach_blockx_215_p_reset = p_reset;
   assign  _seach_blockx_215_m_clock = m_clock;
   assign  _seach_blockx_214_map_block = data_in261;
   assign  _seach_blockx_214_now = 10'b0100000101;
   assign  _seach_blockx_214_in_do = _net_644;
   assign  _seach_blockx_214_p_reset = p_reset;
   assign  _seach_blockx_214_m_clock = m_clock;
   assign  _seach_blockx_213_map_block = data_in260;
   assign  _seach_blockx_213_now = 10'b0100000100;
   assign  _seach_blockx_213_in_do = _net_641;
   assign  _seach_blockx_213_p_reset = p_reset;
   assign  _seach_blockx_213_m_clock = m_clock;
   assign  _seach_blockx_212_map_block = data_in259;
   assign  _seach_blockx_212_now = 10'b0100000011;
   assign  _seach_blockx_212_in_do = _net_638;
   assign  _seach_blockx_212_p_reset = p_reset;
   assign  _seach_blockx_212_m_clock = m_clock;
   assign  _seach_blockx_211_map_block = data_in258;
   assign  _seach_blockx_211_now = 10'b0100000010;
   assign  _seach_blockx_211_in_do = _net_635;
   assign  _seach_blockx_211_p_reset = p_reset;
   assign  _seach_blockx_211_m_clock = m_clock;
   assign  _seach_blockx_210_map_block = data_in257;
   assign  _seach_blockx_210_now = 10'b0100000001;
   assign  _seach_blockx_210_in_do = _net_632;
   assign  _seach_blockx_210_p_reset = p_reset;
   assign  _seach_blockx_210_m_clock = m_clock;
   assign  _seach_blockx_209_map_block = data_in254;
   assign  _seach_blockx_209_now = 10'b0011111110;
   assign  _seach_blockx_209_in_do = _net_629;
   assign  _seach_blockx_209_p_reset = p_reset;
   assign  _seach_blockx_209_m_clock = m_clock;
   assign  _seach_blockx_208_map_block = data_in253;
   assign  _seach_blockx_208_now = 10'b0011111101;
   assign  _seach_blockx_208_in_do = _net_626;
   assign  _seach_blockx_208_p_reset = p_reset;
   assign  _seach_blockx_208_m_clock = m_clock;
   assign  _seach_blockx_207_map_block = data_in252;
   assign  _seach_blockx_207_now = 10'b0011111100;
   assign  _seach_blockx_207_in_do = _net_623;
   assign  _seach_blockx_207_p_reset = p_reset;
   assign  _seach_blockx_207_m_clock = m_clock;
   assign  _seach_blockx_206_map_block = data_in251;
   assign  _seach_blockx_206_now = 10'b0011111011;
   assign  _seach_blockx_206_in_do = _net_620;
   assign  _seach_blockx_206_p_reset = p_reset;
   assign  _seach_blockx_206_m_clock = m_clock;
   assign  _seach_blockx_205_map_block = data_in250;
   assign  _seach_blockx_205_now = 10'b0011111010;
   assign  _seach_blockx_205_in_do = _net_617;
   assign  _seach_blockx_205_p_reset = p_reset;
   assign  _seach_blockx_205_m_clock = m_clock;
   assign  _seach_blockx_204_map_block = data_in249;
   assign  _seach_blockx_204_now = 10'b0011111001;
   assign  _seach_blockx_204_in_do = _net_614;
   assign  _seach_blockx_204_p_reset = p_reset;
   assign  _seach_blockx_204_m_clock = m_clock;
   assign  _seach_blockx_203_map_block = data_in248;
   assign  _seach_blockx_203_now = 10'b0011111000;
   assign  _seach_blockx_203_in_do = _net_611;
   assign  _seach_blockx_203_p_reset = p_reset;
   assign  _seach_blockx_203_m_clock = m_clock;
   assign  _seach_blockx_202_map_block = data_in247;
   assign  _seach_blockx_202_now = 10'b0011110111;
   assign  _seach_blockx_202_in_do = _net_608;
   assign  _seach_blockx_202_p_reset = p_reset;
   assign  _seach_blockx_202_m_clock = m_clock;
   assign  _seach_blockx_201_map_block = data_in246;
   assign  _seach_blockx_201_now = 10'b0011110110;
   assign  _seach_blockx_201_in_do = _net_605;
   assign  _seach_blockx_201_p_reset = p_reset;
   assign  _seach_blockx_201_m_clock = m_clock;
   assign  _seach_blockx_200_map_block = data_in245;
   assign  _seach_blockx_200_now = 10'b0011110101;
   assign  _seach_blockx_200_in_do = _net_602;
   assign  _seach_blockx_200_p_reset = p_reset;
   assign  _seach_blockx_200_m_clock = m_clock;
   assign  _seach_blockx_199_map_block = data_in244;
   assign  _seach_blockx_199_now = 10'b0011110100;
   assign  _seach_blockx_199_in_do = _net_599;
   assign  _seach_blockx_199_p_reset = p_reset;
   assign  _seach_blockx_199_m_clock = m_clock;
   assign  _seach_blockx_198_map_block = data_in243;
   assign  _seach_blockx_198_now = 10'b0011110011;
   assign  _seach_blockx_198_in_do = _net_596;
   assign  _seach_blockx_198_p_reset = p_reset;
   assign  _seach_blockx_198_m_clock = m_clock;
   assign  _seach_blockx_197_map_block = data_in242;
   assign  _seach_blockx_197_now = 10'b0011110010;
   assign  _seach_blockx_197_in_do = _net_593;
   assign  _seach_blockx_197_p_reset = p_reset;
   assign  _seach_blockx_197_m_clock = m_clock;
   assign  _seach_blockx_196_map_block = data_in241;
   assign  _seach_blockx_196_now = 10'b0011110001;
   assign  _seach_blockx_196_in_do = _net_590;
   assign  _seach_blockx_196_p_reset = p_reset;
   assign  _seach_blockx_196_m_clock = m_clock;
   assign  _seach_blockx_195_map_block = data_in240;
   assign  _seach_blockx_195_now = 10'b0011110000;
   assign  _seach_blockx_195_in_do = _net_587;
   assign  _seach_blockx_195_p_reset = p_reset;
   assign  _seach_blockx_195_m_clock = m_clock;
   assign  _seach_blockx_194_map_block = data_in239;
   assign  _seach_blockx_194_now = 10'b0011101111;
   assign  _seach_blockx_194_in_do = _net_584;
   assign  _seach_blockx_194_p_reset = p_reset;
   assign  _seach_blockx_194_m_clock = m_clock;
   assign  _seach_blockx_193_map_block = data_in238;
   assign  _seach_blockx_193_now = 10'b0011101110;
   assign  _seach_blockx_193_in_do = _net_581;
   assign  _seach_blockx_193_p_reset = p_reset;
   assign  _seach_blockx_193_m_clock = m_clock;
   assign  _seach_blockx_192_map_block = data_in237;
   assign  _seach_blockx_192_now = 10'b0011101101;
   assign  _seach_blockx_192_in_do = _net_578;
   assign  _seach_blockx_192_p_reset = p_reset;
   assign  _seach_blockx_192_m_clock = m_clock;
   assign  _seach_blockx_191_map_block = data_in236;
   assign  _seach_blockx_191_now = 10'b0011101100;
   assign  _seach_blockx_191_in_do = _net_575;
   assign  _seach_blockx_191_p_reset = p_reset;
   assign  _seach_blockx_191_m_clock = m_clock;
   assign  _seach_blockx_190_map_block = data_in235;
   assign  _seach_blockx_190_now = 10'b0011101011;
   assign  _seach_blockx_190_in_do = _net_572;
   assign  _seach_blockx_190_p_reset = p_reset;
   assign  _seach_blockx_190_m_clock = m_clock;
   assign  _seach_blockx_189_map_block = data_in234;
   assign  _seach_blockx_189_now = 10'b0011101010;
   assign  _seach_blockx_189_in_do = _net_569;
   assign  _seach_blockx_189_p_reset = p_reset;
   assign  _seach_blockx_189_m_clock = m_clock;
   assign  _seach_blockx_188_map_block = data_in233;
   assign  _seach_blockx_188_now = 10'b0011101001;
   assign  _seach_blockx_188_in_do = _net_566;
   assign  _seach_blockx_188_p_reset = p_reset;
   assign  _seach_blockx_188_m_clock = m_clock;
   assign  _seach_blockx_187_map_block = data_in232;
   assign  _seach_blockx_187_now = 10'b0011101000;
   assign  _seach_blockx_187_in_do = _net_563;
   assign  _seach_blockx_187_p_reset = p_reset;
   assign  _seach_blockx_187_m_clock = m_clock;
   assign  _seach_blockx_186_map_block = data_in231;
   assign  _seach_blockx_186_now = 10'b0011100111;
   assign  _seach_blockx_186_in_do = _net_560;
   assign  _seach_blockx_186_p_reset = p_reset;
   assign  _seach_blockx_186_m_clock = m_clock;
   assign  _seach_blockx_185_map_block = data_in230;
   assign  _seach_blockx_185_now = 10'b0011100110;
   assign  _seach_blockx_185_in_do = _net_557;
   assign  _seach_blockx_185_p_reset = p_reset;
   assign  _seach_blockx_185_m_clock = m_clock;
   assign  _seach_blockx_184_map_block = data_in229;
   assign  _seach_blockx_184_now = 10'b0011100101;
   assign  _seach_blockx_184_in_do = _net_554;
   assign  _seach_blockx_184_p_reset = p_reset;
   assign  _seach_blockx_184_m_clock = m_clock;
   assign  _seach_blockx_183_map_block = data_in228;
   assign  _seach_blockx_183_now = 10'b0011100100;
   assign  _seach_blockx_183_in_do = _net_551;
   assign  _seach_blockx_183_p_reset = p_reset;
   assign  _seach_blockx_183_m_clock = m_clock;
   assign  _seach_blockx_182_map_block = data_in227;
   assign  _seach_blockx_182_now = 10'b0011100011;
   assign  _seach_blockx_182_in_do = _net_548;
   assign  _seach_blockx_182_p_reset = p_reset;
   assign  _seach_blockx_182_m_clock = m_clock;
   assign  _seach_blockx_181_map_block = data_in226;
   assign  _seach_blockx_181_now = 10'b0011100010;
   assign  _seach_blockx_181_in_do = _net_545;
   assign  _seach_blockx_181_p_reset = p_reset;
   assign  _seach_blockx_181_m_clock = m_clock;
   assign  _seach_blockx_180_map_block = data_in225;
   assign  _seach_blockx_180_now = 10'b0011100001;
   assign  _seach_blockx_180_in_do = _net_542;
   assign  _seach_blockx_180_p_reset = p_reset;
   assign  _seach_blockx_180_m_clock = m_clock;
   assign  _seach_blockx_179_map_block = data_in222;
   assign  _seach_blockx_179_now = 10'b0011011110;
   assign  _seach_blockx_179_in_do = _net_539;
   assign  _seach_blockx_179_p_reset = p_reset;
   assign  _seach_blockx_179_m_clock = m_clock;
   assign  _seach_blockx_178_map_block = data_in221;
   assign  _seach_blockx_178_now = 10'b0011011101;
   assign  _seach_blockx_178_in_do = _net_536;
   assign  _seach_blockx_178_p_reset = p_reset;
   assign  _seach_blockx_178_m_clock = m_clock;
   assign  _seach_blockx_177_map_block = data_in220;
   assign  _seach_blockx_177_now = 10'b0011011100;
   assign  _seach_blockx_177_in_do = _net_533;
   assign  _seach_blockx_177_p_reset = p_reset;
   assign  _seach_blockx_177_m_clock = m_clock;
   assign  _seach_blockx_176_map_block = data_in219;
   assign  _seach_blockx_176_now = 10'b0011011011;
   assign  _seach_blockx_176_in_do = _net_530;
   assign  _seach_blockx_176_p_reset = p_reset;
   assign  _seach_blockx_176_m_clock = m_clock;
   assign  _seach_blockx_175_map_block = data_in218;
   assign  _seach_blockx_175_now = 10'b0011011010;
   assign  _seach_blockx_175_in_do = _net_527;
   assign  _seach_blockx_175_p_reset = p_reset;
   assign  _seach_blockx_175_m_clock = m_clock;
   assign  _seach_blockx_174_map_block = data_in217;
   assign  _seach_blockx_174_now = 10'b0011011001;
   assign  _seach_blockx_174_in_do = _net_524;
   assign  _seach_blockx_174_p_reset = p_reset;
   assign  _seach_blockx_174_m_clock = m_clock;
   assign  _seach_blockx_173_map_block = data_in216;
   assign  _seach_blockx_173_now = 10'b0011011000;
   assign  _seach_blockx_173_in_do = _net_521;
   assign  _seach_blockx_173_p_reset = p_reset;
   assign  _seach_blockx_173_m_clock = m_clock;
   assign  _seach_blockx_172_map_block = data_in215;
   assign  _seach_blockx_172_now = 10'b0011010111;
   assign  _seach_blockx_172_in_do = _net_518;
   assign  _seach_blockx_172_p_reset = p_reset;
   assign  _seach_blockx_172_m_clock = m_clock;
   assign  _seach_blockx_171_map_block = data_in214;
   assign  _seach_blockx_171_now = 10'b0011010110;
   assign  _seach_blockx_171_in_do = _net_515;
   assign  _seach_blockx_171_p_reset = p_reset;
   assign  _seach_blockx_171_m_clock = m_clock;
   assign  _seach_blockx_170_map_block = data_in213;
   assign  _seach_blockx_170_now = 10'b0011010101;
   assign  _seach_blockx_170_in_do = _net_512;
   assign  _seach_blockx_170_p_reset = p_reset;
   assign  _seach_blockx_170_m_clock = m_clock;
   assign  _seach_blockx_169_map_block = data_in212;
   assign  _seach_blockx_169_now = 10'b0011010100;
   assign  _seach_blockx_169_in_do = _net_509;
   assign  _seach_blockx_169_p_reset = p_reset;
   assign  _seach_blockx_169_m_clock = m_clock;
   assign  _seach_blockx_168_map_block = data_in211;
   assign  _seach_blockx_168_now = 10'b0011010011;
   assign  _seach_blockx_168_in_do = _net_506;
   assign  _seach_blockx_168_p_reset = p_reset;
   assign  _seach_blockx_168_m_clock = m_clock;
   assign  _seach_blockx_167_map_block = data_in210;
   assign  _seach_blockx_167_now = 10'b0011010010;
   assign  _seach_blockx_167_in_do = _net_503;
   assign  _seach_blockx_167_p_reset = p_reset;
   assign  _seach_blockx_167_m_clock = m_clock;
   assign  _seach_blockx_166_map_block = data_in209;
   assign  _seach_blockx_166_now = 10'b0011010001;
   assign  _seach_blockx_166_in_do = _net_500;
   assign  _seach_blockx_166_p_reset = p_reset;
   assign  _seach_blockx_166_m_clock = m_clock;
   assign  _seach_blockx_165_map_block = data_in208;
   assign  _seach_blockx_165_now = 10'b0011010000;
   assign  _seach_blockx_165_in_do = _net_497;
   assign  _seach_blockx_165_p_reset = p_reset;
   assign  _seach_blockx_165_m_clock = m_clock;
   assign  _seach_blockx_164_map_block = data_in207;
   assign  _seach_blockx_164_now = 10'b0011001111;
   assign  _seach_blockx_164_in_do = _net_494;
   assign  _seach_blockx_164_p_reset = p_reset;
   assign  _seach_blockx_164_m_clock = m_clock;
   assign  _seach_blockx_163_map_block = data_in206;
   assign  _seach_blockx_163_now = 10'b0011001110;
   assign  _seach_blockx_163_in_do = _net_491;
   assign  _seach_blockx_163_p_reset = p_reset;
   assign  _seach_blockx_163_m_clock = m_clock;
   assign  _seach_blockx_162_map_block = data_in205;
   assign  _seach_blockx_162_now = 10'b0011001101;
   assign  _seach_blockx_162_in_do = _net_488;
   assign  _seach_blockx_162_p_reset = p_reset;
   assign  _seach_blockx_162_m_clock = m_clock;
   assign  _seach_blockx_161_map_block = data_in204;
   assign  _seach_blockx_161_now = 10'b0011001100;
   assign  _seach_blockx_161_in_do = _net_485;
   assign  _seach_blockx_161_p_reset = p_reset;
   assign  _seach_blockx_161_m_clock = m_clock;
   assign  _seach_blockx_160_map_block = data_in203;
   assign  _seach_blockx_160_now = 10'b0011001011;
   assign  _seach_blockx_160_in_do = _net_482;
   assign  _seach_blockx_160_p_reset = p_reset;
   assign  _seach_blockx_160_m_clock = m_clock;
   assign  _seach_blockx_159_map_block = data_in202;
   assign  _seach_blockx_159_now = 10'b0011001010;
   assign  _seach_blockx_159_in_do = _net_479;
   assign  _seach_blockx_159_p_reset = p_reset;
   assign  _seach_blockx_159_m_clock = m_clock;
   assign  _seach_blockx_158_map_block = data_in201;
   assign  _seach_blockx_158_now = 10'b0011001001;
   assign  _seach_blockx_158_in_do = _net_476;
   assign  _seach_blockx_158_p_reset = p_reset;
   assign  _seach_blockx_158_m_clock = m_clock;
   assign  _seach_blockx_157_map_block = data_in200;
   assign  _seach_blockx_157_now = 10'b0011001000;
   assign  _seach_blockx_157_in_do = _net_473;
   assign  _seach_blockx_157_p_reset = p_reset;
   assign  _seach_blockx_157_m_clock = m_clock;
   assign  _seach_blockx_156_map_block = data_in199;
   assign  _seach_blockx_156_now = 10'b0011000111;
   assign  _seach_blockx_156_in_do = _net_470;
   assign  _seach_blockx_156_p_reset = p_reset;
   assign  _seach_blockx_156_m_clock = m_clock;
   assign  _seach_blockx_155_map_block = data_in198;
   assign  _seach_blockx_155_now = 10'b0011000110;
   assign  _seach_blockx_155_in_do = _net_467;
   assign  _seach_blockx_155_p_reset = p_reset;
   assign  _seach_blockx_155_m_clock = m_clock;
   assign  _seach_blockx_154_map_block = data_in197;
   assign  _seach_blockx_154_now = 10'b0011000101;
   assign  _seach_blockx_154_in_do = _net_464;
   assign  _seach_blockx_154_p_reset = p_reset;
   assign  _seach_blockx_154_m_clock = m_clock;
   assign  _seach_blockx_153_map_block = data_in196;
   assign  _seach_blockx_153_now = 10'b0011000100;
   assign  _seach_blockx_153_in_do = _net_461;
   assign  _seach_blockx_153_p_reset = p_reset;
   assign  _seach_blockx_153_m_clock = m_clock;
   assign  _seach_blockx_152_map_block = data_in195;
   assign  _seach_blockx_152_now = 10'b0011000011;
   assign  _seach_blockx_152_in_do = _net_458;
   assign  _seach_blockx_152_p_reset = p_reset;
   assign  _seach_blockx_152_m_clock = m_clock;
   assign  _seach_blockx_151_map_block = data_in194;
   assign  _seach_blockx_151_now = 10'b0011000010;
   assign  _seach_blockx_151_in_do = _net_455;
   assign  _seach_blockx_151_p_reset = p_reset;
   assign  _seach_blockx_151_m_clock = m_clock;
   assign  _seach_blockx_150_map_block = data_in193;
   assign  _seach_blockx_150_now = 10'b0011000001;
   assign  _seach_blockx_150_in_do = _net_452;
   assign  _seach_blockx_150_p_reset = p_reset;
   assign  _seach_blockx_150_m_clock = m_clock;
   assign  _seach_blockx_149_map_block = data_in190;
   assign  _seach_blockx_149_now = 10'b0010111110;
   assign  _seach_blockx_149_in_do = _net_449;
   assign  _seach_blockx_149_p_reset = p_reset;
   assign  _seach_blockx_149_m_clock = m_clock;
   assign  _seach_blockx_148_map_block = data_in189;
   assign  _seach_blockx_148_now = 10'b0010111101;
   assign  _seach_blockx_148_in_do = _net_446;
   assign  _seach_blockx_148_p_reset = p_reset;
   assign  _seach_blockx_148_m_clock = m_clock;
   assign  _seach_blockx_147_map_block = data_in188;
   assign  _seach_blockx_147_now = 10'b0010111100;
   assign  _seach_blockx_147_in_do = _net_443;
   assign  _seach_blockx_147_p_reset = p_reset;
   assign  _seach_blockx_147_m_clock = m_clock;
   assign  _seach_blockx_146_map_block = data_in187;
   assign  _seach_blockx_146_now = 10'b0010111011;
   assign  _seach_blockx_146_in_do = _net_440;
   assign  _seach_blockx_146_p_reset = p_reset;
   assign  _seach_blockx_146_m_clock = m_clock;
   assign  _seach_blockx_145_map_block = data_in186;
   assign  _seach_blockx_145_now = 10'b0010111010;
   assign  _seach_blockx_145_in_do = _net_437;
   assign  _seach_blockx_145_p_reset = p_reset;
   assign  _seach_blockx_145_m_clock = m_clock;
   assign  _seach_blockx_144_map_block = data_in185;
   assign  _seach_blockx_144_now = 10'b0010111001;
   assign  _seach_blockx_144_in_do = _net_434;
   assign  _seach_blockx_144_p_reset = p_reset;
   assign  _seach_blockx_144_m_clock = m_clock;
   assign  _seach_blockx_143_map_block = data_in184;
   assign  _seach_blockx_143_now = 10'b0010111000;
   assign  _seach_blockx_143_in_do = _net_431;
   assign  _seach_blockx_143_p_reset = p_reset;
   assign  _seach_blockx_143_m_clock = m_clock;
   assign  _seach_blockx_142_map_block = data_in183;
   assign  _seach_blockx_142_now = 10'b0010110111;
   assign  _seach_blockx_142_in_do = _net_428;
   assign  _seach_blockx_142_p_reset = p_reset;
   assign  _seach_blockx_142_m_clock = m_clock;
   assign  _seach_blockx_141_map_block = data_in182;
   assign  _seach_blockx_141_now = 10'b0010110110;
   assign  _seach_blockx_141_in_do = _net_425;
   assign  _seach_blockx_141_p_reset = p_reset;
   assign  _seach_blockx_141_m_clock = m_clock;
   assign  _seach_blockx_140_map_block = data_in181;
   assign  _seach_blockx_140_now = 10'b0010110101;
   assign  _seach_blockx_140_in_do = _net_422;
   assign  _seach_blockx_140_p_reset = p_reset;
   assign  _seach_blockx_140_m_clock = m_clock;
   assign  _seach_blockx_139_map_block = data_in180;
   assign  _seach_blockx_139_now = 10'b0010110100;
   assign  _seach_blockx_139_in_do = _net_419;
   assign  _seach_blockx_139_p_reset = p_reset;
   assign  _seach_blockx_139_m_clock = m_clock;
   assign  _seach_blockx_138_map_block = data_in179;
   assign  _seach_blockx_138_now = 10'b0010110011;
   assign  _seach_blockx_138_in_do = _net_416;
   assign  _seach_blockx_138_p_reset = p_reset;
   assign  _seach_blockx_138_m_clock = m_clock;
   assign  _seach_blockx_137_map_block = data_in178;
   assign  _seach_blockx_137_now = 10'b0010110010;
   assign  _seach_blockx_137_in_do = _net_413;
   assign  _seach_blockx_137_p_reset = p_reset;
   assign  _seach_blockx_137_m_clock = m_clock;
   assign  _seach_blockx_136_map_block = data_in177;
   assign  _seach_blockx_136_now = 10'b0010110001;
   assign  _seach_blockx_136_in_do = _net_410;
   assign  _seach_blockx_136_p_reset = p_reset;
   assign  _seach_blockx_136_m_clock = m_clock;
   assign  _seach_blockx_135_map_block = data_in176;
   assign  _seach_blockx_135_now = 10'b0010110000;
   assign  _seach_blockx_135_in_do = _net_407;
   assign  _seach_blockx_135_p_reset = p_reset;
   assign  _seach_blockx_135_m_clock = m_clock;
   assign  _seach_blockx_134_map_block = data_in175;
   assign  _seach_blockx_134_now = 10'b0010101111;
   assign  _seach_blockx_134_in_do = _net_404;
   assign  _seach_blockx_134_p_reset = p_reset;
   assign  _seach_blockx_134_m_clock = m_clock;
   assign  _seach_blockx_133_map_block = data_in174;
   assign  _seach_blockx_133_now = 10'b0010101110;
   assign  _seach_blockx_133_in_do = _net_401;
   assign  _seach_blockx_133_p_reset = p_reset;
   assign  _seach_blockx_133_m_clock = m_clock;
   assign  _seach_blockx_132_map_block = data_in173;
   assign  _seach_blockx_132_now = 10'b0010101101;
   assign  _seach_blockx_132_in_do = _net_398;
   assign  _seach_blockx_132_p_reset = p_reset;
   assign  _seach_blockx_132_m_clock = m_clock;
   assign  _seach_blockx_131_map_block = data_in172;
   assign  _seach_blockx_131_now = 10'b0010101100;
   assign  _seach_blockx_131_in_do = _net_395;
   assign  _seach_blockx_131_p_reset = p_reset;
   assign  _seach_blockx_131_m_clock = m_clock;
   assign  _seach_blockx_130_map_block = data_in171;
   assign  _seach_blockx_130_now = 10'b0010101011;
   assign  _seach_blockx_130_in_do = _net_392;
   assign  _seach_blockx_130_p_reset = p_reset;
   assign  _seach_blockx_130_m_clock = m_clock;
   assign  _seach_blockx_129_map_block = data_in170;
   assign  _seach_blockx_129_now = 10'b0010101010;
   assign  _seach_blockx_129_in_do = _net_389;
   assign  _seach_blockx_129_p_reset = p_reset;
   assign  _seach_blockx_129_m_clock = m_clock;
   assign  _seach_blockx_128_map_block = data_in169;
   assign  _seach_blockx_128_now = 10'b0010101001;
   assign  _seach_blockx_128_in_do = _net_386;
   assign  _seach_blockx_128_p_reset = p_reset;
   assign  _seach_blockx_128_m_clock = m_clock;
   assign  _seach_blockx_127_map_block = data_in168;
   assign  _seach_blockx_127_now = 10'b0010101000;
   assign  _seach_blockx_127_in_do = _net_383;
   assign  _seach_blockx_127_p_reset = p_reset;
   assign  _seach_blockx_127_m_clock = m_clock;
   assign  _seach_blockx_126_map_block = data_in167;
   assign  _seach_blockx_126_now = 10'b0010100111;
   assign  _seach_blockx_126_in_do = _net_380;
   assign  _seach_blockx_126_p_reset = p_reset;
   assign  _seach_blockx_126_m_clock = m_clock;
   assign  _seach_blockx_125_map_block = data_in166;
   assign  _seach_blockx_125_now = 10'b0010100110;
   assign  _seach_blockx_125_in_do = _net_377;
   assign  _seach_blockx_125_p_reset = p_reset;
   assign  _seach_blockx_125_m_clock = m_clock;
   assign  _seach_blockx_124_map_block = data_in165;
   assign  _seach_blockx_124_now = 10'b0010100101;
   assign  _seach_blockx_124_in_do = _net_374;
   assign  _seach_blockx_124_p_reset = p_reset;
   assign  _seach_blockx_124_m_clock = m_clock;
   assign  _seach_blockx_123_map_block = data_in164;
   assign  _seach_blockx_123_now = 10'b0010100100;
   assign  _seach_blockx_123_in_do = _net_371;
   assign  _seach_blockx_123_p_reset = p_reset;
   assign  _seach_blockx_123_m_clock = m_clock;
   assign  _seach_blockx_122_map_block = data_in163;
   assign  _seach_blockx_122_now = 10'b0010100011;
   assign  _seach_blockx_122_in_do = _net_368;
   assign  _seach_blockx_122_p_reset = p_reset;
   assign  _seach_blockx_122_m_clock = m_clock;
   assign  _seach_blockx_121_map_block = data_in162;
   assign  _seach_blockx_121_now = 10'b0010100010;
   assign  _seach_blockx_121_in_do = _net_365;
   assign  _seach_blockx_121_p_reset = p_reset;
   assign  _seach_blockx_121_m_clock = m_clock;
   assign  _seach_blockx_120_map_block = data_in161;
   assign  _seach_blockx_120_now = 10'b0010100001;
   assign  _seach_blockx_120_in_do = _net_362;
   assign  _seach_blockx_120_p_reset = p_reset;
   assign  _seach_blockx_120_m_clock = m_clock;
   assign  _seach_blockx_119_map_block = data_in158;
   assign  _seach_blockx_119_now = 10'b0010011110;
   assign  _seach_blockx_119_in_do = _net_359;
   assign  _seach_blockx_119_p_reset = p_reset;
   assign  _seach_blockx_119_m_clock = m_clock;
   assign  _seach_blockx_118_map_block = data_in157;
   assign  _seach_blockx_118_now = 10'b0010011101;
   assign  _seach_blockx_118_in_do = _net_356;
   assign  _seach_blockx_118_p_reset = p_reset;
   assign  _seach_blockx_118_m_clock = m_clock;
   assign  _seach_blockx_117_map_block = data_in156;
   assign  _seach_blockx_117_now = 10'b0010011100;
   assign  _seach_blockx_117_in_do = _net_353;
   assign  _seach_blockx_117_p_reset = p_reset;
   assign  _seach_blockx_117_m_clock = m_clock;
   assign  _seach_blockx_116_map_block = data_in155;
   assign  _seach_blockx_116_now = 10'b0010011011;
   assign  _seach_blockx_116_in_do = _net_350;
   assign  _seach_blockx_116_p_reset = p_reset;
   assign  _seach_blockx_116_m_clock = m_clock;
   assign  _seach_blockx_115_map_block = data_in154;
   assign  _seach_blockx_115_now = 10'b0010011010;
   assign  _seach_blockx_115_in_do = _net_347;
   assign  _seach_blockx_115_p_reset = p_reset;
   assign  _seach_blockx_115_m_clock = m_clock;
   assign  _seach_blockx_114_map_block = data_in153;
   assign  _seach_blockx_114_now = 10'b0010011001;
   assign  _seach_blockx_114_in_do = _net_344;
   assign  _seach_blockx_114_p_reset = p_reset;
   assign  _seach_blockx_114_m_clock = m_clock;
   assign  _seach_blockx_113_map_block = data_in152;
   assign  _seach_blockx_113_now = 10'b0010011000;
   assign  _seach_blockx_113_in_do = _net_341;
   assign  _seach_blockx_113_p_reset = p_reset;
   assign  _seach_blockx_113_m_clock = m_clock;
   assign  _seach_blockx_112_map_block = data_in151;
   assign  _seach_blockx_112_now = 10'b0010010111;
   assign  _seach_blockx_112_in_do = _net_338;
   assign  _seach_blockx_112_p_reset = p_reset;
   assign  _seach_blockx_112_m_clock = m_clock;
   assign  _seach_blockx_111_map_block = data_in150;
   assign  _seach_blockx_111_now = 10'b0010010110;
   assign  _seach_blockx_111_in_do = _net_335;
   assign  _seach_blockx_111_p_reset = p_reset;
   assign  _seach_blockx_111_m_clock = m_clock;
   assign  _seach_blockx_110_map_block = data_in149;
   assign  _seach_blockx_110_now = 10'b0010010101;
   assign  _seach_blockx_110_in_do = _net_332;
   assign  _seach_blockx_110_p_reset = p_reset;
   assign  _seach_blockx_110_m_clock = m_clock;
   assign  _seach_blockx_109_map_block = data_in148;
   assign  _seach_blockx_109_now = 10'b0010010100;
   assign  _seach_blockx_109_in_do = _net_329;
   assign  _seach_blockx_109_p_reset = p_reset;
   assign  _seach_blockx_109_m_clock = m_clock;
   assign  _seach_blockx_108_map_block = data_in147;
   assign  _seach_blockx_108_now = 10'b0010010011;
   assign  _seach_blockx_108_in_do = _net_326;
   assign  _seach_blockx_108_p_reset = p_reset;
   assign  _seach_blockx_108_m_clock = m_clock;
   assign  _seach_blockx_107_map_block = data_in146;
   assign  _seach_blockx_107_now = 10'b0010010010;
   assign  _seach_blockx_107_in_do = _net_323;
   assign  _seach_blockx_107_p_reset = p_reset;
   assign  _seach_blockx_107_m_clock = m_clock;
   assign  _seach_blockx_106_map_block = data_in145;
   assign  _seach_blockx_106_now = 10'b0010010001;
   assign  _seach_blockx_106_in_do = _net_320;
   assign  _seach_blockx_106_p_reset = p_reset;
   assign  _seach_blockx_106_m_clock = m_clock;
   assign  _seach_blockx_105_map_block = data_in144;
   assign  _seach_blockx_105_now = 10'b0010010000;
   assign  _seach_blockx_105_in_do = _net_317;
   assign  _seach_blockx_105_p_reset = p_reset;
   assign  _seach_blockx_105_m_clock = m_clock;
   assign  _seach_blockx_104_map_block = data_in143;
   assign  _seach_blockx_104_now = 10'b0010001111;
   assign  _seach_blockx_104_in_do = _net_314;
   assign  _seach_blockx_104_p_reset = p_reset;
   assign  _seach_blockx_104_m_clock = m_clock;
   assign  _seach_blockx_103_map_block = data_in142;
   assign  _seach_blockx_103_now = 10'b0010001110;
   assign  _seach_blockx_103_in_do = _net_311;
   assign  _seach_blockx_103_p_reset = p_reset;
   assign  _seach_blockx_103_m_clock = m_clock;
   assign  _seach_blockx_102_map_block = data_in141;
   assign  _seach_blockx_102_now = 10'b0010001101;
   assign  _seach_blockx_102_in_do = _net_308;
   assign  _seach_blockx_102_p_reset = p_reset;
   assign  _seach_blockx_102_m_clock = m_clock;
   assign  _seach_blockx_101_map_block = data_in140;
   assign  _seach_blockx_101_now = 10'b0010001100;
   assign  _seach_blockx_101_in_do = _net_305;
   assign  _seach_blockx_101_p_reset = p_reset;
   assign  _seach_blockx_101_m_clock = m_clock;
   assign  _seach_blockx_100_map_block = data_in139;
   assign  _seach_blockx_100_now = 10'b0010001011;
   assign  _seach_blockx_100_in_do = _net_302;
   assign  _seach_blockx_100_p_reset = p_reset;
   assign  _seach_blockx_100_m_clock = m_clock;
   assign  _seach_blockx_99_map_block = data_in138;
   assign  _seach_blockx_99_now = 10'b0010001010;
   assign  _seach_blockx_99_in_do = _net_299;
   assign  _seach_blockx_99_p_reset = p_reset;
   assign  _seach_blockx_99_m_clock = m_clock;
   assign  _seach_blockx_98_map_block = data_in137;
   assign  _seach_blockx_98_now = 10'b0010001001;
   assign  _seach_blockx_98_in_do = _net_296;
   assign  _seach_blockx_98_p_reset = p_reset;
   assign  _seach_blockx_98_m_clock = m_clock;
   assign  _seach_blockx_97_map_block = data_in136;
   assign  _seach_blockx_97_now = 10'b0010001000;
   assign  _seach_blockx_97_in_do = _net_293;
   assign  _seach_blockx_97_p_reset = p_reset;
   assign  _seach_blockx_97_m_clock = m_clock;
   assign  _seach_blockx_96_map_block = data_in135;
   assign  _seach_blockx_96_now = 10'b0010000111;
   assign  _seach_blockx_96_in_do = _net_290;
   assign  _seach_blockx_96_p_reset = p_reset;
   assign  _seach_blockx_96_m_clock = m_clock;
   assign  _seach_blockx_95_map_block = data_in134;
   assign  _seach_blockx_95_now = 10'b0010000110;
   assign  _seach_blockx_95_in_do = _net_287;
   assign  _seach_blockx_95_p_reset = p_reset;
   assign  _seach_blockx_95_m_clock = m_clock;
   assign  _seach_blockx_94_map_block = data_in133;
   assign  _seach_blockx_94_now = 10'b0010000101;
   assign  _seach_blockx_94_in_do = _net_284;
   assign  _seach_blockx_94_p_reset = p_reset;
   assign  _seach_blockx_94_m_clock = m_clock;
   assign  _seach_blockx_93_map_block = data_in132;
   assign  _seach_blockx_93_now = 10'b0010000100;
   assign  _seach_blockx_93_in_do = _net_281;
   assign  _seach_blockx_93_p_reset = p_reset;
   assign  _seach_blockx_93_m_clock = m_clock;
   assign  _seach_blockx_92_map_block = data_in131;
   assign  _seach_blockx_92_now = 10'b0010000011;
   assign  _seach_blockx_92_in_do = _net_278;
   assign  _seach_blockx_92_p_reset = p_reset;
   assign  _seach_blockx_92_m_clock = m_clock;
   assign  _seach_blockx_91_map_block = data_in130;
   assign  _seach_blockx_91_now = 10'b0010000010;
   assign  _seach_blockx_91_in_do = _net_275;
   assign  _seach_blockx_91_p_reset = p_reset;
   assign  _seach_blockx_91_m_clock = m_clock;
   assign  _seach_blockx_90_map_block = data_in129;
   assign  _seach_blockx_90_now = 10'b0010000001;
   assign  _seach_blockx_90_in_do = _net_272;
   assign  _seach_blockx_90_p_reset = p_reset;
   assign  _seach_blockx_90_m_clock = m_clock;
   assign  _seach_blockx_89_map_block = data_in126;
   assign  _seach_blockx_89_now = 10'b0001111110;
   assign  _seach_blockx_89_in_do = _net_269;
   assign  _seach_blockx_89_p_reset = p_reset;
   assign  _seach_blockx_89_m_clock = m_clock;
   assign  _seach_blockx_88_map_block = data_in125;
   assign  _seach_blockx_88_now = 10'b0001111101;
   assign  _seach_blockx_88_in_do = _net_266;
   assign  _seach_blockx_88_p_reset = p_reset;
   assign  _seach_blockx_88_m_clock = m_clock;
   assign  _seach_blockx_87_map_block = data_in124;
   assign  _seach_blockx_87_now = 10'b0001111100;
   assign  _seach_blockx_87_in_do = _net_263;
   assign  _seach_blockx_87_p_reset = p_reset;
   assign  _seach_blockx_87_m_clock = m_clock;
   assign  _seach_blockx_86_map_block = data_in123;
   assign  _seach_blockx_86_now = 10'b0001111011;
   assign  _seach_blockx_86_in_do = _net_260;
   assign  _seach_blockx_86_p_reset = p_reset;
   assign  _seach_blockx_86_m_clock = m_clock;
   assign  _seach_blockx_85_map_block = data_in122;
   assign  _seach_blockx_85_now = 10'b0001111010;
   assign  _seach_blockx_85_in_do = _net_257;
   assign  _seach_blockx_85_p_reset = p_reset;
   assign  _seach_blockx_85_m_clock = m_clock;
   assign  _seach_blockx_84_map_block = data_in121;
   assign  _seach_blockx_84_now = 10'b0001111001;
   assign  _seach_blockx_84_in_do = _net_254;
   assign  _seach_blockx_84_p_reset = p_reset;
   assign  _seach_blockx_84_m_clock = m_clock;
   assign  _seach_blockx_83_map_block = data_in120;
   assign  _seach_blockx_83_now = 10'b0001111000;
   assign  _seach_blockx_83_in_do = _net_251;
   assign  _seach_blockx_83_p_reset = p_reset;
   assign  _seach_blockx_83_m_clock = m_clock;
   assign  _seach_blockx_82_map_block = data_in119;
   assign  _seach_blockx_82_now = 10'b0001110111;
   assign  _seach_blockx_82_in_do = _net_248;
   assign  _seach_blockx_82_p_reset = p_reset;
   assign  _seach_blockx_82_m_clock = m_clock;
   assign  _seach_blockx_81_map_block = data_in118;
   assign  _seach_blockx_81_now = 10'b0001110110;
   assign  _seach_blockx_81_in_do = _net_245;
   assign  _seach_blockx_81_p_reset = p_reset;
   assign  _seach_blockx_81_m_clock = m_clock;
   assign  _seach_blockx_80_map_block = data_in117;
   assign  _seach_blockx_80_now = 10'b0001110101;
   assign  _seach_blockx_80_in_do = _net_242;
   assign  _seach_blockx_80_p_reset = p_reset;
   assign  _seach_blockx_80_m_clock = m_clock;
   assign  _seach_blockx_79_map_block = data_in116;
   assign  _seach_blockx_79_now = 10'b0001110100;
   assign  _seach_blockx_79_in_do = _net_239;
   assign  _seach_blockx_79_p_reset = p_reset;
   assign  _seach_blockx_79_m_clock = m_clock;
   assign  _seach_blockx_78_map_block = data_in115;
   assign  _seach_blockx_78_now = 10'b0001110011;
   assign  _seach_blockx_78_in_do = _net_236;
   assign  _seach_blockx_78_p_reset = p_reset;
   assign  _seach_blockx_78_m_clock = m_clock;
   assign  _seach_blockx_77_map_block = data_in114;
   assign  _seach_blockx_77_now = 10'b0001110010;
   assign  _seach_blockx_77_in_do = _net_233;
   assign  _seach_blockx_77_p_reset = p_reset;
   assign  _seach_blockx_77_m_clock = m_clock;
   assign  _seach_blockx_76_map_block = data_in113;
   assign  _seach_blockx_76_now = 10'b0001110001;
   assign  _seach_blockx_76_in_do = _net_230;
   assign  _seach_blockx_76_p_reset = p_reset;
   assign  _seach_blockx_76_m_clock = m_clock;
   assign  _seach_blockx_75_map_block = data_in112;
   assign  _seach_blockx_75_now = 10'b0001110000;
   assign  _seach_blockx_75_in_do = _net_227;
   assign  _seach_blockx_75_p_reset = p_reset;
   assign  _seach_blockx_75_m_clock = m_clock;
   assign  _seach_blockx_74_map_block = data_in111;
   assign  _seach_blockx_74_now = 10'b0001101111;
   assign  _seach_blockx_74_in_do = _net_224;
   assign  _seach_blockx_74_p_reset = p_reset;
   assign  _seach_blockx_74_m_clock = m_clock;
   assign  _seach_blockx_73_map_block = data_in110;
   assign  _seach_blockx_73_now = 10'b0001101110;
   assign  _seach_blockx_73_in_do = _net_221;
   assign  _seach_blockx_73_p_reset = p_reset;
   assign  _seach_blockx_73_m_clock = m_clock;
   assign  _seach_blockx_72_map_block = data_in109;
   assign  _seach_blockx_72_now = 10'b0001101101;
   assign  _seach_blockx_72_in_do = _net_218;
   assign  _seach_blockx_72_p_reset = p_reset;
   assign  _seach_blockx_72_m_clock = m_clock;
   assign  _seach_blockx_71_map_block = data_in108;
   assign  _seach_blockx_71_now = 10'b0001101100;
   assign  _seach_blockx_71_in_do = _net_215;
   assign  _seach_blockx_71_p_reset = p_reset;
   assign  _seach_blockx_71_m_clock = m_clock;
   assign  _seach_blockx_70_map_block = data_in107;
   assign  _seach_blockx_70_now = 10'b0001101011;
   assign  _seach_blockx_70_in_do = _net_212;
   assign  _seach_blockx_70_p_reset = p_reset;
   assign  _seach_blockx_70_m_clock = m_clock;
   assign  _seach_blockx_69_map_block = data_in106;
   assign  _seach_blockx_69_now = 10'b0001101010;
   assign  _seach_blockx_69_in_do = _net_209;
   assign  _seach_blockx_69_p_reset = p_reset;
   assign  _seach_blockx_69_m_clock = m_clock;
   assign  _seach_blockx_68_map_block = data_in105;
   assign  _seach_blockx_68_now = 10'b0001101001;
   assign  _seach_blockx_68_in_do = _net_206;
   assign  _seach_blockx_68_p_reset = p_reset;
   assign  _seach_blockx_68_m_clock = m_clock;
   assign  _seach_blockx_67_map_block = data_in104;
   assign  _seach_blockx_67_now = 10'b0001101000;
   assign  _seach_blockx_67_in_do = _net_203;
   assign  _seach_blockx_67_p_reset = p_reset;
   assign  _seach_blockx_67_m_clock = m_clock;
   assign  _seach_blockx_66_map_block = data_in103;
   assign  _seach_blockx_66_now = 10'b0001100111;
   assign  _seach_blockx_66_in_do = _net_200;
   assign  _seach_blockx_66_p_reset = p_reset;
   assign  _seach_blockx_66_m_clock = m_clock;
   assign  _seach_blockx_65_map_block = data_in102;
   assign  _seach_blockx_65_now = 10'b0001100110;
   assign  _seach_blockx_65_in_do = _net_197;
   assign  _seach_blockx_65_p_reset = p_reset;
   assign  _seach_blockx_65_m_clock = m_clock;
   assign  _seach_blockx_64_map_block = data_in101;
   assign  _seach_blockx_64_now = 10'b0001100101;
   assign  _seach_blockx_64_in_do = _net_194;
   assign  _seach_blockx_64_p_reset = p_reset;
   assign  _seach_blockx_64_m_clock = m_clock;
   assign  _seach_blockx_63_map_block = data_in100;
   assign  _seach_blockx_63_now = 10'b0001100100;
   assign  _seach_blockx_63_in_do = _net_191;
   assign  _seach_blockx_63_p_reset = p_reset;
   assign  _seach_blockx_63_m_clock = m_clock;
   assign  _seach_blockx_62_map_block = data_in99;
   assign  _seach_blockx_62_now = 10'b0001100011;
   assign  _seach_blockx_62_in_do = _net_188;
   assign  _seach_blockx_62_p_reset = p_reset;
   assign  _seach_blockx_62_m_clock = m_clock;
   assign  _seach_blockx_61_map_block = data_in98;
   assign  _seach_blockx_61_now = 10'b0001100010;
   assign  _seach_blockx_61_in_do = _net_185;
   assign  _seach_blockx_61_p_reset = p_reset;
   assign  _seach_blockx_61_m_clock = m_clock;
   assign  _seach_blockx_60_map_block = data_in97;
   assign  _seach_blockx_60_now = 10'b0001100001;
   assign  _seach_blockx_60_in_do = _net_182;
   assign  _seach_blockx_60_p_reset = p_reset;
   assign  _seach_blockx_60_m_clock = m_clock;
   assign  _seach_blockx_59_map_block = data_in94;
   assign  _seach_blockx_59_now = 10'b0001011110;
   assign  _seach_blockx_59_in_do = _net_179;
   assign  _seach_blockx_59_p_reset = p_reset;
   assign  _seach_blockx_59_m_clock = m_clock;
   assign  _seach_blockx_58_map_block = data_in93;
   assign  _seach_blockx_58_now = 10'b0001011101;
   assign  _seach_blockx_58_in_do = _net_176;
   assign  _seach_blockx_58_p_reset = p_reset;
   assign  _seach_blockx_58_m_clock = m_clock;
   assign  _seach_blockx_57_map_block = data_in92;
   assign  _seach_blockx_57_now = 10'b0001011100;
   assign  _seach_blockx_57_in_do = _net_173;
   assign  _seach_blockx_57_p_reset = p_reset;
   assign  _seach_blockx_57_m_clock = m_clock;
   assign  _seach_blockx_56_map_block = data_in91;
   assign  _seach_blockx_56_now = 10'b0001011011;
   assign  _seach_blockx_56_in_do = _net_170;
   assign  _seach_blockx_56_p_reset = p_reset;
   assign  _seach_blockx_56_m_clock = m_clock;
   assign  _seach_blockx_55_map_block = data_in90;
   assign  _seach_blockx_55_now = 10'b0001011010;
   assign  _seach_blockx_55_in_do = _net_167;
   assign  _seach_blockx_55_p_reset = p_reset;
   assign  _seach_blockx_55_m_clock = m_clock;
   assign  _seach_blockx_54_map_block = data_in89;
   assign  _seach_blockx_54_now = 10'b0001011001;
   assign  _seach_blockx_54_in_do = _net_164;
   assign  _seach_blockx_54_p_reset = p_reset;
   assign  _seach_blockx_54_m_clock = m_clock;
   assign  _seach_blockx_53_map_block = data_in88;
   assign  _seach_blockx_53_now = 10'b0001011000;
   assign  _seach_blockx_53_in_do = _net_161;
   assign  _seach_blockx_53_p_reset = p_reset;
   assign  _seach_blockx_53_m_clock = m_clock;
   assign  _seach_blockx_52_map_block = data_in87;
   assign  _seach_blockx_52_now = 10'b0001010111;
   assign  _seach_blockx_52_in_do = _net_158;
   assign  _seach_blockx_52_p_reset = p_reset;
   assign  _seach_blockx_52_m_clock = m_clock;
   assign  _seach_blockx_51_map_block = data_in86;
   assign  _seach_blockx_51_now = 10'b0001010110;
   assign  _seach_blockx_51_in_do = _net_155;
   assign  _seach_blockx_51_p_reset = p_reset;
   assign  _seach_blockx_51_m_clock = m_clock;
   assign  _seach_blockx_50_map_block = data_in85;
   assign  _seach_blockx_50_now = 10'b0001010101;
   assign  _seach_blockx_50_in_do = _net_152;
   assign  _seach_blockx_50_p_reset = p_reset;
   assign  _seach_blockx_50_m_clock = m_clock;
   assign  _seach_blockx_49_map_block = data_in84;
   assign  _seach_blockx_49_now = 10'b0001010100;
   assign  _seach_blockx_49_in_do = _net_149;
   assign  _seach_blockx_49_p_reset = p_reset;
   assign  _seach_blockx_49_m_clock = m_clock;
   assign  _seach_blockx_48_map_block = data_in83;
   assign  _seach_blockx_48_now = 10'b0001010011;
   assign  _seach_blockx_48_in_do = _net_146;
   assign  _seach_blockx_48_p_reset = p_reset;
   assign  _seach_blockx_48_m_clock = m_clock;
   assign  _seach_blockx_47_map_block = data_in82;
   assign  _seach_blockx_47_now = 10'b0001010010;
   assign  _seach_blockx_47_in_do = _net_143;
   assign  _seach_blockx_47_p_reset = p_reset;
   assign  _seach_blockx_47_m_clock = m_clock;
   assign  _seach_blockx_46_map_block = data_in81;
   assign  _seach_blockx_46_now = 10'b0001010001;
   assign  _seach_blockx_46_in_do = _net_140;
   assign  _seach_blockx_46_p_reset = p_reset;
   assign  _seach_blockx_46_m_clock = m_clock;
   assign  _seach_blockx_45_map_block = data_in80;
   assign  _seach_blockx_45_now = 10'b0001010000;
   assign  _seach_blockx_45_in_do = _net_137;
   assign  _seach_blockx_45_p_reset = p_reset;
   assign  _seach_blockx_45_m_clock = m_clock;
   assign  _seach_blockx_44_map_block = data_in79;
   assign  _seach_blockx_44_now = 10'b0001001111;
   assign  _seach_blockx_44_in_do = _net_134;
   assign  _seach_blockx_44_p_reset = p_reset;
   assign  _seach_blockx_44_m_clock = m_clock;
   assign  _seach_blockx_43_map_block = data_in78;
   assign  _seach_blockx_43_now = 10'b0001001110;
   assign  _seach_blockx_43_in_do = _net_131;
   assign  _seach_blockx_43_p_reset = p_reset;
   assign  _seach_blockx_43_m_clock = m_clock;
   assign  _seach_blockx_42_map_block = data_in77;
   assign  _seach_blockx_42_now = 10'b0001001101;
   assign  _seach_blockx_42_in_do = _net_128;
   assign  _seach_blockx_42_p_reset = p_reset;
   assign  _seach_blockx_42_m_clock = m_clock;
   assign  _seach_blockx_41_map_block = data_in76;
   assign  _seach_blockx_41_now = 10'b0001001100;
   assign  _seach_blockx_41_in_do = _net_125;
   assign  _seach_blockx_41_p_reset = p_reset;
   assign  _seach_blockx_41_m_clock = m_clock;
   assign  _seach_blockx_40_map_block = data_in75;
   assign  _seach_blockx_40_now = 10'b0001001011;
   assign  _seach_blockx_40_in_do = _net_122;
   assign  _seach_blockx_40_p_reset = p_reset;
   assign  _seach_blockx_40_m_clock = m_clock;
   assign  _seach_blockx_39_map_block = data_in74;
   assign  _seach_blockx_39_now = 10'b0001001010;
   assign  _seach_blockx_39_in_do = _net_119;
   assign  _seach_blockx_39_p_reset = p_reset;
   assign  _seach_blockx_39_m_clock = m_clock;
   assign  _seach_blockx_38_map_block = data_in73;
   assign  _seach_blockx_38_now = 10'b0001001001;
   assign  _seach_blockx_38_in_do = _net_116;
   assign  _seach_blockx_38_p_reset = p_reset;
   assign  _seach_blockx_38_m_clock = m_clock;
   assign  _seach_blockx_37_map_block = data_in72;
   assign  _seach_blockx_37_now = 10'b0001001000;
   assign  _seach_blockx_37_in_do = _net_113;
   assign  _seach_blockx_37_p_reset = p_reset;
   assign  _seach_blockx_37_m_clock = m_clock;
   assign  _seach_blockx_36_map_block = data_in71;
   assign  _seach_blockx_36_now = 10'b0001000111;
   assign  _seach_blockx_36_in_do = _net_110;
   assign  _seach_blockx_36_p_reset = p_reset;
   assign  _seach_blockx_36_m_clock = m_clock;
   assign  _seach_blockx_35_map_block = data_in70;
   assign  _seach_blockx_35_now = 10'b0001000110;
   assign  _seach_blockx_35_in_do = _net_107;
   assign  _seach_blockx_35_p_reset = p_reset;
   assign  _seach_blockx_35_m_clock = m_clock;
   assign  _seach_blockx_34_map_block = data_in69;
   assign  _seach_blockx_34_now = 10'b0001000101;
   assign  _seach_blockx_34_in_do = _net_104;
   assign  _seach_blockx_34_p_reset = p_reset;
   assign  _seach_blockx_34_m_clock = m_clock;
   assign  _seach_blockx_33_map_block = data_in68;
   assign  _seach_blockx_33_now = 10'b0001000100;
   assign  _seach_blockx_33_in_do = _net_101;
   assign  _seach_blockx_33_p_reset = p_reset;
   assign  _seach_blockx_33_m_clock = m_clock;
   assign  _seach_blockx_32_map_block = data_in67;
   assign  _seach_blockx_32_now = 10'b0001000011;
   assign  _seach_blockx_32_in_do = _net_98;
   assign  _seach_blockx_32_p_reset = p_reset;
   assign  _seach_blockx_32_m_clock = m_clock;
   assign  _seach_blockx_31_map_block = data_in66;
   assign  _seach_blockx_31_now = 10'b0001000010;
   assign  _seach_blockx_31_in_do = _net_95;
   assign  _seach_blockx_31_p_reset = p_reset;
   assign  _seach_blockx_31_m_clock = m_clock;
   assign  _seach_blockx_30_map_block = data_in65;
   assign  _seach_blockx_30_now = 10'b0001000001;
   assign  _seach_blockx_30_in_do = _net_92;
   assign  _seach_blockx_30_p_reset = p_reset;
   assign  _seach_blockx_30_m_clock = m_clock;
   assign  _seach_blockx_29_map_block = data_in62;
   assign  _seach_blockx_29_now = 10'b0000111110;
   assign  _seach_blockx_29_in_do = _net_89;
   assign  _seach_blockx_29_p_reset = p_reset;
   assign  _seach_blockx_29_m_clock = m_clock;
   assign  _seach_blockx_28_map_block = data_in61;
   assign  _seach_blockx_28_now = 10'b0000111101;
   assign  _seach_blockx_28_in_do = _net_86;
   assign  _seach_blockx_28_p_reset = p_reset;
   assign  _seach_blockx_28_m_clock = m_clock;
   assign  _seach_blockx_27_map_block = data_in60;
   assign  _seach_blockx_27_now = 10'b0000111100;
   assign  _seach_blockx_27_in_do = _net_83;
   assign  _seach_blockx_27_p_reset = p_reset;
   assign  _seach_blockx_27_m_clock = m_clock;
   assign  _seach_blockx_26_map_block = data_in59;
   assign  _seach_blockx_26_now = 10'b0000111011;
   assign  _seach_blockx_26_in_do = _net_80;
   assign  _seach_blockx_26_p_reset = p_reset;
   assign  _seach_blockx_26_m_clock = m_clock;
   assign  _seach_blockx_25_map_block = data_in58;
   assign  _seach_blockx_25_now = 10'b0000111010;
   assign  _seach_blockx_25_in_do = _net_77;
   assign  _seach_blockx_25_p_reset = p_reset;
   assign  _seach_blockx_25_m_clock = m_clock;
   assign  _seach_blockx_24_map_block = data_in57;
   assign  _seach_blockx_24_now = 10'b0000111001;
   assign  _seach_blockx_24_in_do = _net_74;
   assign  _seach_blockx_24_p_reset = p_reset;
   assign  _seach_blockx_24_m_clock = m_clock;
   assign  _seach_blockx_23_map_block = data_in56;
   assign  _seach_blockx_23_now = 10'b0000111000;
   assign  _seach_blockx_23_in_do = _net_71;
   assign  _seach_blockx_23_p_reset = p_reset;
   assign  _seach_blockx_23_m_clock = m_clock;
   assign  _seach_blockx_22_map_block = data_in55;
   assign  _seach_blockx_22_now = 10'b0000110111;
   assign  _seach_blockx_22_in_do = _net_68;
   assign  _seach_blockx_22_p_reset = p_reset;
   assign  _seach_blockx_22_m_clock = m_clock;
   assign  _seach_blockx_21_map_block = data_in54;
   assign  _seach_blockx_21_now = 10'b0000110110;
   assign  _seach_blockx_21_in_do = _net_65;
   assign  _seach_blockx_21_p_reset = p_reset;
   assign  _seach_blockx_21_m_clock = m_clock;
   assign  _seach_blockx_20_map_block = data_in53;
   assign  _seach_blockx_20_now = 10'b0000110101;
   assign  _seach_blockx_20_in_do = _net_62;
   assign  _seach_blockx_20_p_reset = p_reset;
   assign  _seach_blockx_20_m_clock = m_clock;
   assign  _seach_blockx_19_map_block = data_in52;
   assign  _seach_blockx_19_now = 10'b0000110100;
   assign  _seach_blockx_19_in_do = _net_59;
   assign  _seach_blockx_19_p_reset = p_reset;
   assign  _seach_blockx_19_m_clock = m_clock;
   assign  _seach_blockx_18_map_block = data_in51;
   assign  _seach_blockx_18_now = 10'b0000110011;
   assign  _seach_blockx_18_in_do = _net_56;
   assign  _seach_blockx_18_p_reset = p_reset;
   assign  _seach_blockx_18_m_clock = m_clock;
   assign  _seach_blockx_17_map_block = data_in50;
   assign  _seach_blockx_17_now = 10'b0000110010;
   assign  _seach_blockx_17_in_do = _net_53;
   assign  _seach_blockx_17_p_reset = p_reset;
   assign  _seach_blockx_17_m_clock = m_clock;
   assign  _seach_blockx_16_map_block = data_in49;
   assign  _seach_blockx_16_now = 10'b0000110001;
   assign  _seach_blockx_16_in_do = _net_50;
   assign  _seach_blockx_16_p_reset = p_reset;
   assign  _seach_blockx_16_m_clock = m_clock;
   assign  _seach_blockx_15_map_block = data_in48;
   assign  _seach_blockx_15_now = 10'b0000110000;
   assign  _seach_blockx_15_in_do = _net_47;
   assign  _seach_blockx_15_p_reset = p_reset;
   assign  _seach_blockx_15_m_clock = m_clock;
   assign  _seach_blockx_14_map_block = data_in47;
   assign  _seach_blockx_14_now = 10'b0000101111;
   assign  _seach_blockx_14_in_do = _net_44;
   assign  _seach_blockx_14_p_reset = p_reset;
   assign  _seach_blockx_14_m_clock = m_clock;
   assign  _seach_blockx_13_map_block = data_in46;
   assign  _seach_blockx_13_now = 10'b0000101110;
   assign  _seach_blockx_13_in_do = _net_41;
   assign  _seach_blockx_13_p_reset = p_reset;
   assign  _seach_blockx_13_m_clock = m_clock;
   assign  _seach_blockx_12_map_block = data_in45;
   assign  _seach_blockx_12_now = 10'b0000101101;
   assign  _seach_blockx_12_in_do = _net_38;
   assign  _seach_blockx_12_p_reset = p_reset;
   assign  _seach_blockx_12_m_clock = m_clock;
   assign  _seach_blockx_11_map_block = data_in44;
   assign  _seach_blockx_11_now = 10'b0000101100;
   assign  _seach_blockx_11_in_do = _net_35;
   assign  _seach_blockx_11_p_reset = p_reset;
   assign  _seach_blockx_11_m_clock = m_clock;
   assign  _seach_blockx_10_map_block = data_in43;
   assign  _seach_blockx_10_now = 10'b0000101011;
   assign  _seach_blockx_10_in_do = _net_32;
   assign  _seach_blockx_10_p_reset = p_reset;
   assign  _seach_blockx_10_m_clock = m_clock;
   assign  _seach_blockx_9_map_block = data_in42;
   assign  _seach_blockx_9_now = 10'b0000101010;
   assign  _seach_blockx_9_in_do = _net_29;
   assign  _seach_blockx_9_p_reset = p_reset;
   assign  _seach_blockx_9_m_clock = m_clock;
   assign  _seach_blockx_8_map_block = data_in41;
   assign  _seach_blockx_8_now = 10'b0000101001;
   assign  _seach_blockx_8_in_do = _net_26;
   assign  _seach_blockx_8_p_reset = p_reset;
   assign  _seach_blockx_8_m_clock = m_clock;
   assign  _seach_blockx_7_map_block = data_in40;
   assign  _seach_blockx_7_now = 10'b0000101000;
   assign  _seach_blockx_7_in_do = _net_23;
   assign  _seach_blockx_7_p_reset = p_reset;
   assign  _seach_blockx_7_m_clock = m_clock;
   assign  _seach_blockx_6_map_block = data_in39;
   assign  _seach_blockx_6_now = 10'b0000100111;
   assign  _seach_blockx_6_in_do = _net_20;
   assign  _seach_blockx_6_p_reset = p_reset;
   assign  _seach_blockx_6_m_clock = m_clock;
   assign  _seach_blockx_5_map_block = data_in38;
   assign  _seach_blockx_5_now = 10'b0000100110;
   assign  _seach_blockx_5_in_do = _net_17;
   assign  _seach_blockx_5_p_reset = p_reset;
   assign  _seach_blockx_5_m_clock = m_clock;
   assign  _seach_blockx_4_map_block = data_in37;
   assign  _seach_blockx_4_now = 10'b0000100101;
   assign  _seach_blockx_4_in_do = _net_14;
   assign  _seach_blockx_4_p_reset = p_reset;
   assign  _seach_blockx_4_m_clock = m_clock;
   assign  _seach_blockx_3_map_block = data_in36;
   assign  _seach_blockx_3_now = 10'b0000100100;
   assign  _seach_blockx_3_in_do = _net_11;
   assign  _seach_blockx_3_p_reset = p_reset;
   assign  _seach_blockx_3_m_clock = m_clock;
   assign  _seach_blockx_2_map_block = data_in35;
   assign  _seach_blockx_2_now = 10'b0000100011;
   assign  _seach_blockx_2_in_do = _net_8;
   assign  _seach_blockx_2_p_reset = p_reset;
   assign  _seach_blockx_2_m_clock = m_clock;
   assign  _seach_blockx_1_map_block = data_in34;
   assign  _seach_blockx_1_now = 10'b0000100010;
   assign  _seach_blockx_1_in_do = _net_5;
   assign  _seach_blockx_1_p_reset = p_reset;
   assign  _seach_blockx_1_m_clock = m_clock;
   assign  _net_2 = (in_do|_reg_1);
   assign  _net_3 = (in_do|_reg_1);
   assign  _net_4 = (in_do|_reg_1);
   assign  _net_5 = (in_do|_reg_1);
   assign  _net_6 = (in_do|_reg_1);
   assign  _net_7 = (in_do|_reg_1);
   assign  _net_8 = (in_do|_reg_1);
   assign  _net_9 = (in_do|_reg_1);
   assign  _net_10 = (in_do|_reg_1);
   assign  _net_11 = (in_do|_reg_1);
   assign  _net_12 = (in_do|_reg_1);
   assign  _net_13 = (in_do|_reg_1);
   assign  _net_14 = (in_do|_reg_1);
   assign  _net_15 = (in_do|_reg_1);
   assign  _net_16 = (in_do|_reg_1);
   assign  _net_17 = (in_do|_reg_1);
   assign  _net_18 = (in_do|_reg_1);
   assign  _net_19 = (in_do|_reg_1);
   assign  _net_20 = (in_do|_reg_1);
   assign  _net_21 = (in_do|_reg_1);
   assign  _net_22 = (in_do|_reg_1);
   assign  _net_23 = (in_do|_reg_1);
   assign  _net_24 = (in_do|_reg_1);
   assign  _net_25 = (in_do|_reg_1);
   assign  _net_26 = (in_do|_reg_1);
   assign  _net_27 = (in_do|_reg_1);
   assign  _net_28 = (in_do|_reg_1);
   assign  _net_29 = (in_do|_reg_1);
   assign  _net_30 = (in_do|_reg_1);
   assign  _net_31 = (in_do|_reg_1);
   assign  _net_32 = (in_do|_reg_1);
   assign  _net_33 = (in_do|_reg_1);
   assign  _net_34 = (in_do|_reg_1);
   assign  _net_35 = (in_do|_reg_1);
   assign  _net_36 = (in_do|_reg_1);
   assign  _net_37 = (in_do|_reg_1);
   assign  _net_38 = (in_do|_reg_1);
   assign  _net_39 = (in_do|_reg_1);
   assign  _net_40 = (in_do|_reg_1);
   assign  _net_41 = (in_do|_reg_1);
   assign  _net_42 = (in_do|_reg_1);
   assign  _net_43 = (in_do|_reg_1);
   assign  _net_44 = (in_do|_reg_1);
   assign  _net_45 = (in_do|_reg_1);
   assign  _net_46 = (in_do|_reg_1);
   assign  _net_47 = (in_do|_reg_1);
   assign  _net_48 = (in_do|_reg_1);
   assign  _net_49 = (in_do|_reg_1);
   assign  _net_50 = (in_do|_reg_1);
   assign  _net_51 = (in_do|_reg_1);
   assign  _net_52 = (in_do|_reg_1);
   assign  _net_53 = (in_do|_reg_1);
   assign  _net_54 = (in_do|_reg_1);
   assign  _net_55 = (in_do|_reg_1);
   assign  _net_56 = (in_do|_reg_1);
   assign  _net_57 = (in_do|_reg_1);
   assign  _net_58 = (in_do|_reg_1);
   assign  _net_59 = (in_do|_reg_1);
   assign  _net_60 = (in_do|_reg_1);
   assign  _net_61 = (in_do|_reg_1);
   assign  _net_62 = (in_do|_reg_1);
   assign  _net_63 = (in_do|_reg_1);
   assign  _net_64 = (in_do|_reg_1);
   assign  _net_65 = (in_do|_reg_1);
   assign  _net_66 = (in_do|_reg_1);
   assign  _net_67 = (in_do|_reg_1);
   assign  _net_68 = (in_do|_reg_1);
   assign  _net_69 = (in_do|_reg_1);
   assign  _net_70 = (in_do|_reg_1);
   assign  _net_71 = (in_do|_reg_1);
   assign  _net_72 = (in_do|_reg_1);
   assign  _net_73 = (in_do|_reg_1);
   assign  _net_74 = (in_do|_reg_1);
   assign  _net_75 = (in_do|_reg_1);
   assign  _net_76 = (in_do|_reg_1);
   assign  _net_77 = (in_do|_reg_1);
   assign  _net_78 = (in_do|_reg_1);
   assign  _net_79 = (in_do|_reg_1);
   assign  _net_80 = (in_do|_reg_1);
   assign  _net_81 = (in_do|_reg_1);
   assign  _net_82 = (in_do|_reg_1);
   assign  _net_83 = (in_do|_reg_1);
   assign  _net_84 = (in_do|_reg_1);
   assign  _net_85 = (in_do|_reg_1);
   assign  _net_86 = (in_do|_reg_1);
   assign  _net_87 = (in_do|_reg_1);
   assign  _net_88 = (in_do|_reg_1);
   assign  _net_89 = (in_do|_reg_1);
   assign  _net_90 = (in_do|_reg_1);
   assign  _net_91 = (in_do|_reg_1);
   assign  _net_92 = (in_do|_reg_1);
   assign  _net_93 = (in_do|_reg_1);
   assign  _net_94 = (in_do|_reg_1);
   assign  _net_95 = (in_do|_reg_1);
   assign  _net_96 = (in_do|_reg_1);
   assign  _net_97 = (in_do|_reg_1);
   assign  _net_98 = (in_do|_reg_1);
   assign  _net_99 = (in_do|_reg_1);
   assign  _net_100 = (in_do|_reg_1);
   assign  _net_101 = (in_do|_reg_1);
   assign  _net_102 = (in_do|_reg_1);
   assign  _net_103 = (in_do|_reg_1);
   assign  _net_104 = (in_do|_reg_1);
   assign  _net_105 = (in_do|_reg_1);
   assign  _net_106 = (in_do|_reg_1);
   assign  _net_107 = (in_do|_reg_1);
   assign  _net_108 = (in_do|_reg_1);
   assign  _net_109 = (in_do|_reg_1);
   assign  _net_110 = (in_do|_reg_1);
   assign  _net_111 = (in_do|_reg_1);
   assign  _net_112 = (in_do|_reg_1);
   assign  _net_113 = (in_do|_reg_1);
   assign  _net_114 = (in_do|_reg_1);
   assign  _net_115 = (in_do|_reg_1);
   assign  _net_116 = (in_do|_reg_1);
   assign  _net_117 = (in_do|_reg_1);
   assign  _net_118 = (in_do|_reg_1);
   assign  _net_119 = (in_do|_reg_1);
   assign  _net_120 = (in_do|_reg_1);
   assign  _net_121 = (in_do|_reg_1);
   assign  _net_122 = (in_do|_reg_1);
   assign  _net_123 = (in_do|_reg_1);
   assign  _net_124 = (in_do|_reg_1);
   assign  _net_125 = (in_do|_reg_1);
   assign  _net_126 = (in_do|_reg_1);
   assign  _net_127 = (in_do|_reg_1);
   assign  _net_128 = (in_do|_reg_1);
   assign  _net_129 = (in_do|_reg_1);
   assign  _net_130 = (in_do|_reg_1);
   assign  _net_131 = (in_do|_reg_1);
   assign  _net_132 = (in_do|_reg_1);
   assign  _net_133 = (in_do|_reg_1);
   assign  _net_134 = (in_do|_reg_1);
   assign  _net_135 = (in_do|_reg_1);
   assign  _net_136 = (in_do|_reg_1);
   assign  _net_137 = (in_do|_reg_1);
   assign  _net_138 = (in_do|_reg_1);
   assign  _net_139 = (in_do|_reg_1);
   assign  _net_140 = (in_do|_reg_1);
   assign  _net_141 = (in_do|_reg_1);
   assign  _net_142 = (in_do|_reg_1);
   assign  _net_143 = (in_do|_reg_1);
   assign  _net_144 = (in_do|_reg_1);
   assign  _net_145 = (in_do|_reg_1);
   assign  _net_146 = (in_do|_reg_1);
   assign  _net_147 = (in_do|_reg_1);
   assign  _net_148 = (in_do|_reg_1);
   assign  _net_149 = (in_do|_reg_1);
   assign  _net_150 = (in_do|_reg_1);
   assign  _net_151 = (in_do|_reg_1);
   assign  _net_152 = (in_do|_reg_1);
   assign  _net_153 = (in_do|_reg_1);
   assign  _net_154 = (in_do|_reg_1);
   assign  _net_155 = (in_do|_reg_1);
   assign  _net_156 = (in_do|_reg_1);
   assign  _net_157 = (in_do|_reg_1);
   assign  _net_158 = (in_do|_reg_1);
   assign  _net_159 = (in_do|_reg_1);
   assign  _net_160 = (in_do|_reg_1);
   assign  _net_161 = (in_do|_reg_1);
   assign  _net_162 = (in_do|_reg_1);
   assign  _net_163 = (in_do|_reg_1);
   assign  _net_164 = (in_do|_reg_1);
   assign  _net_165 = (in_do|_reg_1);
   assign  _net_166 = (in_do|_reg_1);
   assign  _net_167 = (in_do|_reg_1);
   assign  _net_168 = (in_do|_reg_1);
   assign  _net_169 = (in_do|_reg_1);
   assign  _net_170 = (in_do|_reg_1);
   assign  _net_171 = (in_do|_reg_1);
   assign  _net_172 = (in_do|_reg_1);
   assign  _net_173 = (in_do|_reg_1);
   assign  _net_174 = (in_do|_reg_1);
   assign  _net_175 = (in_do|_reg_1);
   assign  _net_176 = (in_do|_reg_1);
   assign  _net_177 = (in_do|_reg_1);
   assign  _net_178 = (in_do|_reg_1);
   assign  _net_179 = (in_do|_reg_1);
   assign  _net_180 = (in_do|_reg_1);
   assign  _net_181 = (in_do|_reg_1);
   assign  _net_182 = (in_do|_reg_1);
   assign  _net_183 = (in_do|_reg_1);
   assign  _net_184 = (in_do|_reg_1);
   assign  _net_185 = (in_do|_reg_1);
   assign  _net_186 = (in_do|_reg_1);
   assign  _net_187 = (in_do|_reg_1);
   assign  _net_188 = (in_do|_reg_1);
   assign  _net_189 = (in_do|_reg_1);
   assign  _net_190 = (in_do|_reg_1);
   assign  _net_191 = (in_do|_reg_1);
   assign  _net_192 = (in_do|_reg_1);
   assign  _net_193 = (in_do|_reg_1);
   assign  _net_194 = (in_do|_reg_1);
   assign  _net_195 = (in_do|_reg_1);
   assign  _net_196 = (in_do|_reg_1);
   assign  _net_197 = (in_do|_reg_1);
   assign  _net_198 = (in_do|_reg_1);
   assign  _net_199 = (in_do|_reg_1);
   assign  _net_200 = (in_do|_reg_1);
   assign  _net_201 = (in_do|_reg_1);
   assign  _net_202 = (in_do|_reg_1);
   assign  _net_203 = (in_do|_reg_1);
   assign  _net_204 = (in_do|_reg_1);
   assign  _net_205 = (in_do|_reg_1);
   assign  _net_206 = (in_do|_reg_1);
   assign  _net_207 = (in_do|_reg_1);
   assign  _net_208 = (in_do|_reg_1);
   assign  _net_209 = (in_do|_reg_1);
   assign  _net_210 = (in_do|_reg_1);
   assign  _net_211 = (in_do|_reg_1);
   assign  _net_212 = (in_do|_reg_1);
   assign  _net_213 = (in_do|_reg_1);
   assign  _net_214 = (in_do|_reg_1);
   assign  _net_215 = (in_do|_reg_1);
   assign  _net_216 = (in_do|_reg_1);
   assign  _net_217 = (in_do|_reg_1);
   assign  _net_218 = (in_do|_reg_1);
   assign  _net_219 = (in_do|_reg_1);
   assign  _net_220 = (in_do|_reg_1);
   assign  _net_221 = (in_do|_reg_1);
   assign  _net_222 = (in_do|_reg_1);
   assign  _net_223 = (in_do|_reg_1);
   assign  _net_224 = (in_do|_reg_1);
   assign  _net_225 = (in_do|_reg_1);
   assign  _net_226 = (in_do|_reg_1);
   assign  _net_227 = (in_do|_reg_1);
   assign  _net_228 = (in_do|_reg_1);
   assign  _net_229 = (in_do|_reg_1);
   assign  _net_230 = (in_do|_reg_1);
   assign  _net_231 = (in_do|_reg_1);
   assign  _net_232 = (in_do|_reg_1);
   assign  _net_233 = (in_do|_reg_1);
   assign  _net_234 = (in_do|_reg_1);
   assign  _net_235 = (in_do|_reg_1);
   assign  _net_236 = (in_do|_reg_1);
   assign  _net_237 = (in_do|_reg_1);
   assign  _net_238 = (in_do|_reg_1);
   assign  _net_239 = (in_do|_reg_1);
   assign  _net_240 = (in_do|_reg_1);
   assign  _net_241 = (in_do|_reg_1);
   assign  _net_242 = (in_do|_reg_1);
   assign  _net_243 = (in_do|_reg_1);
   assign  _net_244 = (in_do|_reg_1);
   assign  _net_245 = (in_do|_reg_1);
   assign  _net_246 = (in_do|_reg_1);
   assign  _net_247 = (in_do|_reg_1);
   assign  _net_248 = (in_do|_reg_1);
   assign  _net_249 = (in_do|_reg_1);
   assign  _net_250 = (in_do|_reg_1);
   assign  _net_251 = (in_do|_reg_1);
   assign  _net_252 = (in_do|_reg_1);
   assign  _net_253 = (in_do|_reg_1);
   assign  _net_254 = (in_do|_reg_1);
   assign  _net_255 = (in_do|_reg_1);
   assign  _net_256 = (in_do|_reg_1);
   assign  _net_257 = (in_do|_reg_1);
   assign  _net_258 = (in_do|_reg_1);
   assign  _net_259 = (in_do|_reg_1);
   assign  _net_260 = (in_do|_reg_1);
   assign  _net_261 = (in_do|_reg_1);
   assign  _net_262 = (in_do|_reg_1);
   assign  _net_263 = (in_do|_reg_1);
   assign  _net_264 = (in_do|_reg_1);
   assign  _net_265 = (in_do|_reg_1);
   assign  _net_266 = (in_do|_reg_1);
   assign  _net_267 = (in_do|_reg_1);
   assign  _net_268 = (in_do|_reg_1);
   assign  _net_269 = (in_do|_reg_1);
   assign  _net_270 = (in_do|_reg_1);
   assign  _net_271 = (in_do|_reg_1);
   assign  _net_272 = (in_do|_reg_1);
   assign  _net_273 = (in_do|_reg_1);
   assign  _net_274 = (in_do|_reg_1);
   assign  _net_275 = (in_do|_reg_1);
   assign  _net_276 = (in_do|_reg_1);
   assign  _net_277 = (in_do|_reg_1);
   assign  _net_278 = (in_do|_reg_1);
   assign  _net_279 = (in_do|_reg_1);
   assign  _net_280 = (in_do|_reg_1);
   assign  _net_281 = (in_do|_reg_1);
   assign  _net_282 = (in_do|_reg_1);
   assign  _net_283 = (in_do|_reg_1);
   assign  _net_284 = (in_do|_reg_1);
   assign  _net_285 = (in_do|_reg_1);
   assign  _net_286 = (in_do|_reg_1);
   assign  _net_287 = (in_do|_reg_1);
   assign  _net_288 = (in_do|_reg_1);
   assign  _net_289 = (in_do|_reg_1);
   assign  _net_290 = (in_do|_reg_1);
   assign  _net_291 = (in_do|_reg_1);
   assign  _net_292 = (in_do|_reg_1);
   assign  _net_293 = (in_do|_reg_1);
   assign  _net_294 = (in_do|_reg_1);
   assign  _net_295 = (in_do|_reg_1);
   assign  _net_296 = (in_do|_reg_1);
   assign  _net_297 = (in_do|_reg_1);
   assign  _net_298 = (in_do|_reg_1);
   assign  _net_299 = (in_do|_reg_1);
   assign  _net_300 = (in_do|_reg_1);
   assign  _net_301 = (in_do|_reg_1);
   assign  _net_302 = (in_do|_reg_1);
   assign  _net_303 = (in_do|_reg_1);
   assign  _net_304 = (in_do|_reg_1);
   assign  _net_305 = (in_do|_reg_1);
   assign  _net_306 = (in_do|_reg_1);
   assign  _net_307 = (in_do|_reg_1);
   assign  _net_308 = (in_do|_reg_1);
   assign  _net_309 = (in_do|_reg_1);
   assign  _net_310 = (in_do|_reg_1);
   assign  _net_311 = (in_do|_reg_1);
   assign  _net_312 = (in_do|_reg_1);
   assign  _net_313 = (in_do|_reg_1);
   assign  _net_314 = (in_do|_reg_1);
   assign  _net_315 = (in_do|_reg_1);
   assign  _net_316 = (in_do|_reg_1);
   assign  _net_317 = (in_do|_reg_1);
   assign  _net_318 = (in_do|_reg_1);
   assign  _net_319 = (in_do|_reg_1);
   assign  _net_320 = (in_do|_reg_1);
   assign  _net_321 = (in_do|_reg_1);
   assign  _net_322 = (in_do|_reg_1);
   assign  _net_323 = (in_do|_reg_1);
   assign  _net_324 = (in_do|_reg_1);
   assign  _net_325 = (in_do|_reg_1);
   assign  _net_326 = (in_do|_reg_1);
   assign  _net_327 = (in_do|_reg_1);
   assign  _net_328 = (in_do|_reg_1);
   assign  _net_329 = (in_do|_reg_1);
   assign  _net_330 = (in_do|_reg_1);
   assign  _net_331 = (in_do|_reg_1);
   assign  _net_332 = (in_do|_reg_1);
   assign  _net_333 = (in_do|_reg_1);
   assign  _net_334 = (in_do|_reg_1);
   assign  _net_335 = (in_do|_reg_1);
   assign  _net_336 = (in_do|_reg_1);
   assign  _net_337 = (in_do|_reg_1);
   assign  _net_338 = (in_do|_reg_1);
   assign  _net_339 = (in_do|_reg_1);
   assign  _net_340 = (in_do|_reg_1);
   assign  _net_341 = (in_do|_reg_1);
   assign  _net_342 = (in_do|_reg_1);
   assign  _net_343 = (in_do|_reg_1);
   assign  _net_344 = (in_do|_reg_1);
   assign  _net_345 = (in_do|_reg_1);
   assign  _net_346 = (in_do|_reg_1);
   assign  _net_347 = (in_do|_reg_1);
   assign  _net_348 = (in_do|_reg_1);
   assign  _net_349 = (in_do|_reg_1);
   assign  _net_350 = (in_do|_reg_1);
   assign  _net_351 = (in_do|_reg_1);
   assign  _net_352 = (in_do|_reg_1);
   assign  _net_353 = (in_do|_reg_1);
   assign  _net_354 = (in_do|_reg_1);
   assign  _net_355 = (in_do|_reg_1);
   assign  _net_356 = (in_do|_reg_1);
   assign  _net_357 = (in_do|_reg_1);
   assign  _net_358 = (in_do|_reg_1);
   assign  _net_359 = (in_do|_reg_1);
   assign  _net_360 = (in_do|_reg_1);
   assign  _net_361 = (in_do|_reg_1);
   assign  _net_362 = (in_do|_reg_1);
   assign  _net_363 = (in_do|_reg_1);
   assign  _net_364 = (in_do|_reg_1);
   assign  _net_365 = (in_do|_reg_1);
   assign  _net_366 = (in_do|_reg_1);
   assign  _net_367 = (in_do|_reg_1);
   assign  _net_368 = (in_do|_reg_1);
   assign  _net_369 = (in_do|_reg_1);
   assign  _net_370 = (in_do|_reg_1);
   assign  _net_371 = (in_do|_reg_1);
   assign  _net_372 = (in_do|_reg_1);
   assign  _net_373 = (in_do|_reg_1);
   assign  _net_374 = (in_do|_reg_1);
   assign  _net_375 = (in_do|_reg_1);
   assign  _net_376 = (in_do|_reg_1);
   assign  _net_377 = (in_do|_reg_1);
   assign  _net_378 = (in_do|_reg_1);
   assign  _net_379 = (in_do|_reg_1);
   assign  _net_380 = (in_do|_reg_1);
   assign  _net_381 = (in_do|_reg_1);
   assign  _net_382 = (in_do|_reg_1);
   assign  _net_383 = (in_do|_reg_1);
   assign  _net_384 = (in_do|_reg_1);
   assign  _net_385 = (in_do|_reg_1);
   assign  _net_386 = (in_do|_reg_1);
   assign  _net_387 = (in_do|_reg_1);
   assign  _net_388 = (in_do|_reg_1);
   assign  _net_389 = (in_do|_reg_1);
   assign  _net_390 = (in_do|_reg_1);
   assign  _net_391 = (in_do|_reg_1);
   assign  _net_392 = (in_do|_reg_1);
   assign  _net_393 = (in_do|_reg_1);
   assign  _net_394 = (in_do|_reg_1);
   assign  _net_395 = (in_do|_reg_1);
   assign  _net_396 = (in_do|_reg_1);
   assign  _net_397 = (in_do|_reg_1);
   assign  _net_398 = (in_do|_reg_1);
   assign  _net_399 = (in_do|_reg_1);
   assign  _net_400 = (in_do|_reg_1);
   assign  _net_401 = (in_do|_reg_1);
   assign  _net_402 = (in_do|_reg_1);
   assign  _net_403 = (in_do|_reg_1);
   assign  _net_404 = (in_do|_reg_1);
   assign  _net_405 = (in_do|_reg_1);
   assign  _net_406 = (in_do|_reg_1);
   assign  _net_407 = (in_do|_reg_1);
   assign  _net_408 = (in_do|_reg_1);
   assign  _net_409 = (in_do|_reg_1);
   assign  _net_410 = (in_do|_reg_1);
   assign  _net_411 = (in_do|_reg_1);
   assign  _net_412 = (in_do|_reg_1);
   assign  _net_413 = (in_do|_reg_1);
   assign  _net_414 = (in_do|_reg_1);
   assign  _net_415 = (in_do|_reg_1);
   assign  _net_416 = (in_do|_reg_1);
   assign  _net_417 = (in_do|_reg_1);
   assign  _net_418 = (in_do|_reg_1);
   assign  _net_419 = (in_do|_reg_1);
   assign  _net_420 = (in_do|_reg_1);
   assign  _net_421 = (in_do|_reg_1);
   assign  _net_422 = (in_do|_reg_1);
   assign  _net_423 = (in_do|_reg_1);
   assign  _net_424 = (in_do|_reg_1);
   assign  _net_425 = (in_do|_reg_1);
   assign  _net_426 = (in_do|_reg_1);
   assign  _net_427 = (in_do|_reg_1);
   assign  _net_428 = (in_do|_reg_1);
   assign  _net_429 = (in_do|_reg_1);
   assign  _net_430 = (in_do|_reg_1);
   assign  _net_431 = (in_do|_reg_1);
   assign  _net_432 = (in_do|_reg_1);
   assign  _net_433 = (in_do|_reg_1);
   assign  _net_434 = (in_do|_reg_1);
   assign  _net_435 = (in_do|_reg_1);
   assign  _net_436 = (in_do|_reg_1);
   assign  _net_437 = (in_do|_reg_1);
   assign  _net_438 = (in_do|_reg_1);
   assign  _net_439 = (in_do|_reg_1);
   assign  _net_440 = (in_do|_reg_1);
   assign  _net_441 = (in_do|_reg_1);
   assign  _net_442 = (in_do|_reg_1);
   assign  _net_443 = (in_do|_reg_1);
   assign  _net_444 = (in_do|_reg_1);
   assign  _net_445 = (in_do|_reg_1);
   assign  _net_446 = (in_do|_reg_1);
   assign  _net_447 = (in_do|_reg_1);
   assign  _net_448 = (in_do|_reg_1);
   assign  _net_449 = (in_do|_reg_1);
   assign  _net_450 = (in_do|_reg_1);
   assign  _net_451 = (in_do|_reg_1);
   assign  _net_452 = (in_do|_reg_1);
   assign  _net_453 = (in_do|_reg_1);
   assign  _net_454 = (in_do|_reg_1);
   assign  _net_455 = (in_do|_reg_1);
   assign  _net_456 = (in_do|_reg_1);
   assign  _net_457 = (in_do|_reg_1);
   assign  _net_458 = (in_do|_reg_1);
   assign  _net_459 = (in_do|_reg_1);
   assign  _net_460 = (in_do|_reg_1);
   assign  _net_461 = (in_do|_reg_1);
   assign  _net_462 = (in_do|_reg_1);
   assign  _net_463 = (in_do|_reg_1);
   assign  _net_464 = (in_do|_reg_1);
   assign  _net_465 = (in_do|_reg_1);
   assign  _net_466 = (in_do|_reg_1);
   assign  _net_467 = (in_do|_reg_1);
   assign  _net_468 = (in_do|_reg_1);
   assign  _net_469 = (in_do|_reg_1);
   assign  _net_470 = (in_do|_reg_1);
   assign  _net_471 = (in_do|_reg_1);
   assign  _net_472 = (in_do|_reg_1);
   assign  _net_473 = (in_do|_reg_1);
   assign  _net_474 = (in_do|_reg_1);
   assign  _net_475 = (in_do|_reg_1);
   assign  _net_476 = (in_do|_reg_1);
   assign  _net_477 = (in_do|_reg_1);
   assign  _net_478 = (in_do|_reg_1);
   assign  _net_479 = (in_do|_reg_1);
   assign  _net_480 = (in_do|_reg_1);
   assign  _net_481 = (in_do|_reg_1);
   assign  _net_482 = (in_do|_reg_1);
   assign  _net_483 = (in_do|_reg_1);
   assign  _net_484 = (in_do|_reg_1);
   assign  _net_485 = (in_do|_reg_1);
   assign  _net_486 = (in_do|_reg_1);
   assign  _net_487 = (in_do|_reg_1);
   assign  _net_488 = (in_do|_reg_1);
   assign  _net_489 = (in_do|_reg_1);
   assign  _net_490 = (in_do|_reg_1);
   assign  _net_491 = (in_do|_reg_1);
   assign  _net_492 = (in_do|_reg_1);
   assign  _net_493 = (in_do|_reg_1);
   assign  _net_494 = (in_do|_reg_1);
   assign  _net_495 = (in_do|_reg_1);
   assign  _net_496 = (in_do|_reg_1);
   assign  _net_497 = (in_do|_reg_1);
   assign  _net_498 = (in_do|_reg_1);
   assign  _net_499 = (in_do|_reg_1);
   assign  _net_500 = (in_do|_reg_1);
   assign  _net_501 = (in_do|_reg_1);
   assign  _net_502 = (in_do|_reg_1);
   assign  _net_503 = (in_do|_reg_1);
   assign  _net_504 = (in_do|_reg_1);
   assign  _net_505 = (in_do|_reg_1);
   assign  _net_506 = (in_do|_reg_1);
   assign  _net_507 = (in_do|_reg_1);
   assign  _net_508 = (in_do|_reg_1);
   assign  _net_509 = (in_do|_reg_1);
   assign  _net_510 = (in_do|_reg_1);
   assign  _net_511 = (in_do|_reg_1);
   assign  _net_512 = (in_do|_reg_1);
   assign  _net_513 = (in_do|_reg_1);
   assign  _net_514 = (in_do|_reg_1);
   assign  _net_515 = (in_do|_reg_1);
   assign  _net_516 = (in_do|_reg_1);
   assign  _net_517 = (in_do|_reg_1);
   assign  _net_518 = (in_do|_reg_1);
   assign  _net_519 = (in_do|_reg_1);
   assign  _net_520 = (in_do|_reg_1);
   assign  _net_521 = (in_do|_reg_1);
   assign  _net_522 = (in_do|_reg_1);
   assign  _net_523 = (in_do|_reg_1);
   assign  _net_524 = (in_do|_reg_1);
   assign  _net_525 = (in_do|_reg_1);
   assign  _net_526 = (in_do|_reg_1);
   assign  _net_527 = (in_do|_reg_1);
   assign  _net_528 = (in_do|_reg_1);
   assign  _net_529 = (in_do|_reg_1);
   assign  _net_530 = (in_do|_reg_1);
   assign  _net_531 = (in_do|_reg_1);
   assign  _net_532 = (in_do|_reg_1);
   assign  _net_533 = (in_do|_reg_1);
   assign  _net_534 = (in_do|_reg_1);
   assign  _net_535 = (in_do|_reg_1);
   assign  _net_536 = (in_do|_reg_1);
   assign  _net_537 = (in_do|_reg_1);
   assign  _net_538 = (in_do|_reg_1);
   assign  _net_539 = (in_do|_reg_1);
   assign  _net_540 = (in_do|_reg_1);
   assign  _net_541 = (in_do|_reg_1);
   assign  _net_542 = (in_do|_reg_1);
   assign  _net_543 = (in_do|_reg_1);
   assign  _net_544 = (in_do|_reg_1);
   assign  _net_545 = (in_do|_reg_1);
   assign  _net_546 = (in_do|_reg_1);
   assign  _net_547 = (in_do|_reg_1);
   assign  _net_548 = (in_do|_reg_1);
   assign  _net_549 = (in_do|_reg_1);
   assign  _net_550 = (in_do|_reg_1);
   assign  _net_551 = (in_do|_reg_1);
   assign  _net_552 = (in_do|_reg_1);
   assign  _net_553 = (in_do|_reg_1);
   assign  _net_554 = (in_do|_reg_1);
   assign  _net_555 = (in_do|_reg_1);
   assign  _net_556 = (in_do|_reg_1);
   assign  _net_557 = (in_do|_reg_1);
   assign  _net_558 = (in_do|_reg_1);
   assign  _net_559 = (in_do|_reg_1);
   assign  _net_560 = (in_do|_reg_1);
   assign  _net_561 = (in_do|_reg_1);
   assign  _net_562 = (in_do|_reg_1);
   assign  _net_563 = (in_do|_reg_1);
   assign  _net_564 = (in_do|_reg_1);
   assign  _net_565 = (in_do|_reg_1);
   assign  _net_566 = (in_do|_reg_1);
   assign  _net_567 = (in_do|_reg_1);
   assign  _net_568 = (in_do|_reg_1);
   assign  _net_569 = (in_do|_reg_1);
   assign  _net_570 = (in_do|_reg_1);
   assign  _net_571 = (in_do|_reg_1);
   assign  _net_572 = (in_do|_reg_1);
   assign  _net_573 = (in_do|_reg_1);
   assign  _net_574 = (in_do|_reg_1);
   assign  _net_575 = (in_do|_reg_1);
   assign  _net_576 = (in_do|_reg_1);
   assign  _net_577 = (in_do|_reg_1);
   assign  _net_578 = (in_do|_reg_1);
   assign  _net_579 = (in_do|_reg_1);
   assign  _net_580 = (in_do|_reg_1);
   assign  _net_581 = (in_do|_reg_1);
   assign  _net_582 = (in_do|_reg_1);
   assign  _net_583 = (in_do|_reg_1);
   assign  _net_584 = (in_do|_reg_1);
   assign  _net_585 = (in_do|_reg_1);
   assign  _net_586 = (in_do|_reg_1);
   assign  _net_587 = (in_do|_reg_1);
   assign  _net_588 = (in_do|_reg_1);
   assign  _net_589 = (in_do|_reg_1);
   assign  _net_590 = (in_do|_reg_1);
   assign  _net_591 = (in_do|_reg_1);
   assign  _net_592 = (in_do|_reg_1);
   assign  _net_593 = (in_do|_reg_1);
   assign  _net_594 = (in_do|_reg_1);
   assign  _net_595 = (in_do|_reg_1);
   assign  _net_596 = (in_do|_reg_1);
   assign  _net_597 = (in_do|_reg_1);
   assign  _net_598 = (in_do|_reg_1);
   assign  _net_599 = (in_do|_reg_1);
   assign  _net_600 = (in_do|_reg_1);
   assign  _net_601 = (in_do|_reg_1);
   assign  _net_602 = (in_do|_reg_1);
   assign  _net_603 = (in_do|_reg_1);
   assign  _net_604 = (in_do|_reg_1);
   assign  _net_605 = (in_do|_reg_1);
   assign  _net_606 = (in_do|_reg_1);
   assign  _net_607 = (in_do|_reg_1);
   assign  _net_608 = (in_do|_reg_1);
   assign  _net_609 = (in_do|_reg_1);
   assign  _net_610 = (in_do|_reg_1);
   assign  _net_611 = (in_do|_reg_1);
   assign  _net_612 = (in_do|_reg_1);
   assign  _net_613 = (in_do|_reg_1);
   assign  _net_614 = (in_do|_reg_1);
   assign  _net_615 = (in_do|_reg_1);
   assign  _net_616 = (in_do|_reg_1);
   assign  _net_617 = (in_do|_reg_1);
   assign  _net_618 = (in_do|_reg_1);
   assign  _net_619 = (in_do|_reg_1);
   assign  _net_620 = (in_do|_reg_1);
   assign  _net_621 = (in_do|_reg_1);
   assign  _net_622 = (in_do|_reg_1);
   assign  _net_623 = (in_do|_reg_1);
   assign  _net_624 = (in_do|_reg_1);
   assign  _net_625 = (in_do|_reg_1);
   assign  _net_626 = (in_do|_reg_1);
   assign  _net_627 = (in_do|_reg_1);
   assign  _net_628 = (in_do|_reg_1);
   assign  _net_629 = (in_do|_reg_1);
   assign  _net_630 = (in_do|_reg_1);
   assign  _net_631 = (in_do|_reg_1);
   assign  _net_632 = (in_do|_reg_1);
   assign  _net_633 = (in_do|_reg_1);
   assign  _net_634 = (in_do|_reg_1);
   assign  _net_635 = (in_do|_reg_1);
   assign  _net_636 = (in_do|_reg_1);
   assign  _net_637 = (in_do|_reg_1);
   assign  _net_638 = (in_do|_reg_1);
   assign  _net_639 = (in_do|_reg_1);
   assign  _net_640 = (in_do|_reg_1);
   assign  _net_641 = (in_do|_reg_1);
   assign  _net_642 = (in_do|_reg_1);
   assign  _net_643 = (in_do|_reg_1);
   assign  _net_644 = (in_do|_reg_1);
   assign  _net_645 = (in_do|_reg_1);
   assign  _net_646 = (in_do|_reg_1);
   assign  _net_647 = (in_do|_reg_1);
   assign  _net_648 = (in_do|_reg_1);
   assign  _net_649 = (in_do|_reg_1);
   assign  _net_650 = (in_do|_reg_1);
   assign  _net_651 = (in_do|_reg_1);
   assign  _net_652 = (in_do|_reg_1);
   assign  _net_653 = (in_do|_reg_1);
   assign  _net_654 = (in_do|_reg_1);
   assign  _net_655 = (in_do|_reg_1);
   assign  _net_656 = (in_do|_reg_1);
   assign  _net_657 = (in_do|_reg_1);
   assign  _net_658 = (in_do|_reg_1);
   assign  _net_659 = (in_do|_reg_1);
   assign  _net_660 = (in_do|_reg_1);
   assign  _net_661 = (in_do|_reg_1);
   assign  _net_662 = (in_do|_reg_1);
   assign  _net_663 = (in_do|_reg_1);
   assign  _net_664 = (in_do|_reg_1);
   assign  _net_665 = (in_do|_reg_1);
   assign  _net_666 = (in_do|_reg_1);
   assign  _net_667 = (in_do|_reg_1);
   assign  _net_668 = (in_do|_reg_1);
   assign  _net_669 = (in_do|_reg_1);
   assign  _net_670 = (in_do|_reg_1);
   assign  _net_671 = (in_do|_reg_1);
   assign  _net_672 = (in_do|_reg_1);
   assign  _net_673 = (in_do|_reg_1);
   assign  _net_674 = (in_do|_reg_1);
   assign  _net_675 = (in_do|_reg_1);
   assign  _net_676 = (in_do|_reg_1);
   assign  _net_677 = (in_do|_reg_1);
   assign  _net_678 = (in_do|_reg_1);
   assign  _net_679 = (in_do|_reg_1);
   assign  _net_680 = (in_do|_reg_1);
   assign  _net_681 = (in_do|_reg_1);
   assign  _net_682 = (in_do|_reg_1);
   assign  _net_683 = (in_do|_reg_1);
   assign  _net_684 = (in_do|_reg_1);
   assign  _net_685 = (in_do|_reg_1);
   assign  _net_686 = (in_do|_reg_1);
   assign  _net_687 = (in_do|_reg_1);
   assign  _net_688 = (in_do|_reg_1);
   assign  _net_689 = (in_do|_reg_1);
   assign  _net_690 = (in_do|_reg_1);
   assign  _net_691 = (in_do|_reg_1);
   assign  _net_692 = (in_do|_reg_1);
   assign  _net_693 = (in_do|_reg_1);
   assign  _net_694 = (in_do|_reg_1);
   assign  _net_695 = (in_do|_reg_1);
   assign  _net_696 = (in_do|_reg_1);
   assign  _net_697 = (in_do|_reg_1);
   assign  _net_698 = (in_do|_reg_1);
   assign  _net_699 = (in_do|_reg_1);
   assign  _net_700 = (in_do|_reg_1);
   assign  _net_701 = (in_do|_reg_1);
   assign  _net_702 = (in_do|_reg_1);
   assign  _net_703 = (in_do|_reg_1);
   assign  _net_704 = (in_do|_reg_1);
   assign  _net_705 = (in_do|_reg_1);
   assign  _net_706 = (in_do|_reg_1);
   assign  _net_707 = (in_do|_reg_1);
   assign  _net_708 = (in_do|_reg_1);
   assign  _net_709 = (in_do|_reg_1);
   assign  _net_710 = (in_do|_reg_1);
   assign  _net_711 = (in_do|_reg_1);
   assign  _net_712 = (in_do|_reg_1);
   assign  _net_713 = (in_do|_reg_1);
   assign  _net_714 = (in_do|_reg_1);
   assign  _net_715 = (in_do|_reg_1);
   assign  _net_716 = (in_do|_reg_1);
   assign  _net_717 = (in_do|_reg_1);
   assign  _net_718 = (in_do|_reg_1);
   assign  _net_719 = (in_do|_reg_1);
   assign  _net_720 = (in_do|_reg_1);
   assign  _net_721 = (in_do|_reg_1);
   assign  _net_722 = (in_do|_reg_1);
   assign  _net_723 = (in_do|_reg_1);
   assign  _net_724 = (in_do|_reg_1);
   assign  _net_725 = (in_do|_reg_1);
   assign  _net_726 = (in_do|_reg_1);
   assign  _net_727 = (in_do|_reg_1);
   assign  _net_728 = (in_do|_reg_1);
   assign  _net_729 = (in_do|_reg_1);
   assign  _net_730 = (in_do|_reg_1);
   assign  _net_731 = (in_do|_reg_1);
   assign  _net_732 = (in_do|_reg_1);
   assign  _net_733 = (in_do|_reg_1);
   assign  _net_734 = (in_do|_reg_1);
   assign  _net_735 = (in_do|_reg_1);
   assign  _net_736 = (in_do|_reg_1);
   assign  _net_737 = (in_do|_reg_1);
   assign  _net_738 = (in_do|_reg_1);
   assign  _net_739 = (in_do|_reg_1);
   assign  _net_740 = (in_do|_reg_1);
   assign  _net_741 = (in_do|_reg_1);
   assign  _net_742 = (in_do|_reg_1);
   assign  _net_743 = (in_do|_reg_1);
   assign  _net_744 = (in_do|_reg_1);
   assign  _net_745 = (in_do|_reg_1);
   assign  _net_746 = (in_do|_reg_1);
   assign  _net_747 = (in_do|_reg_1);
   assign  _net_748 = (in_do|_reg_1);
   assign  _net_749 = (in_do|_reg_1);
   assign  _net_750 = (in_do|_reg_1);
   assign  _net_751 = (in_do|_reg_1);
   assign  _net_752 = (in_do|_reg_1);
   assign  _net_753 = (in_do|_reg_1);
   assign  _net_754 = (in_do|_reg_1);
   assign  _net_755 = (in_do|_reg_1);
   assign  _net_756 = (in_do|_reg_1);
   assign  _net_757 = (in_do|_reg_1);
   assign  _net_758 = (in_do|_reg_1);
   assign  _net_759 = (in_do|_reg_1);
   assign  _net_760 = (in_do|_reg_1);
   assign  _net_761 = (in_do|_reg_1);
   assign  _net_762 = (in_do|_reg_1);
   assign  _net_763 = (in_do|_reg_1);
   assign  _net_764 = (in_do|_reg_1);
   assign  _net_765 = (in_do|_reg_1);
   assign  _net_766 = (in_do|_reg_1);
   assign  _net_767 = (in_do|_reg_1);
   assign  _net_768 = (in_do|_reg_1);
   assign  _net_769 = (in_do|_reg_1);
   assign  _net_770 = (in_do|_reg_1);
   assign  _net_771 = (in_do|_reg_1);
   assign  _net_772 = (in_do|_reg_1);
   assign  _net_773 = (in_do|_reg_1);
   assign  _net_774 = (in_do|_reg_1);
   assign  _net_775 = (in_do|_reg_1);
   assign  _net_776 = (in_do|_reg_1);
   assign  _net_777 = (in_do|_reg_1);
   assign  _net_778 = (in_do|_reg_1);
   assign  _net_779 = (in_do|_reg_1);
   assign  _net_780 = (in_do|_reg_1);
   assign  _net_781 = (in_do|_reg_1);
   assign  _net_782 = (in_do|_reg_1);
   assign  _net_783 = (in_do|_reg_1);
   assign  _net_784 = (in_do|_reg_1);
   assign  _net_785 = (in_do|_reg_1);
   assign  _net_786 = (in_do|_reg_1);
   assign  _net_787 = (in_do|_reg_1);
   assign  _net_788 = (in_do|_reg_1);
   assign  _net_789 = (in_do|_reg_1);
   assign  _net_790 = (in_do|_reg_1);
   assign  _net_791 = (in_do|_reg_1);
   assign  _net_792 = (in_do|_reg_1);
   assign  _net_793 = (in_do|_reg_1);
   assign  _net_794 = (in_do|_reg_1);
   assign  _net_795 = (in_do|_reg_1);
   assign  _net_796 = (in_do|_reg_1);
   assign  _net_797 = (in_do|_reg_1);
   assign  _net_798 = (in_do|_reg_1);
   assign  _net_799 = (in_do|_reg_1);
   assign  _net_800 = (in_do|_reg_1);
   assign  _net_801 = (in_do|_reg_1);
   assign  _net_802 = (in_do|_reg_1);
   assign  _net_803 = (in_do|_reg_1);
   assign  _net_804 = (in_do|_reg_1);
   assign  _net_805 = (in_do|_reg_1);
   assign  _net_806 = (in_do|_reg_1);
   assign  _net_807 = (in_do|_reg_1);
   assign  _net_808 = (in_do|_reg_1);
   assign  _net_809 = (in_do|_reg_1);
   assign  _net_810 = (in_do|_reg_1);
   assign  _net_811 = (in_do|_reg_1);
   assign  _net_812 = (in_do|_reg_1);
   assign  _net_813 = (in_do|_reg_1);
   assign  _net_814 = (in_do|_reg_1);
   assign  _net_815 = (in_do|_reg_1);
   assign  _net_816 = (in_do|_reg_1);
   assign  _net_817 = (in_do|_reg_1);
   assign  _net_818 = (in_do|_reg_1);
   assign  _net_819 = (in_do|_reg_1);
   assign  _net_820 = (in_do|_reg_1);
   assign  _net_821 = (in_do|_reg_1);
   assign  _net_822 = (in_do|_reg_1);
   assign  _net_823 = (in_do|_reg_1);
   assign  _net_824 = (in_do|_reg_1);
   assign  _net_825 = (in_do|_reg_1);
   assign  _net_826 = (in_do|_reg_1);
   assign  _net_827 = (in_do|_reg_1);
   assign  _net_828 = (in_do|_reg_1);
   assign  _net_829 = (in_do|_reg_1);
   assign  _net_830 = (in_do|_reg_1);
   assign  _net_831 = (in_do|_reg_1);
   assign  _net_832 = (in_do|_reg_1);
   assign  _net_833 = (in_do|_reg_1);
   assign  _net_834 = (in_do|_reg_1);
   assign  _net_835 = (in_do|_reg_1);
   assign  _net_836 = (in_do|_reg_1);
   assign  _net_837 = (in_do|_reg_1);
   assign  _net_838 = (in_do|_reg_1);
   assign  _net_839 = (in_do|_reg_1);
   assign  _net_840 = (in_do|_reg_1);
   assign  _net_841 = (in_do|_reg_1);
   assign  _net_842 = (in_do|_reg_1);
   assign  _net_843 = (in_do|_reg_1);
   assign  _net_844 = (in_do|_reg_1);
   assign  _net_845 = (in_do|_reg_1);
   assign  _net_846 = (in_do|_reg_1);
   assign  _net_847 = (in_do|_reg_1);
   assign  _net_848 = (in_do|_reg_1);
   assign  _net_849 = (in_do|_reg_1);
   assign  _net_850 = (in_do|_reg_1);
   assign  _net_851 = (in_do|_reg_1);
   assign  _net_852 = (in_do|_reg_1);
   assign  _net_853 = (in_do|_reg_1);
   assign  _net_854 = (in_do|_reg_1);
   assign  _net_855 = (in_do|_reg_1);
   assign  _net_856 = (in_do|_reg_1);
   assign  _net_857 = (in_do|_reg_1);
   assign  _net_858 = (in_do|_reg_1);
   assign  _net_859 = (in_do|_reg_1);
   assign  _net_860 = (in_do|_reg_1);
   assign  _net_861 = (in_do|_reg_1);
   assign  _net_862 = (in_do|_reg_1);
   assign  _net_863 = (in_do|_reg_1);
   assign  _net_864 = (in_do|_reg_1);
   assign  _net_865 = (in_do|_reg_1);
   assign  _net_866 = (in_do|_reg_1);
   assign  _net_867 = (in_do|_reg_1);
   assign  _net_868 = (in_do|_reg_1);
   assign  _net_869 = (in_do|_reg_1);
   assign  _net_870 = (in_do|_reg_1);
   assign  _net_871 = (in_do|_reg_1);
   assign  _net_872 = (in_do|_reg_1);
   assign  _net_873 = (in_do|_reg_1);
   assign  _net_874 = (in_do|_reg_1);
   assign  _net_875 = (in_do|_reg_1);
   assign  _net_876 = (in_do|_reg_1);
   assign  _net_877 = (in_do|_reg_1);
   assign  _net_878 = (in_do|_reg_1);
   assign  _net_879 = (in_do|_reg_1);
   assign  _net_880 = (in_do|_reg_1);
   assign  _net_881 = (in_do|_reg_1);
   assign  _net_882 = (in_do|_reg_1);
   assign  _net_883 = (in_do|_reg_1);
   assign  _net_884 = (in_do|_reg_1);
   assign  _net_885 = (in_do|_reg_1);
   assign  _net_886 = (in_do|_reg_1);
   assign  _net_887 = (in_do|_reg_1);
   assign  _net_888 = (in_do|_reg_1);
   assign  _net_889 = (in_do|_reg_1);
   assign  _net_890 = (in_do|_reg_1);
   assign  _net_891 = (in_do|_reg_1);
   assign  _net_892 = (in_do|_reg_1);
   assign  _net_893 = (in_do|_reg_1);
   assign  _net_894 = (in_do|_reg_1);
   assign  _net_895 = (in_do|_reg_1);
   assign  _net_896 = (in_do|_reg_1);
   assign  _net_897 = (in_do|_reg_1);
   assign  _net_898 = (in_do|_reg_1);
   assign  _net_899 = (in_do|_reg_1);
   assign  _net_900 = (in_do|_reg_1);
   assign  _net_901 = (in_do|_reg_1);
   assign  _net_902 = (in_do|_reg_1);
   assign  _net_903 = (in_do|_reg_1);
   assign  _net_904 = (in_do|_reg_1);
   assign  _net_905 = (in_do|_reg_1);
   assign  _net_906 = (in_do|_reg_1);
   assign  _net_907 = (in_do|_reg_1);
   assign  _net_908 = (in_do|_reg_1);
   assign  _net_909 = (in_do|_reg_1);
   assign  _net_910 = (in_do|_reg_1);
   assign  _net_911 = (in_do|_reg_1);
   assign  _net_912 = (in_do|_reg_1);
   assign  _net_913 = (in_do|_reg_1);
   assign  _net_914 = (in_do|_reg_1);
   assign  _net_915 = (in_do|_reg_1);
   assign  _net_916 = (in_do|_reg_1);
   assign  _net_917 = (in_do|_reg_1);
   assign  _net_918 = (in_do|_reg_1);
   assign  _net_919 = (in_do|_reg_1);
   assign  _net_920 = (in_do|_reg_1);
   assign  _net_921 = (in_do|_reg_1);
   assign  _net_922 = (in_do|_reg_1);
   assign  _net_923 = (in_do|_reg_1);
   assign  _net_924 = (in_do|_reg_1);
   assign  _net_925 = (in_do|_reg_1);
   assign  _net_926 = (in_do|_reg_1);
   assign  _net_927 = (in_do|_reg_1);
   assign  _net_928 = (in_do|_reg_1);
   assign  _net_929 = (in_do|_reg_1);
   assign  _net_930 = (in_do|_reg_1);
   assign  _net_931 = (in_do|_reg_1);
   assign  _net_932 = (in_do|_reg_1);
   assign  _net_933 = (in_do|_reg_1);
   assign  _net_934 = (in_do|_reg_1);
   assign  _net_935 = (in_do|_reg_1);
   assign  _net_936 = (in_do|_reg_1);
   assign  _net_937 = (in_do|_reg_1);
   assign  _net_938 = (in_do|_reg_1);
   assign  _net_939 = (in_do|_reg_1);
   assign  _net_940 = (in_do|_reg_1);
   assign  _net_941 = (in_do|_reg_1);
   assign  _net_942 = (in_do|_reg_1);
   assign  _net_943 = (in_do|_reg_1);
   assign  _net_944 = (in_do|_reg_1);
   assign  _net_945 = (in_do|_reg_1);
   assign  _net_946 = (in_do|_reg_1);
   assign  _net_947 = (in_do|_reg_1);
   assign  _net_948 = (in_do|_reg_1);
   assign  _net_949 = (in_do|_reg_1);
   assign  _net_950 = (in_do|_reg_1);
   assign  _net_951 = (in_do|_reg_1);
   assign  _net_952 = (in_do|_reg_1);
   assign  _net_953 = (in_do|_reg_1);
   assign  _net_954 = (in_do|_reg_1);
   assign  _net_955 = (in_do|_reg_1);
   assign  _net_956 = (in_do|_reg_1);
   assign  _net_957 = (in_do|_reg_1);
   assign  _net_958 = (in_do|_reg_1);
   assign  _net_959 = (in_do|_reg_1);
   assign  _net_960 = (in_do|_reg_1);
   assign  _net_961 = (in_do|_reg_1);
   assign  _net_962 = (in_do|_reg_1);
   assign  _net_963 = (in_do|_reg_1);
   assign  _net_964 = (in_do|_reg_1);
   assign  _net_965 = (in_do|_reg_1);
   assign  _net_966 = (in_do|_reg_1);
   assign  _net_967 = (in_do|_reg_1);
   assign  _net_968 = (in_do|_reg_1);
   assign  _net_969 = (in_do|_reg_1);
   assign  _net_970 = (in_do|_reg_1);
   assign  _net_971 = (in_do|_reg_1);
   assign  _net_972 = (in_do|_reg_1);
   assign  _net_973 = (in_do|_reg_1);
   assign  _net_974 = (in_do|_reg_1);
   assign  _net_975 = (in_do|_reg_1);
   assign  _net_976 = (in_do|_reg_1);
   assign  _net_977 = (in_do|_reg_1);
   assign  _net_978 = (in_do|_reg_1);
   assign  _net_979 = (in_do|_reg_1);
   assign  _net_980 = (in_do|_reg_1);
   assign  _net_981 = (in_do|_reg_1);
   assign  _net_982 = (in_do|_reg_1);
   assign  _net_983 = (in_do|_reg_1);
   assign  _net_984 = (in_do|_reg_1);
   assign  _net_985 = (in_do|_reg_1);
   assign  _net_986 = (in_do|_reg_1);
   assign  _net_987 = (in_do|_reg_1);
   assign  _net_988 = (in_do|_reg_1);
   assign  _net_989 = (in_do|_reg_1);
   assign  _net_990 = (in_do|_reg_1);
   assign  _net_991 = (in_do|_reg_1);
   assign  _net_992 = (in_do|_reg_1);
   assign  _net_993 = (in_do|_reg_1);
   assign  _net_994 = (in_do|_reg_1);
   assign  _net_995 = (in_do|_reg_1);
   assign  _net_996 = (in_do|_reg_1);
   assign  _net_997 = (in_do|_reg_1);
   assign  _net_998 = (in_do|_reg_1);
   assign  _net_999 = (in_do|_reg_1);
   assign  _net_1000 = (in_do|_reg_1);
   assign  _net_1001 = (in_do|_reg_1);
   assign  _net_1002 = (in_do|_reg_1);
   assign  _net_1003 = (in_do|_reg_1);
   assign  _net_1004 = (in_do|_reg_1);
   assign  _net_1005 = (in_do|_reg_1);
   assign  _net_1006 = (in_do|_reg_1);
   assign  _net_1007 = (in_do|_reg_1);
   assign  _net_1008 = (in_do|_reg_1);
   assign  _net_1009 = (in_do|_reg_1);
   assign  _net_1010 = (in_do|_reg_1);
   assign  _net_1011 = (in_do|_reg_1);
   assign  _net_1012 = (in_do|_reg_1);
   assign  _net_1013 = (in_do|_reg_1);
   assign  _net_1014 = (in_do|_reg_1);
   assign  _net_1015 = (in_do|_reg_1);
   assign  _net_1016 = (in_do|_reg_1);
   assign  _net_1017 = (in_do|_reg_1);
   assign  _net_1018 = (in_do|_reg_1);
   assign  _net_1019 = (in_do|_reg_1);
   assign  _net_1020 = (in_do|_reg_1);
   assign  _net_1021 = (in_do|_reg_1);
   assign  _net_1022 = (in_do|_reg_1);
   assign  _net_1023 = (in_do|_reg_1);
   assign  _net_1024 = (in_do|_reg_1);
   assign  _net_1025 = (in_do|_reg_1);
   assign  _net_1026 = (in_do|_reg_1);
   assign  _net_1027 = (in_do|_reg_1);
   assign  _net_1028 = (in_do|_reg_1);
   assign  _net_1029 = (in_do|_reg_1);
   assign  _net_1030 = (in_do|_reg_1);
   assign  _net_1031 = (in_do|_reg_1);
   assign  _net_1032 = (in_do|_reg_1);
   assign  _net_1033 = (in_do|_reg_1);
   assign  _net_1034 = (in_do|_reg_1);
   assign  _net_1035 = (in_do|_reg_1);
   assign  _net_1036 = (in_do|_reg_1);
   assign  _net_1037 = (in_do|_reg_1);
   assign  _net_1038 = (in_do|_reg_1);
   assign  _net_1039 = (in_do|_reg_1);
   assign  _net_1040 = (in_do|_reg_1);
   assign  _net_1041 = (in_do|_reg_1);
   assign  _net_1042 = (in_do|_reg_1);
   assign  _net_1043 = (in_do|_reg_1);
   assign  _net_1044 = (in_do|_reg_1);
   assign  _net_1045 = (in_do|_reg_1);
   assign  _net_1046 = (in_do|_reg_1);
   assign  _net_1047 = (in_do|_reg_1);
   assign  _net_1048 = (in_do|_reg_1);
   assign  _net_1049 = (in_do|_reg_1);
   assign  _net_1050 = (in_do|_reg_1);
   assign  _net_1051 = (in_do|_reg_1);
   assign  _net_1052 = (in_do|_reg_1);
   assign  _net_1053 = (in_do|_reg_1);
   assign  _net_1054 = (in_do|_reg_1);
   assign  _net_1055 = (in_do|_reg_1);
   assign  _net_1056 = (in_do|_reg_1);
   assign  _net_1057 = (in_do|_reg_1);
   assign  _net_1058 = (in_do|_reg_1);
   assign  _net_1059 = (in_do|_reg_1);
   assign  _net_1060 = (in_do|_reg_1);
   assign  _net_1061 = (in_do|_reg_1);
   assign  _net_1062 = (in_do|_reg_1);
   assign  _net_1063 = (in_do|_reg_1);
   assign  _net_1064 = (in_do|_reg_1);
   assign  _net_1065 = (in_do|_reg_1);
   assign  _net_1066 = (in_do|_reg_1);
   assign  _net_1067 = (in_do|_reg_1);
   assign  _net_1068 = (in_do|_reg_1);
   assign  _net_1069 = (in_do|_reg_1);
   assign  _net_1070 = (in_do|_reg_1);
   assign  _net_1071 = (in_do|_reg_1);
   assign  _net_1072 = (in_do|_reg_1);
   assign  _net_1073 = (in_do|_reg_1);
   assign  _net_1074 = (in_do|_reg_1);
   assign  _net_1075 = (in_do|_reg_1);
   assign  _net_1076 = (in_do|_reg_1);
   assign  _net_1077 = (in_do|_reg_1);
   assign  _net_1078 = (in_do|_reg_1);
   assign  _net_1079 = (in_do|_reg_1);
   assign  _net_1080 = (in_do|_reg_1);
   assign  _net_1081 = (in_do|_reg_1);
   assign  _net_1082 = (in_do|_reg_1);
   assign  _net_1083 = (in_do|_reg_1);
   assign  _net_1084 = (in_do|_reg_1);
   assign  _net_1085 = (in_do|_reg_1);
   assign  _net_1086 = (in_do|_reg_1);
   assign  _net_1087 = (in_do|_reg_1);
   assign  _net_1088 = (in_do|_reg_1);
   assign  _net_1089 = (in_do|_reg_1);
   assign  _net_1090 = (in_do|_reg_1);
   assign  _net_1091 = (in_do|_reg_1);
   assign  _net_1092 = (in_do|_reg_1);
   assign  _net_1093 = (in_do|_reg_1);
   assign  _net_1094 = (in_do|_reg_1);
   assign  _net_1095 = (in_do|_reg_1);
   assign  _net_1096 = (in_do|_reg_1);
   assign  _net_1097 = (in_do|_reg_1);
   assign  _net_1098 = (in_do|_reg_1);
   assign  _net_1099 = (in_do|_reg_1);
   assign  _net_1100 = (in_do|_reg_1);
   assign  _net_1101 = (in_do|_reg_1);
   assign  _net_1102 = (in_do|_reg_1);
   assign  _net_1103 = (in_do|_reg_1);
   assign  _net_1104 = (in_do|_reg_1);
   assign  _net_1105 = (in_do|_reg_1);
   assign  _net_1106 = (in_do|_reg_1);
   assign  _net_1107 = (in_do|_reg_1);
   assign  _net_1108 = (in_do|_reg_1);
   assign  _net_1109 = (in_do|_reg_1);
   assign  _net_1110 = (in_do|_reg_1);
   assign  _net_1111 = (in_do|_reg_1);
   assign  _net_1112 = (in_do|_reg_1);
   assign  _net_1113 = (in_do|_reg_1);
   assign  _net_1114 = (in_do|_reg_1);
   assign  _net_1115 = (in_do|_reg_1);
   assign  _net_1116 = (in_do|_reg_1);
   assign  _net_1117 = (in_do|_reg_1);
   assign  _net_1118 = (in_do|_reg_1);
   assign  _net_1119 = (in_do|_reg_1);
   assign  _net_1120 = (in_do|_reg_1);
   assign  _net_1121 = (in_do|_reg_1);
   assign  _net_1122 = (in_do|_reg_1);
   assign  _net_1123 = (in_do|_reg_1);
   assign  _net_1124 = (in_do|_reg_1);
   assign  _net_1125 = (in_do|_reg_1);
   assign  _net_1126 = (in_do|_reg_1);
   assign  _net_1127 = (in_do|_reg_1);
   assign  _net_1128 = (in_do|_reg_1);
   assign  _net_1129 = (in_do|_reg_1);
   assign  _net_1130 = (in_do|_reg_1);
   assign  _net_1131 = (in_do|_reg_1);
   assign  _net_1132 = (in_do|_reg_1);
   assign  _net_1133 = (in_do|_reg_1);
   assign  _net_1134 = (in_do|_reg_1);
   assign  _net_1135 = (in_do|_reg_1);
   assign  _net_1136 = (in_do|_reg_1);
   assign  _net_1137 = (in_do|_reg_1);
   assign  _net_1138 = (in_do|_reg_1);
   assign  _net_1139 = (in_do|_reg_1);
   assign  _net_1140 = (in_do|_reg_1);
   assign  _net_1141 = (in_do|_reg_1);
   assign  _net_1142 = (in_do|_reg_1);
   assign  _net_1143 = (in_do|_reg_1);
   assign  _net_1144 = (in_do|_reg_1);
   assign  _net_1145 = (in_do|_reg_1);
   assign  _net_1146 = (in_do|_reg_1);
   assign  _net_1147 = (in_do|_reg_1);
   assign  _net_1148 = (in_do|_reg_1);
   assign  _net_1149 = (in_do|_reg_1);
   assign  _net_1150 = (in_do|_reg_1);
   assign  _net_1151 = (in_do|_reg_1);
   assign  _net_1152 = (in_do|_reg_1);
   assign  _net_1153 = (in_do|_reg_1);
   assign  _net_1154 = (in_do|_reg_1);
   assign  _net_1155 = (in_do|_reg_1);
   assign  _net_1156 = (in_do|_reg_1);
   assign  _net_1157 = (in_do|_reg_1);
   assign  _net_1158 = (in_do|_reg_1);
   assign  _net_1159 = (in_do|_reg_1);
   assign  _net_1160 = (in_do|_reg_1);
   assign  _net_1161 = (in_do|_reg_1);
   assign  _net_1162 = (in_do|_reg_1);
   assign  _net_1163 = (in_do|_reg_1);
   assign  _net_1164 = (in_do|_reg_1);
   assign  _net_1165 = (in_do|_reg_1);
   assign  _net_1166 = (in_do|_reg_1);
   assign  _net_1167 = (in_do|_reg_1);
   assign  _net_1168 = (in_do|_reg_1);
   assign  _net_1169 = (in_do|_reg_1);
   assign  _net_1170 = (in_do|_reg_1);
   assign  _net_1171 = (in_do|_reg_1);
   assign  _net_1172 = (in_do|_reg_1);
   assign  _net_1173 = (in_do|_reg_1);
   assign  _net_1174 = (in_do|_reg_1);
   assign  _net_1175 = (in_do|_reg_1);
   assign  _net_1176 = (in_do|_reg_1);
   assign  _net_1177 = (in_do|_reg_1);
   assign  _net_1178 = (in_do|_reg_1);
   assign  _net_1179 = (in_do|_reg_1);
   assign  _net_1180 = (in_do|_reg_1);
   assign  _net_1181 = (in_do|_reg_1);
   assign  _net_1182 = (in_do|_reg_1);
   assign  _net_1183 = (in_do|_reg_1);
   assign  _net_1184 = (in_do|_reg_1);
   assign  _net_1185 = (in_do|_reg_1);
   assign  _net_1186 = (in_do|_reg_1);
   assign  _net_1187 = (in_do|_reg_1);
   assign  _net_1188 = (in_do|_reg_1);
   assign  _net_1189 = (in_do|_reg_1);
   assign  _net_1190 = (in_do|_reg_1);
   assign  _net_1191 = (in_do|_reg_1);
   assign  _net_1192 = (in_do|_reg_1);
   assign  _net_1193 = (in_do|_reg_1);
   assign  _net_1194 = (in_do|_reg_1);
   assign  _net_1195 = (in_do|_reg_1);
   assign  _net_1196 = (in_do|_reg_1);
   assign  _net_1197 = (in_do|_reg_1);
   assign  _net_1198 = (in_do|_reg_1);
   assign  _net_1199 = (in_do|_reg_1);
   assign  _net_1200 = (in_do|_reg_1);
   assign  _net_1201 = (in_do|_reg_1);
   assign  _net_1202 = (in_do|_reg_1);
   assign  _net_1203 = (in_do|_reg_1);
   assign  _net_1204 = (in_do|_reg_1);
   assign  _net_1205 = (in_do|_reg_1);
   assign  _net_1206 = (in_do|_reg_1);
   assign  _net_1207 = (in_do|_reg_1);
   assign  _net_1208 = (in_do|_reg_1);
   assign  _net_1209 = (in_do|_reg_1);
   assign  _net_1210 = (in_do|_reg_1);
   assign  _net_1211 = (in_do|_reg_1);
   assign  _net_1212 = (in_do|_reg_1);
   assign  _net_1213 = (in_do|_reg_1);
   assign  _net_1214 = (in_do|_reg_1);
   assign  _net_1215 = (in_do|_reg_1);
   assign  _net_1216 = (in_do|_reg_1);
   assign  _net_1217 = (in_do|_reg_1);
   assign  _net_1218 = (in_do|_reg_1);
   assign  _net_1219 = (in_do|_reg_1);
   assign  _net_1220 = (in_do|_reg_1);
   assign  _net_1221 = (in_do|_reg_1);
   assign  _net_1222 = (in_do|_reg_1);
   assign  _net_1223 = (in_do|_reg_1);
   assign  _net_1224 = (in_do|_reg_1);
   assign  _net_1225 = (in_do|_reg_1);
   assign  _net_1226 = (in_do|_reg_1);
   assign  _net_1227 = (in_do|_reg_1);
   assign  _net_1228 = (in_do|_reg_1);
   assign  _net_1229 = (in_do|_reg_1);
   assign  _net_1230 = (in_do|_reg_1);
   assign  _net_1231 = (in_do|_reg_1);
   assign  _net_1232 = (in_do|_reg_1);
   assign  _net_1233 = (in_do|_reg_1);
   assign  _net_1234 = (in_do|_reg_1);
   assign  _net_1235 = (in_do|_reg_1);
   assign  _net_1236 = (in_do|_reg_1);
   assign  _net_1237 = (in_do|_reg_1);
   assign  _net_1238 = (in_do|_reg_1);
   assign  _net_1239 = (in_do|_reg_1);
   assign  _net_1240 = (in_do|_reg_1);
   assign  _net_1241 = (in_do|_reg_1);
   assign  _net_1242 = (in_do|_reg_1);
   assign  _net_1243 = (in_do|_reg_1);
   assign  _net_1244 = (in_do|_reg_1);
   assign  _net_1245 = (in_do|_reg_1);
   assign  _net_1246 = (in_do|_reg_1);
   assign  _net_1247 = (in_do|_reg_1);
   assign  _net_1248 = (in_do|_reg_1);
   assign  _net_1249 = (in_do|_reg_1);
   assign  _net_1250 = (in_do|_reg_1);
   assign  _net_1251 = (in_do|_reg_1);
   assign  _net_1252 = (in_do|_reg_1);
   assign  _net_1253 = (in_do|_reg_1);
   assign  _net_1254 = (in_do|_reg_1);
   assign  _net_1255 = (in_do|_reg_1);
   assign  _net_1256 = (in_do|_reg_1);
   assign  _net_1257 = (in_do|_reg_1);
   assign  _net_1258 = (in_do|_reg_1);
   assign  _net_1259 = (in_do|_reg_1);
   assign  _net_1260 = (in_do|_reg_1);
   assign  _net_1261 = (in_do|_reg_1);
   assign  _net_1262 = (in_do|_reg_1);
   assign  _net_1263 = (in_do|_reg_1);
   assign  _net_1264 = (in_do|(_reg_0|_reg_1));
   assign  data_out33 = _seach_blockx_data_out;
   assign  data_out34 = _seach_blockx_1_data_out;
   assign  data_out35 = _seach_blockx_2_data_out;
   assign  data_out36 = _seach_blockx_3_data_out;
   assign  data_out37 = _seach_blockx_4_data_out;
   assign  data_out38 = _seach_blockx_5_data_out;
   assign  data_out39 = _seach_blockx_6_data_out;
   assign  data_out40 = _seach_blockx_7_data_out;
   assign  data_out41 = _seach_blockx_8_data_out;
   assign  data_out42 = _seach_blockx_9_data_out;
   assign  data_out43 = _seach_blockx_10_data_out;
   assign  data_out44 = _seach_blockx_11_data_out;
   assign  data_out45 = _seach_blockx_12_data_out;
   assign  data_out46 = _seach_blockx_13_data_out;
   assign  data_out47 = _seach_blockx_14_data_out;
   assign  data_out48 = _seach_blockx_15_data_out;
   assign  data_out49 = _seach_blockx_16_data_out;
   assign  data_out50 = _seach_blockx_17_data_out;
   assign  data_out51 = _seach_blockx_18_data_out;
   assign  data_out52 = _seach_blockx_19_data_out;
   assign  data_out53 = _seach_blockx_20_data_out;
   assign  data_out54 = _seach_blockx_21_data_out;
   assign  data_out55 = _seach_blockx_22_data_out;
   assign  data_out56 = _seach_blockx_23_data_out;
   assign  data_out57 = _seach_blockx_24_data_out;
   assign  data_out58 = _seach_blockx_25_data_out;
   assign  data_out59 = _seach_blockx_26_data_out;
   assign  data_out60 = _seach_blockx_27_data_out;
   assign  data_out61 = _seach_blockx_28_data_out;
   assign  data_out62 = _seach_blockx_29_data_out;
   assign  data_out65 = _seach_blockx_30_data_out;
   assign  data_out66 = _seach_blockx_31_data_out;
   assign  data_out67 = _seach_blockx_32_data_out;
   assign  data_out68 = _seach_blockx_33_data_out;
   assign  data_out69 = _seach_blockx_34_data_out;
   assign  data_out70 = _seach_blockx_35_data_out;
   assign  data_out71 = _seach_blockx_36_data_out;
   assign  data_out72 = _seach_blockx_37_data_out;
   assign  data_out73 = _seach_blockx_38_data_out;
   assign  data_out74 = _seach_blockx_39_data_out;
   assign  data_out75 = _seach_blockx_40_data_out;
   assign  data_out76 = _seach_blockx_41_data_out;
   assign  data_out77 = _seach_blockx_42_data_out;
   assign  data_out78 = _seach_blockx_43_data_out;
   assign  data_out79 = _seach_blockx_44_data_out;
   assign  data_out80 = _seach_blockx_45_data_out;
   assign  data_out81 = _seach_blockx_46_data_out;
   assign  data_out82 = _seach_blockx_47_data_out;
   assign  data_out83 = _seach_blockx_48_data_out;
   assign  data_out84 = _seach_blockx_49_data_out;
   assign  data_out85 = _seach_blockx_50_data_out;
   assign  data_out86 = _seach_blockx_51_data_out;
   assign  data_out87 = _seach_blockx_52_data_out;
   assign  data_out88 = _seach_blockx_53_data_out;
   assign  data_out89 = _seach_blockx_54_data_out;
   assign  data_out90 = _seach_blockx_55_data_out;
   assign  data_out91 = _seach_blockx_56_data_out;
   assign  data_out92 = _seach_blockx_57_data_out;
   assign  data_out93 = _seach_blockx_58_data_out;
   assign  data_out94 = _seach_blockx_59_data_out;
   assign  data_out97 = _seach_blockx_60_data_out;
   assign  data_out98 = _seach_blockx_61_data_out;
   assign  data_out99 = _seach_blockx_62_data_out;
   assign  data_out100 = _seach_blockx_63_data_out;
   assign  data_out101 = _seach_blockx_64_data_out;
   assign  data_out102 = _seach_blockx_65_data_out;
   assign  data_out103 = _seach_blockx_66_data_out;
   assign  data_out104 = _seach_blockx_67_data_out;
   assign  data_out105 = _seach_blockx_68_data_out;
   assign  data_out106 = _seach_blockx_69_data_out;
   assign  data_out107 = _seach_blockx_70_data_out;
   assign  data_out108 = _seach_blockx_71_data_out;
   assign  data_out109 = _seach_blockx_72_data_out;
   assign  data_out110 = _seach_blockx_73_data_out;
   assign  data_out111 = _seach_blockx_74_data_out;
   assign  data_out112 = _seach_blockx_75_data_out;
   assign  data_out113 = _seach_blockx_76_data_out;
   assign  data_out114 = _seach_blockx_77_data_out;
   assign  data_out115 = _seach_blockx_78_data_out;
   assign  data_out116 = _seach_blockx_79_data_out;
   assign  data_out117 = _seach_blockx_80_data_out;
   assign  data_out118 = _seach_blockx_81_data_out;
   assign  data_out119 = _seach_blockx_82_data_out;
   assign  data_out120 = _seach_blockx_83_data_out;
   assign  data_out121 = _seach_blockx_84_data_out;
   assign  data_out122 = _seach_blockx_85_data_out;
   assign  data_out123 = _seach_blockx_86_data_out;
   assign  data_out124 = _seach_blockx_87_data_out;
   assign  data_out125 = _seach_blockx_88_data_out;
   assign  data_out126 = _seach_blockx_89_data_out;
   assign  data_out129 = _seach_blockx_90_data_out;
   assign  data_out130 = _seach_blockx_91_data_out;
   assign  data_out131 = _seach_blockx_92_data_out;
   assign  data_out132 = _seach_blockx_93_data_out;
   assign  data_out133 = _seach_blockx_94_data_out;
   assign  data_out134 = _seach_blockx_95_data_out;
   assign  data_out135 = _seach_blockx_96_data_out;
   assign  data_out136 = _seach_blockx_97_data_out;
   assign  data_out137 = _seach_blockx_98_data_out;
   assign  data_out138 = _seach_blockx_99_data_out;
   assign  data_out139 = _seach_blockx_100_data_out;
   assign  data_out140 = _seach_blockx_101_data_out;
   assign  data_out141 = _seach_blockx_102_data_out;
   assign  data_out142 = _seach_blockx_103_data_out;
   assign  data_out143 = _seach_blockx_104_data_out;
   assign  data_out144 = _seach_blockx_105_data_out;
   assign  data_out145 = _seach_blockx_106_data_out;
   assign  data_out146 = _seach_blockx_107_data_out;
   assign  data_out147 = _seach_blockx_108_data_out;
   assign  data_out148 = _seach_blockx_109_data_out;
   assign  data_out149 = _seach_blockx_110_data_out;
   assign  data_out150 = _seach_blockx_111_data_out;
   assign  data_out151 = _seach_blockx_112_data_out;
   assign  data_out152 = _seach_blockx_113_data_out;
   assign  data_out153 = _seach_blockx_114_data_out;
   assign  data_out154 = _seach_blockx_115_data_out;
   assign  data_out155 = _seach_blockx_116_data_out;
   assign  data_out156 = _seach_blockx_117_data_out;
   assign  data_out157 = _seach_blockx_118_data_out;
   assign  data_out158 = _seach_blockx_119_data_out;
   assign  data_out161 = _seach_blockx_120_data_out;
   assign  data_out162 = _seach_blockx_121_data_out;
   assign  data_out163 = _seach_blockx_122_data_out;
   assign  data_out164 = _seach_blockx_123_data_out;
   assign  data_out165 = _seach_blockx_124_data_out;
   assign  data_out166 = _seach_blockx_125_data_out;
   assign  data_out167 = _seach_blockx_126_data_out;
   assign  data_out168 = _seach_blockx_127_data_out;
   assign  data_out169 = _seach_blockx_128_data_out;
   assign  data_out170 = _seach_blockx_129_data_out;
   assign  data_out171 = _seach_blockx_130_data_out;
   assign  data_out172 = _seach_blockx_131_data_out;
   assign  data_out173 = _seach_blockx_132_data_out;
   assign  data_out174 = _seach_blockx_133_data_out;
   assign  data_out175 = _seach_blockx_134_data_out;
   assign  data_out176 = _seach_blockx_135_data_out;
   assign  data_out177 = _seach_blockx_136_data_out;
   assign  data_out178 = _seach_blockx_137_data_out;
   assign  data_out179 = _seach_blockx_138_data_out;
   assign  data_out180 = _seach_blockx_139_data_out;
   assign  data_out181 = _seach_blockx_140_data_out;
   assign  data_out182 = _seach_blockx_141_data_out;
   assign  data_out183 = _seach_blockx_142_data_out;
   assign  data_out184 = _seach_blockx_143_data_out;
   assign  data_out185 = _seach_blockx_144_data_out;
   assign  data_out186 = _seach_blockx_145_data_out;
   assign  data_out187 = _seach_blockx_146_data_out;
   assign  data_out188 = _seach_blockx_147_data_out;
   assign  data_out189 = _seach_blockx_148_data_out;
   assign  data_out190 = _seach_blockx_149_data_out;
   assign  data_out193 = _seach_blockx_150_data_out;
   assign  data_out194 = _seach_blockx_151_data_out;
   assign  data_out195 = _seach_blockx_152_data_out;
   assign  data_out196 = _seach_blockx_153_data_out;
   assign  data_out197 = _seach_blockx_154_data_out;
   assign  data_out198 = _seach_blockx_155_data_out;
   assign  data_out199 = _seach_blockx_156_data_out;
   assign  data_out200 = _seach_blockx_157_data_out;
   assign  data_out201 = _seach_blockx_158_data_out;
   assign  data_out202 = _seach_blockx_159_data_out;
   assign  data_out203 = _seach_blockx_160_data_out;
   assign  data_out204 = _seach_blockx_161_data_out;
   assign  data_out205 = _seach_blockx_162_data_out;
   assign  data_out206 = _seach_blockx_163_data_out;
   assign  data_out207 = _seach_blockx_164_data_out;
   assign  data_out208 = _seach_blockx_165_data_out;
   assign  data_out209 = _seach_blockx_166_data_out;
   assign  data_out210 = _seach_blockx_167_data_out;
   assign  data_out211 = _seach_blockx_168_data_out;
   assign  data_out212 = _seach_blockx_169_data_out;
   assign  data_out213 = _seach_blockx_170_data_out;
   assign  data_out214 = _seach_blockx_171_data_out;
   assign  data_out215 = _seach_blockx_172_data_out;
   assign  data_out216 = _seach_blockx_173_data_out;
   assign  data_out217 = _seach_blockx_174_data_out;
   assign  data_out218 = _seach_blockx_175_data_out;
   assign  data_out219 = _seach_blockx_176_data_out;
   assign  data_out220 = _seach_blockx_177_data_out;
   assign  data_out221 = _seach_blockx_178_data_out;
   assign  data_out222 = _seach_blockx_179_data_out;
   assign  data_out225 = _seach_blockx_180_data_out;
   assign  data_out226 = _seach_blockx_181_data_out;
   assign  data_out227 = _seach_blockx_182_data_out;
   assign  data_out228 = _seach_blockx_183_data_out;
   assign  data_out229 = _seach_blockx_184_data_out;
   assign  data_out230 = _seach_blockx_185_data_out;
   assign  data_out231 = _seach_blockx_186_data_out;
   assign  data_out232 = _seach_blockx_187_data_out;
   assign  data_out233 = _seach_blockx_188_data_out;
   assign  data_out234 = _seach_blockx_189_data_out;
   assign  data_out235 = _seach_blockx_190_data_out;
   assign  data_out236 = _seach_blockx_191_data_out;
   assign  data_out237 = _seach_blockx_192_data_out;
   assign  data_out238 = _seach_blockx_193_data_out;
   assign  data_out239 = _seach_blockx_194_data_out;
   assign  data_out240 = _seach_blockx_195_data_out;
   assign  data_out241 = _seach_blockx_196_data_out;
   assign  data_out242 = _seach_blockx_197_data_out;
   assign  data_out243 = _seach_blockx_198_data_out;
   assign  data_out244 = _seach_blockx_199_data_out;
   assign  data_out245 = _seach_blockx_200_data_out;
   assign  data_out246 = _seach_blockx_201_data_out;
   assign  data_out247 = _seach_blockx_202_data_out;
   assign  data_out248 = _seach_blockx_203_data_out;
   assign  data_out249 = _seach_blockx_204_data_out;
   assign  data_out250 = _seach_blockx_205_data_out;
   assign  data_out251 = _seach_blockx_206_data_out;
   assign  data_out252 = _seach_blockx_207_data_out;
   assign  data_out253 = _seach_blockx_208_data_out;
   assign  data_out254 = _seach_blockx_209_data_out;
   assign  data_out257 = _seach_blockx_210_data_out;
   assign  data_out258 = _seach_blockx_211_data_out;
   assign  data_out259 = _seach_blockx_212_data_out;
   assign  data_out260 = _seach_blockx_213_data_out;
   assign  data_out261 = _seach_blockx_214_data_out;
   assign  data_out262 = _seach_blockx_215_data_out;
   assign  data_out263 = _seach_blockx_216_data_out;
   assign  data_out264 = _seach_blockx_217_data_out;
   assign  data_out265 = _seach_blockx_218_data_out;
   assign  data_out266 = _seach_blockx_219_data_out;
   assign  data_out267 = _seach_blockx_220_data_out;
   assign  data_out268 = _seach_blockx_221_data_out;
   assign  data_out269 = _seach_blockx_222_data_out;
   assign  data_out270 = _seach_blockx_223_data_out;
   assign  data_out271 = _seach_blockx_224_data_out;
   assign  data_out272 = _seach_blockx_225_data_out;
   assign  data_out273 = _seach_blockx_226_data_out;
   assign  data_out274 = _seach_blockx_227_data_out;
   assign  data_out275 = _seach_blockx_228_data_out;
   assign  data_out276 = _seach_blockx_229_data_out;
   assign  data_out277 = _seach_blockx_230_data_out;
   assign  data_out278 = _seach_blockx_231_data_out;
   assign  data_out279 = _seach_blockx_232_data_out;
   assign  data_out280 = _seach_blockx_233_data_out;
   assign  data_out281 = _seach_blockx_234_data_out;
   assign  data_out282 = _seach_blockx_235_data_out;
   assign  data_out283 = _seach_blockx_236_data_out;
   assign  data_out284 = _seach_blockx_237_data_out;
   assign  data_out285 = _seach_blockx_238_data_out;
   assign  data_out286 = _seach_blockx_239_data_out;
   assign  data_out289 = _seach_blockx_240_data_out;
   assign  data_out290 = _seach_blockx_241_data_out;
   assign  data_out291 = _seach_blockx_242_data_out;
   assign  data_out292 = _seach_blockx_243_data_out;
   assign  data_out293 = _seach_blockx_244_data_out;
   assign  data_out294 = _seach_blockx_245_data_out;
   assign  data_out295 = _seach_blockx_246_data_out;
   assign  data_out296 = _seach_blockx_247_data_out;
   assign  data_out297 = _seach_blockx_248_data_out;
   assign  data_out298 = _seach_blockx_249_data_out;
   assign  data_out299 = _seach_blockx_250_data_out;
   assign  data_out300 = _seach_blockx_251_data_out;
   assign  data_out301 = _seach_blockx_252_data_out;
   assign  data_out302 = _seach_blockx_253_data_out;
   assign  data_out303 = _seach_blockx_254_data_out;
   assign  data_out304 = _seach_blockx_255_data_out;
   assign  data_out305 = _seach_blockx_256_data_out;
   assign  data_out306 = _seach_blockx_257_data_out;
   assign  data_out307 = _seach_blockx_258_data_out;
   assign  data_out308 = _seach_blockx_259_data_out;
   assign  data_out309 = _seach_blockx_260_data_out;
   assign  data_out310 = _seach_blockx_261_data_out;
   assign  data_out311 = _seach_blockx_262_data_out;
   assign  data_out312 = _seach_blockx_263_data_out;
   assign  data_out313 = _seach_blockx_264_data_out;
   assign  data_out314 = _seach_blockx_265_data_out;
   assign  data_out315 = _seach_blockx_266_data_out;
   assign  data_out316 = _seach_blockx_267_data_out;
   assign  data_out317 = _seach_blockx_268_data_out;
   assign  data_out318 = _seach_blockx_269_data_out;
   assign  data_out321 = _seach_blockx_270_data_out;
   assign  data_out322 = _seach_blockx_271_data_out;
   assign  data_out323 = _seach_blockx_272_data_out;
   assign  data_out324 = _seach_blockx_273_data_out;
   assign  data_out325 = _seach_blockx_274_data_out;
   assign  data_out326 = _seach_blockx_275_data_out;
   assign  data_out327 = _seach_blockx_276_data_out;
   assign  data_out328 = _seach_blockx_277_data_out;
   assign  data_out329 = _seach_blockx_278_data_out;
   assign  data_out330 = _seach_blockx_279_data_out;
   assign  data_out331 = _seach_blockx_280_data_out;
   assign  data_out332 = _seach_blockx_281_data_out;
   assign  data_out333 = _seach_blockx_282_data_out;
   assign  data_out334 = _seach_blockx_283_data_out;
   assign  data_out335 = _seach_blockx_284_data_out;
   assign  data_out336 = _seach_blockx_285_data_out;
   assign  data_out337 = _seach_blockx_286_data_out;
   assign  data_out338 = _seach_blockx_287_data_out;
   assign  data_out339 = _seach_blockx_288_data_out;
   assign  data_out340 = _seach_blockx_289_data_out;
   assign  data_out341 = _seach_blockx_290_data_out;
   assign  data_out342 = _seach_blockx_291_data_out;
   assign  data_out343 = _seach_blockx_292_data_out;
   assign  data_out344 = _seach_blockx_293_data_out;
   assign  data_out345 = _seach_blockx_294_data_out;
   assign  data_out346 = _seach_blockx_295_data_out;
   assign  data_out347 = _seach_blockx_296_data_out;
   assign  data_out348 = _seach_blockx_297_data_out;
   assign  data_out349 = _seach_blockx_298_data_out;
   assign  data_out350 = _seach_blockx_299_data_out;
   assign  data_out353 = _seach_blockx_300_data_out;
   assign  data_out354 = _seach_blockx_301_data_out;
   assign  data_out355 = _seach_blockx_302_data_out;
   assign  data_out356 = _seach_blockx_303_data_out;
   assign  data_out357 = _seach_blockx_304_data_out;
   assign  data_out358 = _seach_blockx_305_data_out;
   assign  data_out359 = _seach_blockx_306_data_out;
   assign  data_out360 = _seach_blockx_307_data_out;
   assign  data_out361 = _seach_blockx_308_data_out;
   assign  data_out362 = _seach_blockx_309_data_out;
   assign  data_out363 = _seach_blockx_310_data_out;
   assign  data_out364 = _seach_blockx_311_data_out;
   assign  data_out365 = _seach_blockx_312_data_out;
   assign  data_out366 = _seach_blockx_313_data_out;
   assign  data_out367 = _seach_blockx_314_data_out;
   assign  data_out368 = _seach_blockx_315_data_out;
   assign  data_out369 = _seach_blockx_316_data_out;
   assign  data_out370 = _seach_blockx_317_data_out;
   assign  data_out371 = _seach_blockx_318_data_out;
   assign  data_out372 = _seach_blockx_319_data_out;
   assign  data_out373 = _seach_blockx_320_data_out;
   assign  data_out374 = _seach_blockx_321_data_out;
   assign  data_out375 = _seach_blockx_322_data_out;
   assign  data_out376 = _seach_blockx_323_data_out;
   assign  data_out377 = _seach_blockx_324_data_out;
   assign  data_out378 = _seach_blockx_325_data_out;
   assign  data_out379 = _seach_blockx_326_data_out;
   assign  data_out380 = _seach_blockx_327_data_out;
   assign  data_out381 = _seach_blockx_328_data_out;
   assign  data_out382 = _seach_blockx_329_data_out;
   assign  data_out385 = _seach_blockx_330_data_out;
   assign  data_out386 = _seach_blockx_331_data_out;
   assign  data_out387 = _seach_blockx_332_data_out;
   assign  data_out388 = _seach_blockx_333_data_out;
   assign  data_out389 = _seach_blockx_334_data_out;
   assign  data_out390 = _seach_blockx_335_data_out;
   assign  data_out391 = _seach_blockx_336_data_out;
   assign  data_out392 = _seach_blockx_337_data_out;
   assign  data_out393 = _seach_blockx_338_data_out;
   assign  data_out394 = _seach_blockx_339_data_out;
   assign  data_out395 = _seach_blockx_340_data_out;
   assign  data_out396 = _seach_blockx_341_data_out;
   assign  data_out397 = _seach_blockx_342_data_out;
   assign  data_out398 = _seach_blockx_343_data_out;
   assign  data_out399 = _seach_blockx_344_data_out;
   assign  data_out400 = _seach_blockx_345_data_out;
   assign  data_out401 = _seach_blockx_346_data_out;
   assign  data_out402 = _seach_blockx_347_data_out;
   assign  data_out403 = _seach_blockx_348_data_out;
   assign  data_out404 = _seach_blockx_349_data_out;
   assign  data_out405 = _seach_blockx_350_data_out;
   assign  data_out406 = _seach_blockx_351_data_out;
   assign  data_out407 = _seach_blockx_352_data_out;
   assign  data_out408 = _seach_blockx_353_data_out;
   assign  data_out409 = _seach_blockx_354_data_out;
   assign  data_out410 = _seach_blockx_355_data_out;
   assign  data_out411 = _seach_blockx_356_data_out;
   assign  data_out412 = _seach_blockx_357_data_out;
   assign  data_out413 = _seach_blockx_358_data_out;
   assign  data_out414 = _seach_blockx_359_data_out;
   assign  data_out417 = _seach_blockx_360_data_out;
   assign  data_out418 = _seach_blockx_361_data_out;
   assign  data_out419 = _seach_blockx_362_data_out;
   assign  data_out420 = _seach_blockx_363_data_out;
   assign  data_out421 = _seach_blockx_364_data_out;
   assign  data_out422 = _seach_blockx_365_data_out;
   assign  data_out423 = _seach_blockx_366_data_out;
   assign  data_out424 = _seach_blockx_367_data_out;
   assign  data_out425 = _seach_blockx_368_data_out;
   assign  data_out426 = _seach_blockx_369_data_out;
   assign  data_out427 = _seach_blockx_370_data_out;
   assign  data_out428 = _seach_blockx_371_data_out;
   assign  data_out429 = _seach_blockx_372_data_out;
   assign  data_out430 = _seach_blockx_373_data_out;
   assign  data_out431 = _seach_blockx_374_data_out;
   assign  data_out432 = _seach_blockx_375_data_out;
   assign  data_out433 = _seach_blockx_376_data_out;
   assign  data_out434 = _seach_blockx_377_data_out;
   assign  data_out435 = _seach_blockx_378_data_out;
   assign  data_out436 = _seach_blockx_379_data_out;
   assign  data_out437 = _seach_blockx_380_data_out;
   assign  data_out438 = _seach_blockx_381_data_out;
   assign  data_out439 = _seach_blockx_382_data_out;
   assign  data_out440 = _seach_blockx_383_data_out;
   assign  data_out441 = _seach_blockx_384_data_out;
   assign  data_out442 = _seach_blockx_385_data_out;
   assign  data_out443 = _seach_blockx_386_data_out;
   assign  data_out444 = _seach_blockx_387_data_out;
   assign  data_out445 = _seach_blockx_388_data_out;
   assign  data_out446 = _seach_blockx_389_data_out;
   assign  data_out449 = _seach_blockx_390_data_out;
   assign  data_out450 = _seach_blockx_391_data_out;
   assign  data_out451 = _seach_blockx_392_data_out;
   assign  data_out452 = _seach_blockx_393_data_out;
   assign  data_out453 = _seach_blockx_394_data_out;
   assign  data_out454 = _seach_blockx_395_data_out;
   assign  data_out455 = _seach_blockx_396_data_out;
   assign  data_out456 = _seach_blockx_397_data_out;
   assign  data_out457 = _seach_blockx_398_data_out;
   assign  data_out458 = _seach_blockx_399_data_out;
   assign  data_out459 = _seach_blockx_400_data_out;
   assign  data_out460 = _seach_blockx_401_data_out;
   assign  data_out461 = _seach_blockx_402_data_out;
   assign  data_out462 = _seach_blockx_403_data_out;
   assign  data_out463 = _seach_blockx_404_data_out;
   assign  data_out464 = _seach_blockx_405_data_out;
   assign  data_out465 = _seach_blockx_406_data_out;
   assign  data_out466 = _seach_blockx_407_data_out;
   assign  data_out467 = _seach_blockx_408_data_out;
   assign  data_out468 = _seach_blockx_409_data_out;
   assign  data_out469 = _seach_blockx_410_data_out;
   assign  data_out470 = _seach_blockx_411_data_out;
   assign  data_out471 = _seach_blockx_412_data_out;
   assign  data_out472 = _seach_blockx_413_data_out;
   assign  data_out473 = _seach_blockx_414_data_out;
   assign  data_out474 = _seach_blockx_415_data_out;
   assign  data_out475 = _seach_blockx_416_data_out;
   assign  data_out476 = _seach_blockx_417_data_out;
   assign  data_out477 = _seach_blockx_418_data_out;
   assign  data_out478 = _seach_blockx_419_data_out;
   assign  startplot = startplot_reg;
   assign  goalplot = goalplot_reg;
   assign  out_do = _reg_0;
   assign  out_data = 1'b1;
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     startplot_reg <= 10'b0000000000;
else if ((_net_1262)) 
      startplot_reg <= (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_seach_blockx_start|_seach_blockx_1_start)|_seach_blockx_2_start)|_seach_blockx_3_start)|_seach_blockx_4_start)|_seach_blockx_5_start)|_seach_blockx_6_start)|_seach_blockx_7_start)|_seach_blockx_8_start)|_seach_blockx_9_start)|_seach_blockx_10_start)|_seach_blockx_11_start)|_seach_blockx_12_start)|_seach_blockx_13_start)|_seach_blockx_14_start)|_seach_blockx_15_start)|_seach_blockx_16_start)|_seach_blockx_17_start)|_seach_blockx_18_start)|_seach_blockx_19_start)|_seach_blockx_20_start)|_seach_blockx_21_start)|_seach_blockx_22_start)|_seach_blockx_23_start)|_seach_blockx_24_start)|_seach_blockx_25_start)|_seach_blockx_26_start)|_seach_blockx_27_start)|_seach_blockx_28_start)|_seach_blockx_29_start)|_seach_blockx_30_start)|_seach_blockx_31_start)|_seach_blockx_32_start)|_seach_blockx_33_start)|_seach_blockx_34_start)|_seach_blockx_35_start)|_seach_blockx_36_start)|_seach_blockx_37_start)|_seach_blockx_38_start)|_seach_blockx_39_start)|_seach_blockx_40_start)|_seach_blockx_41_start)|_seach_blockx_42_start)|_seach_blockx_43_start)|_seach_blockx_44_start)|_seach_blockx_45_start)|_seach_blockx_46_start)|_seach_blockx_47_start)|_seach_blockx_48_start)|_seach_blockx_49_start)|_seach_blockx_50_start)|_seach_blockx_51_start)|_seach_blockx_52_start)|_seach_blockx_53_start)|_seach_blockx_54_start)|_seach_blockx_55_start)|_seach_blockx_56_start)|_seach_blockx_57_start)|_seach_blockx_58_start)|_seach_blockx_59_start)|_seach_blockx_60_start)|_seach_blockx_61_start)|_seach_blockx_62_start)|_seach_blockx_63_start)|_seach_blockx_64_start)|_seach_blockx_65_start)|_seach_blockx_66_start)|_seach_blockx_67_start)|_seach_blockx_68_start)|_seach_blockx_69_start)|_seach_blockx_70_start)|_seach_blockx_71_start)|_seach_blockx_72_start)|_seach_blockx_73_start)|_seach_blockx_74_start)|_seach_blockx_75_start)|_seach_blockx_76_start)|_seach_blockx_77_start)|_seach_blockx_78_start)|_seach_blockx_79_start)|_seach_blockx_80_start)|_seach_blockx_81_start)|_seach_blockx_82_start)|_seach_blockx_83_start)|_seach_blockx_84_start)|_seach_blockx_85_start)|_seach_blockx_86_start)|_seach_blockx_87_start)|_seach_blockx_88_start)|_seach_blockx_89_start)|_seach_blockx_90_start)|_seach_blockx_91_start)|_seach_blockx_92_start)|_seach_blockx_93_start)|_seach_blockx_94_start)|_seach_blockx_95_start)|_seach_blockx_96_start)|_seach_blockx_97_start)|_seach_blockx_98_start)|_seach_blockx_99_start)|_seach_blockx_100_start)|_seach_blockx_101_start)|_seach_blockx_102_start)|_seach_blockx_103_start)|_seach_blockx_104_start)|_seach_blockx_105_start)|_seach_blockx_106_start)|_seach_blockx_107_start)|_seach_blockx_108_start)|_seach_blockx_109_start)|_seach_blockx_110_start)|_seach_blockx_111_start)|_seach_blockx_112_start)|_seach_blockx_113_start)|_seach_blockx_114_start)|_seach_blockx_115_start)|_seach_blockx_116_start)|_seach_blockx_117_start)|_seach_blockx_118_start)|_seach_blockx_119_start)|_seach_blockx_120_start)|_seach_blockx_121_start)|_seach_blockx_122_start)|_seach_blockx_123_start)|_seach_blockx_124_start)|_seach_blockx_125_start)|_seach_blockx_126_start)|_seach_blockx_127_start)|_seach_blockx_128_start)|_seach_blockx_129_start)|_seach_blockx_130_start)|_seach_blockx_131_start)|_seach_blockx_132_start)|_seach_blockx_133_start)|_seach_blockx_134_start)|_seach_blockx_135_start)|_seach_blockx_136_start)|_seach_blockx_137_start)|_seach_blockx_138_start)|_seach_blockx_139_start)|_seach_blockx_140_start)|_seach_blockx_141_start)|_seach_blockx_142_start)|_seach_blockx_143_start)|_seach_blockx_144_start)|_seach_blockx_145_start)|_seach_blockx_146_start)|_seach_blockx_147_start)|_seach_blockx_148_start)|_seach_blockx_149_start)|_seach_blockx_150_start)|_seach_blockx_151_start)|_seach_blockx_152_start)|_seach_blockx_153_start)|_seach_blockx_154_start)|_seach_blockx_155_start)|_seach_blockx_156_start)|_seach_blockx_157_start)|_seach_blockx_158_start)|_seach_blockx_159_start)|_seach_blockx_160_start)|_seach_blockx_161_start)|_seach_blockx_162_start)|_seach_blockx_163_start)|_seach_blockx_164_start)|_seach_blockx_165_start)|_seach_blockx_166_start)|_seach_blockx_167_start)|_seach_blockx_168_start)|_seach_blockx_169_start)|_seach_blockx_170_start)|_seach_blockx_171_start)|_seach_blockx_172_start)|_seach_blockx_173_start)|_seach_blockx_174_start)|_seach_blockx_175_start)|_seach_blockx_176_start)|_seach_blockx_177_start)|_seach_blockx_178_start)|_seach_blockx_179_start)|_seach_blockx_180_start)|_seach_blockx_181_start)|_seach_blockx_182_start)|_seach_blockx_183_start)|_seach_blockx_184_start)|_seach_blockx_185_start)|_seach_blockx_186_start)|_seach_blockx_187_start)|_seach_blockx_188_start)|_seach_blockx_189_start)|_seach_blockx_190_start)|_seach_blockx_191_start)|_seach_blockx_192_start)|_seach_blockx_193_start)|_seach_blockx_194_start)|_seach_blockx_195_start)|_seach_blockx_196_start)|_seach_blockx_197_start)|_seach_blockx_198_start)|_seach_blockx_199_start)|_seach_blockx_200_start)|_seach_blockx_201_start)|_seach_blockx_202_start)|_seach_blockx_203_start)|_seach_blockx_204_start)|_seach_blockx_205_start)|_seach_blockx_206_start)|_seach_blockx_207_start)|_seach_blockx_208_start)|_seach_blockx_209_start)|_seach_blockx_210_start)|_seach_blockx_211_start)|_seach_blockx_212_start)|_seach_blockx_213_start)|_seach_blockx_214_start)|_seach_blockx_215_start)|_seach_blockx_216_start)|_seach_blockx_217_start)|_seach_blockx_218_start)|_seach_blockx_219_start)|_seach_blockx_220_start)|_seach_blockx_221_start)|_seach_blockx_222_start)|_seach_blockx_223_start)|_seach_blockx_224_start)|_seach_blockx_225_start)|_seach_blockx_226_start)|_seach_blockx_227_start)|_seach_blockx_228_start)|_seach_blockx_229_start)|_seach_blockx_230_start)|_seach_blockx_231_start)|_seach_blockx_232_start)|_seach_blockx_233_start)|_seach_blockx_234_start)|_seach_blockx_235_start)|_seach_blockx_236_start)|_seach_blockx_237_start)|_seach_blockx_238_start)|_seach_blockx_239_start)|_seach_blockx_240_start)|_seach_blockx_241_start)|_seach_blockx_242_start)|_seach_blockx_243_start)|_seach_blockx_244_start)|_seach_blockx_245_start)|_seach_blockx_246_start)|_seach_blockx_247_start)|_seach_blockx_248_start)|_seach_blockx_249_start)|_seach_blockx_250_start)|_seach_blockx_251_start)|_seach_blockx_252_start)|_seach_blockx_253_start)|_seach_blockx_254_start)|_seach_blockx_255_start)|_seach_blockx_256_start)|_seach_blockx_257_start)|_seach_blockx_258_start)|_seach_blockx_259_start)|_seach_blockx_260_start)|_seach_blockx_261_start)|_seach_blockx_262_start)|_seach_blockx_263_start)|_seach_blockx_264_start)|_seach_blockx_265_start)|_seach_blockx_266_start)|_seach_blockx_267_start)|_seach_blockx_268_start)|_seach_blockx_269_start)|_seach_blockx_270_start)|_seach_blockx_271_start)|_seach_blockx_272_start)|_seach_blockx_273_start)|_seach_blockx_274_start)|_seach_blockx_275_start)|_seach_blockx_276_start)|_seach_blockx_277_start)|_seach_blockx_278_start)|_seach_blockx_279_start)|_seach_blockx_280_start)|_seach_blockx_281_start)|_seach_blockx_282_start)|_seach_blockx_283_start)|_seach_blockx_284_start)|_seach_blockx_285_start)|_seach_blockx_286_start)|_seach_blockx_287_start)|_seach_blockx_288_start)|_seach_blockx_289_start)|_seach_blockx_290_start)|_seach_blockx_291_start)|_seach_blockx_292_start)|_seach_blockx_293_start)|_seach_blockx_294_start)|_seach_blockx_295_start)|_seach_blockx_296_start)|_seach_blockx_297_start)|_seach_blockx_298_start)|_seach_blockx_299_start)|_seach_blockx_300_start)|_seach_blockx_301_start)|_seach_blockx_302_start)|_seach_blockx_303_start)|_seach_blockx_304_start)|_seach_blockx_305_start)|_seach_blockx_306_start)|_seach_blockx_307_start)|_seach_blockx_308_start)|_seach_blockx_309_start)|_seach_blockx_310_start)|_seach_blockx_311_start)|_seach_blockx_312_start)|_seach_blockx_313_start)|_seach_blockx_314_start)|_seach_blockx_315_start)|_seach_blockx_316_start)|_seach_blockx_317_start)|_seach_blockx_318_start)|_seach_blockx_319_start)|_seach_blockx_320_start)|_seach_blockx_321_start)|_seach_blockx_322_start)|_seach_blockx_323_start)|_seach_blockx_324_start)|_seach_blockx_325_start)|_seach_blockx_326_start)|_seach_blockx_327_start)|_seach_blockx_328_start)|_seach_blockx_329_start)|_seach_blockx_330_start)|_seach_blockx_331_start)|_seach_blockx_332_start)|_seach_blockx_333_start)|_seach_blockx_334_start)|_seach_blockx_335_start)|_seach_blockx_336_start)|_seach_blockx_337_start)|_seach_blockx_338_start)|_seach_blockx_339_start)|_seach_blockx_340_start)|_seach_blockx_341_start)|_seach_blockx_342_start)|_seach_blockx_343_start)|_seach_blockx_344_start)|_seach_blockx_345_start)|_seach_blockx_346_start)|_seach_blockx_347_start)|_seach_blockx_348_start)|_seach_blockx_349_start)|_seach_blockx_350_start)|_seach_blockx_351_start)|_seach_blockx_352_start)|_seach_blockx_353_start)|_seach_blockx_354_start)|_seach_blockx_355_start)|_seach_blockx_356_start)|_seach_blockx_357_start)|_seach_blockx_358_start)|_seach_blockx_359_start)|_seach_blockx_360_start)|_seach_blockx_361_start)|_seach_blockx_362_start)|_seach_blockx_363_start)|_seach_blockx_364_start)|_seach_blockx_365_start)|_seach_blockx_366_start)|_seach_blockx_367_start)|_seach_blockx_368_start)|_seach_blockx_369_start)|_seach_blockx_370_start)|_seach_blockx_371_start)|_seach_blockx_372_start)|_seach_blockx_373_start)|_seach_blockx_374_start)|_seach_blockx_375_start)|_seach_blockx_376_start)|_seach_blockx_377_start)|_seach_blockx_378_start)|_seach_blockx_379_start)|_seach_blockx_380_start)|_seach_blockx_381_start)|_seach_blockx_382_start)|_seach_blockx_383_start)|_seach_blockx_384_start)|_seach_blockx_385_start)|_seach_blockx_386_start)|_seach_blockx_387_start)|_seach_blockx_388_start)|_seach_blockx_389_start)|_seach_blockx_390_start)|_seach_blockx_391_start)|_seach_blockx_392_start)|_seach_blockx_393_start)|_seach_blockx_394_start)|_seach_blockx_395_start)|_seach_blockx_396_start)|_seach_blockx_397_start)|_seach_blockx_398_start)|_seach_blockx_399_start)|_seach_blockx_400_start)|_seach_blockx_401_start)|_seach_blockx_402_start)|_seach_blockx_403_start)|_seach_blockx_404_start)|_seach_blockx_405_start)|_seach_blockx_406_start)|_seach_blockx_407_start)|_seach_blockx_408_start)|_seach_blockx_409_start)|_seach_blockx_410_start)|_seach_blockx_411_start)|_seach_blockx_412_start)|_seach_blockx_413_start)|_seach_blockx_414_start)|_seach_blockx_415_start)|_seach_blockx_416_start)|_seach_blockx_417_start)|_seach_blockx_418_start)|_seach_blockx_419_start);
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     goalplot_reg <= 10'b0000000000;
else if ((_net_1263)) 
      goalplot_reg <= (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_seach_blockx_goal|_seach_blockx_1_goal)|_seach_blockx_2_goal)|_seach_blockx_3_goal)|_seach_blockx_4_goal)|_seach_blockx_5_goal)|_seach_blockx_6_goal)|_seach_blockx_7_goal)|_seach_blockx_8_goal)|_seach_blockx_9_goal)|_seach_blockx_10_goal)|_seach_blockx_11_goal)|_seach_blockx_12_goal)|_seach_blockx_13_goal)|_seach_blockx_14_goal)|_seach_blockx_15_goal)|_seach_blockx_16_goal)|_seach_blockx_17_goal)|_seach_blockx_18_goal)|_seach_blockx_19_goal)|_seach_blockx_20_goal)|_seach_blockx_21_goal)|_seach_blockx_22_goal)|_seach_blockx_23_goal)|_seach_blockx_24_goal)|_seach_blockx_25_goal)|_seach_blockx_26_goal)|_seach_blockx_27_goal)|_seach_blockx_28_goal)|_seach_blockx_29_goal)|_seach_blockx_30_goal)|_seach_blockx_31_goal)|_seach_blockx_32_goal)|_seach_blockx_33_goal)|_seach_blockx_34_goal)|_seach_blockx_35_goal)|_seach_blockx_36_goal)|_seach_blockx_37_goal)|_seach_blockx_38_goal)|_seach_blockx_39_goal)|_seach_blockx_40_goal)|_seach_blockx_41_goal)|_seach_blockx_42_goal)|_seach_blockx_43_goal)|_seach_blockx_44_goal)|_seach_blockx_45_goal)|_seach_blockx_46_goal)|_seach_blockx_47_goal)|_seach_blockx_48_goal)|_seach_blockx_49_goal)|_seach_blockx_50_goal)|_seach_blockx_51_goal)|_seach_blockx_52_goal)|_seach_blockx_53_goal)|_seach_blockx_54_goal)|_seach_blockx_55_goal)|_seach_blockx_56_goal)|_seach_blockx_57_goal)|_seach_blockx_58_goal)|_seach_blockx_59_goal)|_seach_blockx_60_goal)|_seach_blockx_61_goal)|_seach_blockx_62_goal)|_seach_blockx_63_goal)|_seach_blockx_64_goal)|_seach_blockx_65_goal)|_seach_blockx_66_goal)|_seach_blockx_67_goal)|_seach_blockx_68_goal)|_seach_blockx_69_goal)|_seach_blockx_70_goal)|_seach_blockx_71_goal)|_seach_blockx_72_goal)|_seach_blockx_73_goal)|_seach_blockx_74_goal)|_seach_blockx_75_goal)|_seach_blockx_76_goal)|_seach_blockx_77_goal)|_seach_blockx_78_goal)|_seach_blockx_79_goal)|_seach_blockx_80_goal)|_seach_blockx_81_goal)|_seach_blockx_82_goal)|_seach_blockx_83_goal)|_seach_blockx_84_goal)|_seach_blockx_85_goal)|_seach_blockx_86_goal)|_seach_blockx_87_goal)|_seach_blockx_88_goal)|_seach_blockx_89_goal)|_seach_blockx_90_goal)|_seach_blockx_91_goal)|_seach_blockx_92_goal)|_seach_blockx_93_goal)|_seach_blockx_94_goal)|_seach_blockx_95_goal)|_seach_blockx_96_goal)|_seach_blockx_97_goal)|_seach_blockx_98_goal)|_seach_blockx_99_goal)|_seach_blockx_100_goal)|_seach_blockx_101_goal)|_seach_blockx_102_goal)|_seach_blockx_103_goal)|_seach_blockx_104_goal)|_seach_blockx_105_goal)|_seach_blockx_106_goal)|_seach_blockx_107_goal)|_seach_blockx_108_goal)|_seach_blockx_109_goal)|_seach_blockx_110_goal)|_seach_blockx_111_goal)|_seach_blockx_112_goal)|_seach_blockx_113_goal)|_seach_blockx_114_goal)|_seach_blockx_115_goal)|_seach_blockx_116_goal)|_seach_blockx_117_goal)|_seach_blockx_118_goal)|_seach_blockx_119_goal)|_seach_blockx_120_goal)|_seach_blockx_121_goal)|_seach_blockx_122_goal)|_seach_blockx_123_goal)|_seach_blockx_124_goal)|_seach_blockx_125_goal)|_seach_blockx_126_goal)|_seach_blockx_127_goal)|_seach_blockx_128_goal)|_seach_blockx_129_goal)|_seach_blockx_130_goal)|_seach_blockx_131_goal)|_seach_blockx_132_goal)|_seach_blockx_133_goal)|_seach_blockx_134_goal)|_seach_blockx_135_goal)|_seach_blockx_136_goal)|_seach_blockx_137_goal)|_seach_blockx_138_goal)|_seach_blockx_139_goal)|_seach_blockx_140_goal)|_seach_blockx_141_goal)|_seach_blockx_142_goal)|_seach_blockx_143_goal)|_seach_blockx_144_goal)|_seach_blockx_145_goal)|_seach_blockx_146_goal)|_seach_blockx_147_goal)|_seach_blockx_148_goal)|_seach_blockx_149_goal)|_seach_blockx_150_goal)|_seach_blockx_151_goal)|_seach_blockx_152_goal)|_seach_blockx_153_goal)|_seach_blockx_154_goal)|_seach_blockx_155_goal)|_seach_blockx_156_goal)|_seach_blockx_157_goal)|_seach_blockx_158_goal)|_seach_blockx_159_goal)|_seach_blockx_160_goal)|_seach_blockx_161_goal)|_seach_blockx_162_goal)|_seach_blockx_163_goal)|_seach_blockx_164_goal)|_seach_blockx_165_goal)|_seach_blockx_166_goal)|_seach_blockx_167_goal)|_seach_blockx_168_goal)|_seach_blockx_169_goal)|_seach_blockx_170_goal)|_seach_blockx_171_goal)|_seach_blockx_172_goal)|_seach_blockx_173_goal)|_seach_blockx_174_goal)|_seach_blockx_175_goal)|_seach_blockx_176_goal)|_seach_blockx_177_goal)|_seach_blockx_178_goal)|_seach_blockx_179_goal)|_seach_blockx_180_goal)|_seach_blockx_181_goal)|_seach_blockx_182_goal)|_seach_blockx_183_goal)|_seach_blockx_184_goal)|_seach_blockx_185_goal)|_seach_blockx_186_goal)|_seach_blockx_187_goal)|_seach_blockx_188_goal)|_seach_blockx_189_goal)|_seach_blockx_190_goal)|_seach_blockx_191_goal)|_seach_blockx_192_goal)|_seach_blockx_193_goal)|_seach_blockx_194_goal)|_seach_blockx_195_goal)|_seach_blockx_196_goal)|_seach_blockx_197_goal)|_seach_blockx_198_goal)|_seach_blockx_199_goal)|_seach_blockx_200_goal)|_seach_blockx_201_goal)|_seach_blockx_202_goal)|_seach_blockx_203_goal)|_seach_blockx_204_goal)|_seach_blockx_205_goal)|_seach_blockx_206_goal)|_seach_blockx_207_goal)|_seach_blockx_208_goal)|_seach_blockx_209_goal)|_seach_blockx_210_goal)|_seach_blockx_211_goal)|_seach_blockx_212_goal)|_seach_blockx_213_goal)|_seach_blockx_214_goal)|_seach_blockx_215_goal)|_seach_blockx_216_goal)|_seach_blockx_217_goal)|_seach_blockx_218_goal)|_seach_blockx_219_goal)|_seach_blockx_220_goal)|_seach_blockx_221_goal)|_seach_blockx_222_goal)|_seach_blockx_223_goal)|_seach_blockx_224_goal)|_seach_blockx_225_goal)|_seach_blockx_226_goal)|_seach_blockx_227_goal)|_seach_blockx_228_goal)|_seach_blockx_229_goal)|_seach_blockx_230_goal)|_seach_blockx_231_goal)|_seach_blockx_232_goal)|_seach_blockx_233_goal)|_seach_blockx_234_goal)|_seach_blockx_235_goal)|_seach_blockx_236_goal)|_seach_blockx_237_goal)|_seach_blockx_238_goal)|_seach_blockx_239_goal)|_seach_blockx_240_goal)|_seach_blockx_241_goal)|_seach_blockx_242_goal)|_seach_blockx_243_goal)|_seach_blockx_244_goal)|_seach_blockx_245_goal)|_seach_blockx_246_goal)|_seach_blockx_247_goal)|_seach_blockx_248_goal)|_seach_blockx_249_goal)|_seach_blockx_250_goal)|_seach_blockx_251_goal)|_seach_blockx_252_goal)|_seach_blockx_253_goal)|_seach_blockx_254_goal)|_seach_blockx_255_goal)|_seach_blockx_256_goal)|_seach_blockx_257_goal)|_seach_blockx_258_goal)|_seach_blockx_259_goal)|_seach_blockx_260_goal)|_seach_blockx_261_goal)|_seach_blockx_262_goal)|_seach_blockx_263_goal)|_seach_blockx_264_goal)|_seach_blockx_265_goal)|_seach_blockx_266_goal)|_seach_blockx_267_goal)|_seach_blockx_268_goal)|_seach_blockx_269_goal)|_seach_blockx_270_goal)|_seach_blockx_271_goal)|_seach_blockx_272_goal)|_seach_blockx_273_goal)|_seach_blockx_274_goal)|_seach_blockx_275_goal)|_seach_blockx_276_goal)|_seach_blockx_277_goal)|_seach_blockx_278_goal)|_seach_blockx_279_goal)|_seach_blockx_280_goal)|_seach_blockx_281_goal)|_seach_blockx_282_goal)|_seach_blockx_283_goal)|_seach_blockx_284_goal)|_seach_blockx_285_goal)|_seach_blockx_286_goal)|_seach_blockx_287_goal)|_seach_blockx_288_goal)|_seach_blockx_289_goal)|_seach_blockx_290_goal)|_seach_blockx_291_goal)|_seach_blockx_292_goal)|_seach_blockx_293_goal)|_seach_blockx_294_goal)|_seach_blockx_295_goal)|_seach_blockx_296_goal)|_seach_blockx_297_goal)|_seach_blockx_298_goal)|_seach_blockx_299_goal)|_seach_blockx_300_goal)|_seach_blockx_301_goal)|_seach_blockx_302_goal)|_seach_blockx_303_goal)|_seach_blockx_304_goal)|_seach_blockx_305_goal)|_seach_blockx_306_goal)|_seach_blockx_307_goal)|_seach_blockx_308_goal)|_seach_blockx_309_goal)|_seach_blockx_310_goal)|_seach_blockx_311_goal)|_seach_blockx_312_goal)|_seach_blockx_313_goal)|_seach_blockx_314_goal)|_seach_blockx_315_goal)|_seach_blockx_316_goal)|_seach_blockx_317_goal)|_seach_blockx_318_goal)|_seach_blockx_319_goal)|_seach_blockx_320_goal)|_seach_blockx_321_goal)|_seach_blockx_322_goal)|_seach_blockx_323_goal)|_seach_blockx_324_goal)|_seach_blockx_325_goal)|_seach_blockx_326_goal)|_seach_blockx_327_goal)|_seach_blockx_328_goal)|_seach_blockx_329_goal)|_seach_blockx_330_goal)|_seach_blockx_331_goal)|_seach_blockx_332_goal)|_seach_blockx_333_goal)|_seach_blockx_334_goal)|_seach_blockx_335_goal)|_seach_blockx_336_goal)|_seach_blockx_337_goal)|_seach_blockx_338_goal)|_seach_blockx_339_goal)|_seach_blockx_340_goal)|_seach_blockx_341_goal)|_seach_blockx_342_goal)|_seach_blockx_343_goal)|_seach_blockx_344_goal)|_seach_blockx_345_goal)|_seach_blockx_346_goal)|_seach_blockx_347_goal)|_seach_blockx_348_goal)|_seach_blockx_349_goal)|_seach_blockx_350_goal)|_seach_blockx_351_goal)|_seach_blockx_352_goal)|_seach_blockx_353_goal)|_seach_blockx_354_goal)|_seach_blockx_355_goal)|_seach_blockx_356_goal)|_seach_blockx_357_goal)|_seach_blockx_358_goal)|_seach_blockx_359_goal)|_seach_blockx_360_goal)|_seach_blockx_361_goal)|_seach_blockx_362_goal)|_seach_blockx_363_goal)|_seach_blockx_364_goal)|_seach_blockx_365_goal)|_seach_blockx_366_goal)|_seach_blockx_367_goal)|_seach_blockx_368_goal)|_seach_blockx_369_goal)|_seach_blockx_370_goal)|_seach_blockx_371_goal)|_seach_blockx_372_goal)|_seach_blockx_373_goal)|_seach_blockx_374_goal)|_seach_blockx_375_goal)|_seach_blockx_376_goal)|_seach_blockx_377_goal)|_seach_blockx_378_goal)|_seach_blockx_379_goal)|_seach_blockx_380_goal)|_seach_blockx_381_goal)|_seach_blockx_382_goal)|_seach_blockx_383_goal)|_seach_blockx_384_goal)|_seach_blockx_385_goal)|_seach_blockx_386_goal)|_seach_blockx_387_goal)|_seach_blockx_388_goal)|_seach_blockx_389_goal)|_seach_blockx_390_goal)|_seach_blockx_391_goal)|_seach_blockx_392_goal)|_seach_blockx_393_goal)|_seach_blockx_394_goal)|_seach_blockx_395_goal)|_seach_blockx_396_goal)|_seach_blockx_397_goal)|_seach_blockx_398_goal)|_seach_blockx_399_goal)|_seach_blockx_400_goal)|_seach_blockx_401_goal)|_seach_blockx_402_goal)|_seach_blockx_403_goal)|_seach_blockx_404_goal)|_seach_blockx_405_goal)|_seach_blockx_406_goal)|_seach_blockx_407_goal)|_seach_blockx_408_goal)|_seach_blockx_409_goal)|_seach_blockx_410_goal)|_seach_blockx_411_goal)|_seach_blockx_412_goal)|_seach_blockx_413_goal)|_seach_blockx_414_goal)|_seach_blockx_415_goal)|_seach_blockx_416_goal)|_seach_blockx_417_goal)|_seach_blockx_418_goal)|_seach_blockx_419_goal);
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_0 <= 1'b0;
else if ((_net_1264)) 
      _reg_0 <= (_reg_1|in_do);
end
always @(posedge m_clock or negedge p_reset)
  begin
if (~p_reset)
     _reg_1 <= 1'b0;
else if ((_reg_1)) 
      _reg_1 <= 1'b0;
end
endmodule

/*Produced by NSL Core(version=20211030), IP ARCH, Inc. Mon Jan  9 14:47:40 2023
 Licensed to :EVALUATION USER*/
